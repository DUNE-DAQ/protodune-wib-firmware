// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QLCndKoxh7fSN142Agx4VfdHIkeza1evxb+0EbB0bSq3NkobWqXERDNZOL/fBEJY
GUC3KYCJrrdYTcSS93s/+N9/UPWCDWUM9ZwbO4vQ8FWNcyXX627oQ3C+pIvAUpVw
6vA8zzoBfAoaIu6Cj4CotWodT61nTBeofDa8ddkCXW4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7536)
2uNFqB+1Jxgy7YGmJjHz01iUS0uaoYZVWJIbnpZNvbJk3JcnvjzOiT4Uo6r3SYSd
GN2LJo+7CX7QVlE41nbwvG5rZQ5wfgE2tKWnsKuiL+Ld0DJwumX17ay65pXL7+ZJ
8bIZolqLjph1bdNqGYA3wMWdd7tI77uDg4i9G6dlK2LAxZ2qP3oyZwiY4yMofkCW
ne18R51rv6+kZyUWTch4Ir0JbK85PoK1kiQ58HK4YGospcUgs9tztoy6MfWuAEF8
hfuPTQYTtRzeHmGkynMp5qPF8Y6zgIasjhrDBb/uX1IzF5OU8u9q95/U4jIkB6Rx
Pyr7pYx1xMgU5bVCftnq5WS1RSa80MTJnVRt+rXIqq7v0tSkyHdQ0CCBZb6Wm5AF
weh72gIkdfNr3DVXuSJZ5kZonm/dA5FTsvHmQlUPO+yK3r120KobCmR8BBOI9PVr
O63wiqcQPk7gRxz0PD2skyXqrOkasK25BfwGyp5Teg0jkw5QaV6ezU93dubpySS5
zciMpMDEUf5Xk3bSQ7WSwqoZ3t7E1CIXJb8eA/sxObAfpzbug0b63oMF75JdIdeB
KyuVWgvsFW+gdczoB8TAO7tn2Lsd0sJE7LeAndWGwgjC0VlEEBSKd0Sne2M483r2
gi2veLm0fRk9D0thMXYG1prhhg6bRGM5tda+N4ZR3ijAwjsI0U2j1UwmkC9ZQ+dQ
inNyE1ZpIMmX5nyvZxD8a0jMJBnNpqFYYLmpdBSYqE66jcz3IyU7dLobKOWoQH05
5qlP9p/44YiBwfSV2IijZbbl8lXAf6bd4lXWDIKUZ32+uS08HIA2KQloHA2Ns7KZ
C/TVrDEc610LImaMQAhx336ytwpcOGV8G15uDQgSf6M8faiNY7cw5x60O4nRQ4wL
OIDaE8LXDRbcPO5M8o2VAEyaPIO7Om5G8T0SZYgcQ+B1L4TacFKd+wk4M+/mrJ4w
nz8vTQqS/9Wd9icuNcEt3tHZce735ZDxwnM9Jqt5x1o8sYCnUEqEwpOYdwUarX5N
K+qY6mbwVsXrVRTzYgqiQhX1c5oBO30ZUDYeIcnG6MMGUsvng4VEfzIcsAP3w+K2
myZxtleXX+z6bb36p5tByrcqGBEemcoT8BJ/B4QdNG+j8LQphFvmRMk4XFp82jaE
kG52w7SEmJZF/aHrR3C8yWw958BnygWQzc25nJ5tw36HGvL9xJ5YMFB5bmZsIdZG
tUBtjvkgP4t3YaBxQxANI4sC4N21fjM/pfUlpkkFijgKC4CShh/pGRqR6y/xRGOt
1nXS562mUbciDRwEn2FNWXaiPiQg8nVfptxWenf4BvJlBqW6x2FH1KqTLTQE1ktE
hOwbljSZvOMMPzgWCmsnFKvNrf/qdwAzMmXqIB3tT21IsiMSqMafVmpLrmsiD8Eq
yF3niG1oooa7IBNpqUFjBWpykaLYZ+VrdWCMV9ACH1QCRan4EFcuJDzCtvzOdkIU
kBE0aRxiJ9UG58uXwbbDaAUKgMckuwGR+7i7LFM4ZBJ5ZEy4rm+HfWM9DZuuBh6/
uP4joIKRNh86hg6fW9CWjxB3T6do8bheEFcrsoJQH35Fkktt+AqJEDY2jTd+K1oo
hVd8fmP5i03LAXvtqsbUY8ytnkcx01h8szOTGD4dLZ0B/C21pUR81roub0skSbxS
zIDO0F/zVSDkeyvQuU4aBMRLwndgDURFyUxuY43p5CUGgAJYW0gRlzT2klKPJDhl
GbNXUldXjE96kfV7maM6RUN7V8VYkc6Wmv3mrWx9sT0mRGWVd00NSePNV0pwX6wB
MVqfUpxJLifQEW4Zw3ehzrQCW7V5ba51n2cl+yTp1QC3zzqW5VgYzLnZUI85Cc/N
QIDd4Gfc0jPjJngD0BPu8tXnB9cqYn68WEE+dkB/7DmBzxyI2v9haJ8Dh8P/+rO+
nT3stSD/4yd2UCzvhCoUeHVKqe4WNeUv5q1CTDrJ/HIMgSa5DhAlZnYvxQQIVV6M
2IQzXVmfYngD04A/RLfqlGT+qQ9SMn9GtK7JYk9il5euR71PCsDuGjVsNZm/5srm
yZWzYBnScvmTW6FH7YlfFC2qpU07veJWoFBd1FF7Jbo5I6dtJlKvlxRBJ5CBUAi8
5MkvCZ40+eJrvpd0N4NoUtFv5CPQtMjNUry/+Tvsq+W8QN9VFeg4HUIyOdJ0z12p
Q39j71zv9nNxbVAMdLlCSkavfd2Jrg0xeYFYHEdL3RNw7WjA629g4Z5DMicutMBU
z5VPoKAuEzfaR0spSZHeqFP1Ebv9E76geUrjHhvYqI/4tArgVuNXL+eVwEk0XE5+
f54Wtfb4RxfjM/Xp0taYutz0RwenViy9qGO56mpKCmBNNWDY4hW1YJ0HbbU1/DVx
jIfQwGmVfcydzXB0L2I2g7O+GPhD1mShHi67g4/wedMlroVNVJl3LHREeOOhsXxW
rtZM2d+afzj7VgumXVVcn/IfKWm+BTGoZnZhKYbPUeXUT5AAgrS0/e5bdUS1En0x
IuPMc+VXO6kdjyvSSU/I19SO0re1SisOQtxKlGKr3UNTyHQoAbfBahTBQXGGcF4a
n691tdwFoy2VwzMVtEPPqqFWfMttLDSbaCymJZxfPxuEjibOMKkeMitOThWZHBQC
sULDqWbmCmF/RLVdNfI/Daw71BlfPTgxY2pcmAtHP5s+G7LNo4hVSsAMzmlDbhOy
Yj2MNFMVjFhDU//zbqsWRcbs+DR40pswXI4nHKQgVJZX97bbVxGU5YdATWIam3Zx
DM03gfkTwuwwBOvvhy+cwjtKxeaKqop5JKcIysQhK0LlBRvk/Cp/eBEpxZEcrAEE
ks2j0085di16Utsx+vZYqnJ3vosngXD+vdE3ThyIh8cE14wdpmRTpA9pHISFZnZu
gdN6MD5LAjsD+/HXTnVOmvis282YquzVmdqC72qO6K9V6lh+bptJet73w6sc9aXh
JvEi8Byahj8Pi0xvuuM/1U30eXimNCqZH+7QNmimwsBDLrXM2iAo7iTQKscwNagF
TP8bRK38Y80Ss3XhyzHRUaERw8fALwq8H/sg4YiVPXqZcUqNipFe1OVbbYUKSNOW
wOuI7KG4fy7Jgt5exMUX5/L1kHzaj5zsthsXenQoEo8jnAK0LE6VUlDpKq7iUH2f
GVmvSZZQcf9OOqrX94mvqP5RCteeH+5nj6yhCbwggQkilI49W4YYV4OBDJI+D3Um
vATukcjEqceYWltgRlX8HQWPdEDGCYx2aNjmwdE/nS+lG4U6tfYo4Wj0Xo1UuiX3
Q2VSK/sJ/3rsuefZj2MnBq62MGe3n1+K14I5V8OWS3ojpNq2IU9um2+3qAbNytuc
yKodbJGZbWPYBd9GTIXuXIFpW4x48TF2NrNmnjKizNOGXStUIjvUlT4soBGpSlX1
1dZo9M7z0SMHuX3TC3Q5vmblRMF7zvktK+8g/V+xcNoI0BJG5ytgOSHqHqf1TQsl
ILYSlr4LuCx8Ow00D9Jk5+GoTxPQgsZVk8jlbIBMytIhz3NMBZUvIa3OXl9c54+J
G4jzv4T5zEX63H8Xcbl1j+ZR3kNDm5yiKR2JIMnvUwGWvf7JWjwwXjfVz6nIvpDT
x9yan1QyHPBrsr2gf65MjfpTZxT5ZARI56t1zXgMWgk+DLVOmeEFRdPf4K4MhgcG
AcHnUD5oqxzRRAslOKepD/my0VY0X9xfrZ+7Wb2bNnQjE6CJOLCzjdvuVJqfEyxU
zXm5pyXOTj0HjNkgmbG2mpUpgUGj2ZZ4b+1hDN+vZYDH3use+GctKeGq6tHt8i0a
Ahvq7dD9SaAbGaOZGODasQwcfTXAWaRt1kafvCqYDUIJRdiIfsbZUAtPzCNE2csN
fayJ9cR7UUUpxmI1gC4LfT+ZhdWfBqjrVCJIcTw4x3KsakX5SEMWbvibX14UQtfa
sQH03KvKUiAUvhuVCxxzEONCt9TY1XPLcuBVPRZZLpy4AxNj0xBtLhRRrkaa8UBA
2Uft/FrIKo8cNbAYVTlha3vI49hkG+IkfBEndmWnPEIm5fVaJtr5w8lUBBquHVFV
TyszA69ROicPtbOS6guEhz9EG6QNHCYsY9mNwCI6nKWFcVJpBGKQXuu7AKLqwgjC
DI6bo1/MK2qKeJMbcDE4UyJuy3fqH4cPtBkG8054PL+vr0fndbiG3s6+n8d9SX4A
9c8+u5GzyQZF9VErw/8va2HEwnCO0KQQbbQ7za4j9AbPr6vEAoytxymIwiv9bRu8
QJzjPG3kLyvVP3ceQainGKIJzJsuuZVCwcpxR6Zz5yMm64rA2HBP7pjjDHc9Nivv
wH6QW4Rp0sKhEP/U0wDC3/+B5MxdV3CQoTrgEL3l+SsQaaDNcnN2tRutml9tr8WN
RQlC70um3TY8GUVmpLm+K3yxv3m+ySEO4yWcpnEhNV12pFdNs8h73Ne3dVy3BpBv
OT9EDep8SEn53jxT7ussYRGbo2mjo8zi6uuxgBqJobyR4CoOtC74WjtQZepfNJDn
39XxNhUiz+uyzlUH3Zwf2VyZYX9/8oCH8icf38KNoEoeDYhyqzQ8JuqBeGfErpkc
5uqLjD1ptiIhZoOuFVphnyo2Wo90YI+hoK1NAurc1Y87Uoew6t21lUyRwJjJUlaI
Kb5CE8Zi4Mv5Ac8aYeqLjgjQ4EZPnM7kZVciSmqhjHdiWOJYUVnqZX2aAysNyJUW
0Zn7+WEL7QVxozpwE+NtaDGjsZ25qg65LJxRHf2XFA5OgHvC9SkL8LjDiWEJJjzG
4385a6nvqodzUz8wbhIKDdZ8rKZdHe/QjNGEiMUpgVLWdl/LEOUV6CgIXoDhmJHh
NTBgWu8WZpTua4C0b4jgIkIyBsEMk6FAOpYiEeMYWtc4PR9RVKCEPFVnbvEoVZCW
m5MV/b45k6jfL7UXmmXvJ5prI5+02vop717BYhyvTQKX3V+maaAFThw/B/+5RGJx
RKcH7+McEktQKIMVmLGnjFOt9zMoOXYHONNNt5Q1I3m8KQPVsbAEsVoyL+sEtUki
Z1GP5OVaksyEQMDSUizrCLI5HkhNoRWFW8pDQMgD8Xz1YJV5TT95M6Rp9QUPzXbb
ypci0Y4BOKhm/P41M5t986s5LqRfjBGXSgHk8Zlxbjxqr3DKj71Ai+OrjNrE1Fem
wCEJm+OWItvVWnbTIOsrTvM/bRDaOTy7RuZdxYQ7Elm/APfC7k3akxLuQkWE2J3l
vvm2B6FkfYxZLOP1o87tSnTryFAcvmFNMf62LHEK2OtJp59oMFF2vctTt2HRajjI
Qp1IYg19QwvzMTigmVlNnoMUtntNXfmY/0MLrRqYOPir2hgyI8jjtVzHZCt+QSft
U+58FEBSnNP+BzqQVh5u11xQrS2Etx/ZQeiT00FLgvrM50fP+nPir6A5wE5XzhLR
Xv3ZYFE57OWduqWNqQWc5AvgV5EJvR4bD6cMHtldFforSIWrmiSML17e2vH12+27
C+jTukVzdlpNUJGQ2StR4FVsRG62yJrXrotzLhWog6NJ71GBcMG5H/ntXNeSOVF2
zfOAhDxZS5STT8vAU/d+Xu0i5eq2VSDoLoJT8qK2V0NuqIZzYYrnhlzUfh/2RPwD
7zdqp2VHkhpST6t5aaQDfl5lRZboAO+Zu/hf4n8ZtmVVwuHzdFAmbWikTRifn1S8
SGV+qUBVJNgRLDauI0NFKddF5S0cb+Ky1QXqzM9Ywr1f2saVNUj7QMVa3BwTYQ6p
x7eI+2BTdWUgb8VzSW4i4iVZijwljZfe5VGEXPHTXT0yXQWIR8+iUJEzmZy2YWWE
nYWpn2NTDE8ANOtYyUvllDQ/VFHPNZhC31AiLkyL5Ds+BZWZLtojc0h6QW4zS7pZ
RQZSxXJsSFcGOjOTOJh8cfj97vqiKVby3E57/+hiNi6kROB34FseHq5jP+AIhtE4
pfTFYC+j9fXCX/d/Ii8U6s+P13rq7XgK7wFES9ClFkpZgnPqFJ+m3dgU157axszn
ucfbAfQcs+Jz4IltyoVoLe7TiIC2+xdR8oA8tVuRxQjj42Wu2+x/gphL0L4uMjZj
Fl6wFrt7CVfwihL9Re+bAJ3IhW51EPkxeYnOj+WZccn+w89pIrt+kr1vnmeRwJ1s
ARaOv4yv0av/fPUgICHvBgMdrePiAUxFj58C24/ouKwYk2avsVt7p+Ig+8SQzmi4
fx5pjQapLtFnYE6BCKmcOxjzPbhpFI/zmAIsyRsJ4OKqKgJIv7hIAn3rSwuSCXDF
7hzXAl1YMnKgHNyPHoKc4dW+OyhFccRl3IAdmtRZE+nmzS1p6gbgJtFAvo4pXdAV
j2ix8Qu1x5ZX1/rFGMEsmD0WfahpXuppFijALvuDRTQcQTdi4+bcov/ehwKfuomp
z7XEV+Q02mN/sr7XlDfyxRUc625G66r8QsyOdUx/7XJsQWD+WSjjIWJ+A3A0qFIc
hw3GTQhnfmttxkO5L8Q+qYl50QjxCTrIj0ZwgMfMhbWrk0xfRAC/Zsp69pVc0FIA
9Thhtr5mKJfJeqsaQz6Ut3s3Ng3Q+fnUawLQjkavY/8bL3lX+EOaoGDpmeLatXU2
vlivKQ5+WIA4J5LX6qrKFQaAxvZ7y2VT6PEzH8OlZsORRnsMv5mVuUWuwFM97cUq
BKT7z25wAgzVuAhfpRqADawCe3NKkTJYMgK6e4oasVgC3RC0XGbdWM+TRkFiFGSm
Dro5cI3TEC28x+VdSa8Os/J7URWVe33lOMg4++AoGnoT1RXf6VjlDxZLRq0fTJO+
xKafA/goh3EfleQZiN7W3peYGgLSc1vTV9OA6E1VbsQ7lToPv387ga0gPwkILeaS
flxtnAstr7DzEI6SH5c3NWVTJ7W6WWnZ2hUKY49nqkNT7ax1PW3uEUsZRnl0Shxg
WbXfcraQeVsI5+7dkzrvbKaCrJHrLrR+J0LT5GNSF6yjlVfgTU1m3EamUr9XYe++
ViYtavQWxJNfmAtjKOS5eDnbijv9ZSkoOFI8aDRE8GrWm68j6bT4mGA9nqDi1x3/
OC6DL22bcEAy/EpY3rlyc4oszWuPMiMBh8jLlfON1E16XxjV47dBGDZr40xcS9jy
GoBG7inFGt1z3pr/Ts/25XQ7EJJ4KaTt+vCO+UQEIX4U7GKF2WK3aLTgLoKzx+pa
K9SQRInEVtlLSwTiSwNJAljbyDoTXK2TzpWVxHtjq9l6uaf49R4Sa8AP8w/ZdA+K
zFoiXYQVWUvZtZxGmkD6X/3lO3FY0MqVwK6BYfy870l+bOjAuucJ8xQEI+qvyUhh
I8te1aQ0tG0ZeWWeJ4AGKp/yaCasjbwo84yeOmXFeJYUh2+cjIgkj3K507ZTWwZY
Gc+BMH84KOKD8KwBVt7ifzLrARoxTSSV0si2qZWk9GNeJlrkJ++UGMY2jwn0NmHZ
rvuH6+TOJLX81+/1ZbaM9j+lqR2gKJgj74MMMaI2hq6y6FTrk+2MA8fGXErk3olB
bSXU+TD3x8MT0sEqk8iC4gKarFD9/BiMaEqKTKbqU1iZMy/cG42THNNUbNjMQ/3c
zfNrbqd8YbRsaonWY2PurovuQGKmRpsEGRDwL9sOwgh15h4aqPJeJ+xvhJXOIZxx
M2Itq+HqqU6ETCKIaeKOsZXzTgduOTXEd8hTqQ3lHx8b9mm+Oc6/mks0sZXlxTrL
eTy47zjAQbVSNjVVX9ohT9PBdCaw8gGXnGu4YQDqJ+f4K2vU5uHg8hmPubIG88Um
yNWd5L0Wc0f8fb2EHSjrCl4etWnvtxra7nMaCpkFEHyIrKS6EKdrgMaWk/y5o173
Vpc/Fwt8d5b1laFtFi/gJpd4XDeJES22zASYrovRUI7n3RqzmfLbPo7w3TTK8jT9
X72b86Aa23nbZOiUfrv8D4cnMHBGs8imLqulAtxI2ZQdaomE3DqvLR/GbiFzy/o0
u0yEakbl7Cz269RXhzE4Gwk+5fnslp33q9FxhiATAOjJC8KULTt1HdnAH6YPr0pB
nW1wCAY1rEGy9ArBxf4V7gHQ4MHIP9YhJeA4aSPHYdkOvHjDsJ72bfFkxuw48uN0
NZY8WHrl6022gC88Q0UXL22J2crUXamz32IIpLuI9xRGtKUcUEuZwdMLmx0mnO/7
u3xx2yLo110hCSdlrc6iA7o8WQBUjDwaGZ2C7EM9fEzQ15SKeqGAeG0nXEMEzSqZ
p+VoBZxlk9FM23VtLlkQ6gVYcm/Mcdkkq66d36itdBE64XJX7/IhzIsVgSzE23XP
sVs1tSzRd7ZemjYpwmBUrTC8ABi97UsCSUiVlUltJxtt4rGcHBiypRaDGy152Jk5
Tx8ffl6KvcIJ//OFvXtsrcBsUJSO0XHKhtWepxqH6DQ8dCoK1ir+CSmEl3dCF5Fo
/OhvgXkAuI2UZyC1x3UT/R8BkcRMZkMMmQR21urXO00lkD/L+6neZOIirZYd1n4v
A3q10cZk2SD88cq25/sTXVwK4WNOxpq7J3tc98VLKYropC1mTIZQ6nKrgkFWKrqw
3yu+Wxs7NT7UXOn+9La7dJ+XypXVwpIk9eE4HhR/oJPII/L596cQJfYeIu5vkLlJ
CG4gRSK7NmbcWnNr1obGo4vXbr1xQ1XXX0M619KfnKNPP9oE7bBdp+ykct8Ddtbz
O0Z7521jybYvjmDS+aSoqdVi3MH/Gr0WkzoxcwuiN0b8uamOGNTfMX+ZOrSc836S
ZNw9tJJjH0uBiWkOojJpXvRQGWyDpvQF6zsv8lcwzehAbEIR/BVHvuzXIOiiIjrf
b/5P5e+rRV6lo7B2Yqai0fqJkiPUXwimGrQtf8x67zh+dIZ0VZM+deKYLgUXvOnz
oeYqMQqzGyFDayTc7OgatMg+GVfy0YrIdAFVolIDg3J6BbtqJ1Rv2Xry6dQB2qif
rjVGAAMYoYQqTxgI6HBokB4dJUaeAiOaORYPY3nDfxgloUnVxQnZ3DDLANwrT/Wi
dIp959FnvFyhlRhnGGK9g8wk5I6DnbaNLRR5rW6QY7ms9e4TkqRu7IMbQF2lfJ//
XG/JVifs4Sxn2Ah2LubKewEGbS4pjEC2e8tMpWnXjQH2AwXWuDK8UN+DlF7jI1//
JXvXH/QuUA7BvXeqqakkxmwu9JBefXseptXvwlEAdrbdqA66bcduH5Q0sqq93L1Z
6+8OHiVHBOXoQVqBSfEBRCpHjjN7kf1vITLIrzFLnhogxkhNX6fXQFfDvJ4VzxHm
QZbO9tf9PcXNSjNy7eedPcROarCz+fkNTkyvJdocnMCkPoRY8ozR1PHG2eChnn6R
B7v4mYthpQg8HqAlgqRN2oWNj54wXf6BpHcworqWwRjBVxSAB+o/pcoBmtU2az/N
io0zPHKKZu9X19ZHCejxUdEJmaLFIpmAyYUexeT8M5iXFwII1/9vX83IjXqnZibV
uJjGJ3T7AgpcW0lHUKS6H2mvf2lBifbuW5e2i/wmCn7OZbNUhS13EVzPHRWx9J/V
gv/vTSMd194wkbUIM3/1SpVCOceHuAK0/wdbywFgb9xwKpesqpO/ZktFnVoy3GlX
krGTbsK267Qd3q3CJPFKo0VA00MVvu9YwKr49otCiNzTcWPgolft5Vh/7DE/R0rN
7Nt9nE29/3bstWo3S2CcZXaRMt47idllAMNX5s7/KcezKZ33l0rUXmRoFQqPK2dC
SyBM7L2AqnN6363mDg1YjMcfy/Pyh9J5fQ9hj9BhWmoPJmbAAyj9Cqx5cdpY5hjf
81ZrU+Svo+6HJRbNwJD5HuUGu1iQe1cXNl/O5N8bIFfFNDSWEmqVp1tPtJwdkkae
XMuqMukdf2fDou1oITiZIG2wPi//mp46LzEqxxF+cXtgOHLVZpX9xTznCPbWgVlG
bgcWfZ+aI4dd9pNQJpacOtrFgpJe2sC5gZjHXCgzNHtZA2AnOednNSMhtk0wbLjE
I90hG0sDG0aok278wX40tFQCocgRZE+ymyEHIDF2JuqLVu/gF2eM0JTf/razEGJt
FoJAAwlv+kYWch/eplKdOJjQxPgQXxmDjlhzGr39roLEAymReLC2svzMGnRGRhq5
MzneLamS2RxDdtb3IR0B0fjrqY2zmxt+M4IBi7JYhG/KY2WhlKg/O3vw8ufoy2Ou
`pragma protect end_protected
