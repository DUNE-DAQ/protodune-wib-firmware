// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EAgpPoFCOh7ztTgFrn7TDeukzx5oF2v8bx0t7r8RacAULX0D1nrEE6VTvdZ319AJ
Rque7Ixjy2DAM8GmdmqTOzA4UZL1SrXZ9IMYqWlBya/sHa/zLYSsN7iHihT/GUHQ
nE06jE5EN4nOb/dxiNZLYwKc36s7oIpxjO/WSzpm1Is=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15376)
5Uw3NCVdMBO7D3f7gvWJ8LKx/myB36LMXi52FIAXS1hWu8ZF6eui5PGF3mBBtrqK
KZxu8XxiPnsvQTUD+3J6of6G6WwawZoP3V4Azs1kV/KGddJr+ifPT9WA3bgp/WY9
QDuJ6aRR3czrXEVl2LR4KAMvdCvn4FyVLHPdkshI6s7Qqk3Kk6fxoPjTqsiFqZW2
fHdqIaJOjmLyRGXRKxF+YaIHDuKx2pSeD4s98g/4KXQgJc+mW+mXX/x+2zzcfki0
v3j8skCWO3wPUYTTpDC0Kq1T14nyJTKWZeER8xtjWxpXQvWCxpxB6FjEvApsweCu
YHg+EdQ8OQmXm404sR7J6GFVitN0wmNV242nWq5cR5Yzcec5UsKynB/169P/8k9m
ZbDXk3R5OTc4LSv8+XUQ//FcJW21JLl4z2jJ1S29RPojPDV7ulozVWeKIkSFLs8a
36JnKN/CQnvcXnsRfKCnboFRbykNI51isfPvKpPZ/8tRIltYGI2KTG/ohrg2lao8
02ndl+V300lTvtpTXPp56JvGvYjG1hqpGGAtKsbJnlF2NP5avcBhU9MamtkEMfar
LWBbuSTvL319YnMLrqxdJlmJku6LDfnSNPuv5sqTckB5C1vZr+aosUpm0mQPoQUf
QAZipsQGIGge/bMLBaezBqECH9BOYncDYTeZRa6DVpap7ybziLVwHsMqDVENz+qF
rOicLU8PeS8b5fpezZo8YVvrt1Avdd+6IS3NCMKABv9+kA64i0CWwdhz15D0MZAn
2WqQQNmLdD6Mrc7WJ6D+G0ZvYuDw4RvnxENs4wpH3QG9eDjCj+J0DWkI8ctJMzT6
E9mxLJvhT4e9YEpjdPY/kN2vjYu6XO+dhEJ8qYT3xzdhwnFVT8jH+KgyxEf4xiQY
SkiuPYvhoDdi74Op5TSLSrOTM0cNL9IaF7mBGdQInxK60UHdJZ+i4Y/LTxCJVHCA
FVaYJLxr9HwdLOVma1v+vge/Uq7FI9s+V3nSy84B36ghF2awi6Stv1v1rmh2DVT9
/cBUWFUadaOifa/L3+u3nxRzO/XLZju7gZaPk/y2WM3XKoc/jRbvmk/lGh3PzHly
2HaLghAuhEOw/UH7iu1wfffp4V1EcwsQMWnmWnSuEz5tJrwD60rLM98p3pmUgIfP
Kq3YKL8kIjBqOyOLgNq7gTl1c5HBlke/8ikzX6EL6WUQcRJC/Ok4ZJQgih4JY8fV
fGYZ4DEmHvsTq1I4W7V/zkqlfXt+rSV89ekBkL0wNsjaYp70J3KdKXaPeYEK17tJ
hBcpcn0BKGKvdJy6zmXRmTiPCKjnIRHuSH6VH/evvlaHcCEPTxOm6YxrtMBIuADa
pJOZDVQJemTOdsF0ooQ9hXU/WRTytp8x1/RTGHFoZyP5dafdQHqCjcPF14QvqZgo
8YfDFJQVdDh8T0fifFck2UGoBpLQE77UGFY7Cv9mGEQA5EsDaBaDu4auRU/djK35
rR0WY/NNMxUV4ICKUeVSXzM4SrmA9gvG06OtQ4YNU3T5P5kC/t18nMfsfXA/YR8e
iAurzr9qZhwENsIIgSEsd76JuiR2vN8yFZ9qod5+T4eVCxv5O/Tdpm8/o42PvGKq
7B7GTYAKncxt9aJu4bmKSfx9owEy0ci/rjhOLzgKqXJX3drhTjKkNZwpNZU7PAjy
cPI8/htjCRWi092SEEnnX1aeloQ9MDvftvs6/OSgPUshynwZzpI0nYFKlQ5yexq2
k9YevPE02XOuoua6CBq/snbMA6pq14aGIivvNEqWPNo+sqRnyOaL5u0O51fAJgcB
3BWMLduWO6q+FuyWrUc78S6TnSBh8Jz1Ki7KGCZkPD8I7wf9pob1Nu21Cekyh9bL
Q86irYiDbfppnv02JXwZQaxIwE4Cwcx4ECE85yfaCQ+tj1iJLl5zRwwREHMufnhm
VcWEX17uH3rp2VXVS1EaxOd30jA8Sx4VXX6EmZHcbK+bdmL44kd4IJZv9B9Cm8YH
YUQCIMswOC83016H1q36HAc0vcazOt0LgPs79eTNE4WJWe4vNMjfyxov0TdXA020
tzmu07ooXdqCUWLrfyfFYF6++eJ1ZjzT7I8XfejdXXuBBtQqTXUkCskiThR/YmCS
XOKdlllJp+HUTldH0PIZlhCNOaivwO9HjqKCe/ypBBWT5n1Xe+aEnyDBD4cfIoDO
JISj6JHF9kLQ1Gv6gsQETHBT5N7xtcdjroQLAWpEIoRiQRRYHwpM9MXrbVYEVL0G
maS7hay+GPUrFYE5ELOOG5ulxQdrb+gRtOgOgNvepfyC6L9SXvcyLLKW50Pzjvsd
Hc4zKQgLPFq2gPswLuSKVm1PDGpMcIkiqLIEYkosc/JcaWcN/McFWQ2xoRZ/vini
SRnibu3XY+3UxVuz1LFF4jwMHGqcFAZtVnrP8fqUGDe4blzxhcs8PdLQVkf0LfQ3
AsdlPwy+Nmt3TmJux8ohi5iiUp1OVsH7QT7Hb5U7N+1oprXB55kaj2aKubaxOrwI
1EYtAraWDLUbRw9YjKiLBDjZ+VRJQLm9TMMb4hGNeof0D2p4BGdG+LBDuAc4oBg0
ixpFDFpLQBjoFZLRk+c/wa+lFndACkPxTdFO8LrYt4b2O8MjOl6HZf36G75GPDiK
Ccao7JsX8DgPgoucTJQbgIzwcy2LnTgw/idJh7PGYQkCYb7zV6tkvkgL9pPKfSCI
bnsSoU7eAQrT4jm4AhnpqpMsR7wKbjx0KPGbMHAsWE5tk33Q3cgqlKVFRy0944/B
4Y9DMegRpar7yzokc18TdfVIXaARPf70J37u/jn8MJBUGvBdPZ87XoSmOQdp5B9+
pjKHjusAXVv4OYcXvNmhOGBm/oj80tw7XGqJqBVj00Uplb7nauEvu3vMcXTpxG4T
KF8XRVWA48/jC0bRcWXzaKOZaQMdwUKx0ZoD/zcmk9rQ3ALGMUPJre1HcFgXYga+
1K1EBnbb26tWG46s081XnEUdSGV+6UpUb2fJW6/ydrbCKqCmB5l03+lmt911Ax17
RSl5bpnkCdN2HENZZVI3dc8c4Ee8b90Rv94rE748r2n5cesqMhbG3pCNZGvqbLfD
ta7frYrOq3mAoq7/PdO2yuBCCUA4n/Hpq9aImjy9/DHILtb1S2teQsOzp1OoTFOs
hUH3ndpHd79tdXkSFOj0ZefvJV4NyACX3kjh9EDKo+DF3PIW3CXn1kWxG+y/3gi6
cQtXTcau12tBHw7wkyKTmWs9KTyzJnz7m5d2csO6wVhSQtE1YWD3xhrYH3UMfOG0
Ydi4m8rj75lMnZ1l15HK2RGmMpH5nGqf/9bpfw98eTfFosXJa3l46DvfQiV7Ednp
SJ80XIZQWoriDkFrvHPvJvKHbAK+UOjjTENHVB5Mel0lhoeQSMhSYYz57Itb1Am0
K+jkX4WgQPWeWR5ujmmclHsIWeA/GBfmx6aGsP0T1n3Zs+UBo0OmSU/qJOPdEgOB
olWPn7Pkg3oMI9WCXt0BWYKDT7XlGigmHEtoeAIfYvBB6hq5AEZRVWvJFjtpSws/
NB272Ppv8zmu/Mia61qbgAma+1X44SbNV5ErMCARAae+mK70LgJy5T49GBZjsRn1
n8JwKpytH7cyxrtMlNx07ZgZdbTy7wPObiVM1jpl1bmFmKh9h/H/LOKU9Pg3kkmt
g/uj2RiN3mKJdlk8R6l+FGKIAJKX9VNrd+PkxHWZR8B5WppMuY+XPAYMKsx+tclZ
tfhMQJwpSyh5SttvdNqzItu4p9HESwd/SvkoO/c0VrmC1pz6NS4SuxCuNU0vDosp
jAFiQEpEYzWcw+0j0X6MD76l3I2vdD90iBLbqsCQ9X7Oh9qDdXz4iLDuj0NluTmB
7LMZrZDwpZ+Vsivho1VGCSLftVgp3ot6UOI4K7LOQhCreoYf0d7aSpOP/Gz9XBEH
7bBT/9Nhwt2QIIiTjLa4J5V3OT5Z+UK93PenIFgfduRIk/PlqmxqYicvGX2J8Io7
std/iVULXgQOtQZIpRYLjXkPBleFlfsa/1FHC+w38w8Hsa2b6nFsRHd2Vh2eJdwV
LAxyWmSP/lXsgCxIhiVfwC84TtMDpsz6bZUOJnKMEJDgg5WEEs+prEMhKR6KT4nN
LgdOvMj+sQGUG+UMHrj7WpdFKY7Mt9YB0sR95qUxLtUXMBiYxOIlYhg8VBsIqQBN
nSOvXGTK5b0G0rE35RmFrUAGCYMaijil/ECz+AZ4bLjy6lmktn8QThQqc1mRj+ND
PANfHwujrer2gg3nuxOQVsLA+O6uCxSZkNt7rLyOkHrr4VDonOWolaqMk/bsVitB
xD9uDjowWMkfVa10N1ol2Q8cyUFEXyz5hZePMhEcHx/lR56uXQhWc0RvrDZndPo5
/rvpH5gGSMSHUzxaL/tWrMhaJ+2o1vP22M+CMM/4wYwM78bDuz1/tvPJhbt86UB+
mul4pZUcQltSm8mVMQt/lIWYLWN38G/7IeMeVweseg7uHwR0NOMosM4Zyystfn5A
i9/f38eA1Z7Ad053H/jEvfRsBeZuPv93ENcoa+9acoOc+p2ue0lz4CaVCraU0Uw9
lrHcHJAfMBOP5MUtwZtPr2bB+8vjzzuuqIyvpyMw0wv+hFVFcA7fYx534tjrL01L
rUfgTliMK9vEE0AijsdpDn9u5XbrcZQxrAYo54Zw5OE/hQzV3FqGRmXtoKVRDiA1
wKxhXf2slhN0HIja8eqSrN6rX3FHR87IHjMtfO3LulFKoSXYwPbwijJ/GcIiGba7
XD5/pceQjR9xyJ8G/orp6uck/g2C1eYaM2zsurYBIGsaqNI2usxXws5M6jkmsQio
4614R5kAhyWQCa/8t3edKi0RFBFXXmK2K2DXHyFi428xYyPP0m5eiBM75FxSKQHx
6HiU43mZM/g39x07tdhFEQvNkOgXxg1kjpral8xGy5Ltr14c0q5ZgdYyhQrW2RAi
MbNwbMtMQpp8BxPN0SL5GmndtnYClCh2TN1mgWHIZTPp6miG+JtBKyCMmt7CKRUk
V5mfH+dAYTM6Avcny4U3zjT4wX3YAiWCrTnrZk6ttHlftqZT9skHeNOXh1M0tEnS
xTc0RNDQiZO7VJGPZVSWAzAalO6bOIyWx1SjprnTYpUCoXdEaS5r428qpSW7vcyZ
P+sNHmeg4ZnTytGjUz8Ff2UoiI6LG1wq3I1D2MKjeUWR6MKsFNfXUrYiHnq3Tupv
2NN2oqe00vhFQxzS4vlYGsUoI9wnHrqSyY9roaaTv49Ynapzley4m2E82p+BT2mo
kVot2yYZJEYnUZa5seHWEswz4ad9qFbuIbquhGjzd75JQKQie6kgQb0iX7IaRvb9
YzcxJwxzhpGy76CltzIdcbQGa0/nqcXrqv7FaGFAxgg+aK/kbLj4lpsJYA/S4qZ8
0rWV7Q6h+yYtnPCqQAfZl52bmLKNbpfWa7LrSbDOKroTJO9ObLnTcMZcc2BBat+b
oiB6mCGmRIQh6AXaGXUEsqG7E+fYgKwsR3Tpn13jv1zete3/7fbdJO3rnGtOy67q
XnKdPHB5DGID+qYTqYtqFkuzwSo0fC1ZWOQA63jjCzgYh+NV/JjJWqe8Xl8AhD7v
qY8QrK4TKaPpz6smjyPTPNOzhzqFPPR/+qxZQfeeELWv9QumGYAjeHkEXsUs+rOI
AcgXUSZeI8WVp9vN1J13eGjFs/3w+pKxd5fVxFg6fzZa27R0IRA3MPxqc4UBydNU
EXohIHHk8gS/J84150UE3e5kOkmKXTSGRhuT/zz848Pi5m6IcjW4XYcTMZMseWtY
mwUxBb6rGRsHnhsbOuYrePowDNgUM8U8NvPQKshg6e1PDNMm+eg9+g4Hum5KCvqU
EHwAwCewvE8X3D0SGY1QQBfxhkR023box1AB93jvStKSXfUpcj4s2lmMuZ9xeiro
4A1Sk7Ctq2BM3Vg3NYiApcmyCKGgn0jdaySS3fzTU5dekHTRdocIVvNfYxlbHBdc
1IgXIMRLWxpPoSKvG3YmXo2j/Bi+0SWo+YPjsm/CCfUZ9ac1S1aMzF4CKC4nHzhY
baBHynqnETaFbqdilqQxvVzSOjpXZRaDJca5JVK/rnSVp6vWahsFpYRwKH5C+9jw
GWXawBcnSMw5ebTn4S1wogLOoSMdNxAfdC73KvDyVP00E2TMSryYuxhlH24/RiXn
kKOJFzXvOHlaA2T4Wp9mZq5y7dasTBrvQje64r5xmKzS6G5udZiIey1sYK7iZ1mj
6NH2ERXlPQtz/PmviFbuX41tPMnLtgJXPKWDbDXLgpmnee5lPtOwMHkcTgyYm1EZ
RAPh6C1onZmqkmcSVajaD2P5dLQXCxsHcNqRo/CEreTbAkXYbkpEM/ESDRxrt2ie
460XcRqza4ujqrh9rtskwC6eu1Nd/5fgbiw7CXXffHOyhIP/+uXd7edbV+ELuBg2
h7eGgQKBhmc8GxrYUGWXBSpibUahukcvh9sQigpnKXcsZ+vISTiie4kASmD1f/GS
udvtbN4m7uAjWYvpOXIDMApBDCXsTBu7p7I5/E2eNf+ff6UrifP+G5OJQE+EzRpd
PmCxd8h+7yhPdLMt9DrXebIFy7rl4ZwX5MRZv7kf1UI1aviCPUVDlc8Ujh8bjJaY
PO2CfTAjaCgIt3O9g3M00P9JiBtU+1s2LTGohHtYtk8d3YsCZ6LYv0BOWex0u8b0
lxobicu/d29GPV7dmeJNpNpApaR3BnDtviyLVCtfNDZ3DssDWUIK+cbuzdVfqWTF
o1SVGZrGLSDaaf7HNvzhczkiWJhM6JDd5ilPjA2GsJ6xznDtuJxAs74BIASCT7lA
2YgB+z3g/aJIdXxXcEjC6D933tE5LSYsh/0HKY5K4T6b8eKWaiBIFpel4GFYcASm
90iTNJAjg/e0KUO6flehPOu5TcAPhz8xJL3vuueqx5BnpJAwAHLkdAz78gytkVE2
Wnj8p1BgeqREmlGvTwS+Iw05+2XZEfSLQBnB4by4z79nPPM1sf+PSZbgOB3YFKhK
EEj1Qyl+lSC0cn2SLkRrHYja789KbfKBk3OK9KsC+YQzo+KoRJgvLR0RpPLDgE94
2xiGEaQjoxZcbbuTkkGbrBGkClxOx9/Z5pCG+bEPCx9rCvzMMxatqca02DQ7e6Wv
KDpPmOZnunU9344N3bs+mZdaT0RrRuBwODFOaPdaRx2H1DXqnRnLoJnGm4odGgh6
uH2t0DQuW7s8496NIXlfqz2qDM/mgjHZ4tskhPMmoazKDIV8K+hQnwTd8zlFNTC1
k9iYgQOW09QtRQBdK24jGEhFoZKWn8o+aP8vu65I4Jwe04KRX03p8D97DTu3moPS
qmQouLQU6y1cEbLaNJNKi+zBUCWIwx7GMTA+5pnpK3JfKaZVJFP/cUw7I1JIuoVg
l1h9NcMpP5EF/kjb2FLM4yzXxgNBY8HufbV6ryhTf0HpDtQ4P1f61DXtJcqWCVxq
3k0sjLgGlFFXZq00LmJhBg2B21THleyQ+7OVhtOOih/vE6CFkLdxFUl6AwjCWaM0
bj9xLkhkCkv27gf3AUsFPcicHDCWNVT9Fg8Xu+Hn1skMU6aOUd2Lh2JeSkWDAJOk
pMVAkI+s3frJSR3WHQmVo838wSlSJpEt7fMC3NIzBvVz9oYV8mS6MVgXQDmnX7ZM
JCNyPVt0JgRDuNHQ9rWJPM1wNWidWtPiCIQg8ynsb71ukHhquGsazcvqdHSE947v
s4jt7NhmVrN3H0sGCU1m8SHkQLZaJRZMWVQXp6rIKn0rfm/b7RvPj0aFkBZuzpNo
Mj8z0kNJtM61R5GRv5PEgt6Xo/m2HHk9fZLBIpRg+l0z4ZH11yiqART5zlJ/kmNr
mJ9M8Js4q0nZ71zjYf+rNtnxIpOcnS0boOkeSHLIFJVsLfDOmhnBiFlfIttce62p
Gh+WSyjDFUazbzm7cfFTOiO7OsAahxxcuG339jBFgJAJg7y4wPakXUotYaOATEew
/kFXCQYYPRfWHHG/YaQojlhPBxqTpcFFcBOOyichzXCe1rJTKN6MMjBhMqnJdX6Q
x6ZdyLRA29JGAm55va5XfMZdGBfqnVXvnx4IiyIXkjzF81syzaq4RKmmsCXG4EBM
Ks62Mnha/5qegQEYaf4eNJ5ae/hlIiNbwYgzJjGLtlgJ3JSib1YxqsSqTHE/gub2
zkFxgj4QQD1cinuMcpJIMM0gPdcjI19qHjsoG/LGK4m5mlfJCA+IaGmBLZfNgPto
utMxrz9PQkvEFTOFTOHg2N38U1qJyDpG1MtZvF/VpCEGP5gHaFJt2Yqf7HWld5Fp
/tpPVpQCDOiZwioJTgvsVbYreIFGcYh9UvTgQg+1eBaI/XHyo//r9LU67+xdnW8C
6ZYGmlQhPqXzZqf2betO2xjdtx82R+HmEK12P1M6Paruifo+u/3CYmF1wKhM/Th8
8YNl/TaNvalc7az6dSIpz9hjb7Yt7D0yt/D2Z30Pa4VJKXs5D2dtU/Z3txHY7YMO
G8UtXIsuSNw2bkHWJUbpTo3Go78W9Auw9D6Gyt8VsCjEyQ6bZ89Vw0MA/5BFjdHs
dpAsj+0SNxCHuV3c+HOwQyTFlv4b40jNHFpLVpfqKE2rBExJ0k60hLQpNc3HlLgN
IxWiJNejyAEI1fLyoDWxanzS/odEQxKvaidPvJoHpGLY4ltqdq9eyOdQtorPQKh2
DrsE5SqjO1+JhCyTX+zJYGWqbShpI76OEwJECQIUTkJRaYb8u8P9RqezSOmKZjNx
qhBBIdiOl3EaS/HYQoAieIryKWBIQy9zViBhZdbt6p9vGdW60mMNaD8v26QGNi6s
41IIRG2SvwFlfGo/Fb+f6Hckm5W+wKfO8RD9OeyPz58Sqwl0tsDGEBQo9Dtj4Brq
Ne5qYB9KylWZme501XSs/ZblRmd7hC99lnKJpN8ICSxPziQ4U09NQHCMWXLqR/51
ygr3dCTPAzd1rujyHxlho48iJJQo9PtprQt3/4DtbdgIRBFMCN4ePSsxCZAfpWt4
EjKYWFBKJmwCRMsU6inBi01AAid6QeMDDlV8brJ5JBqjvoMv2NloF5FVZ/HDSu0I
KuJTyl6Y5dcsJ8ePdwb+vm7sRPMQaOx9t0JQguLIwSgy/VVaUb+YhBLlGAqj/hgT
a1KB/igBTsz36LRFJz6UHW04xFsF7dh0t23/HZj1J9Bsa4cierVkEIH/HnfGErQh
X5OHegygFiqUVN0l6bZdKVKm6TxJgL55qhXdlKxaX9DTmM3WNrxyGd2Bu/5adAJl
1LJXYPA4VYKwX/nEb0wrVJgIRV09g546YxIUGqbhiFlPeQqSexph9QjFTsDj4yso
y6c/NX0REos1z4Vg14K5/iVi0lEvLhmX4mphvOwMtLlkuurjRrV6H0r+/i6RRiOv
MbdyKgwqf+xPHN5EWCFmdyRC4049hF+cUvDuxiF34KfQkXN+iuYp96eykNggJDtq
gvEcfvaLapRinwGsPIDYFhf13/chpqRUYvgBi0zVKyhxEXXHfWznchRqYjqKU1Nk
IzHx9z3GKgcjP3evCLSDwdAfQzEbz4ynBJNTvcavhqHdjmWh1f+iVb/nYotsiUdH
awcyhutsDkGXa3O7CjvMG/UZy3HZbgn3bf3AZB3ukZss97KW6EM8EyQbSwaJfgds
8QR8kx+rzzG4HdPkw4A/J1YY3PwjgqLAD/NYDeFSwgExwtuDY/j39JhVNA4HRJC8
vtF5rDw+isiL5F7paPPisMjpyKR94SAenk6s0K21Es6U/ZBLdqt+D2DJjCnwiga/
IclHQqWvqGxUdTKbZIBNcfkJ/Ad0rrUkayUjp3fEAOhRr7WiTUJCxzEXltw/gvEK
Ld0Xeqlarc/UDqw9hLK/fzdf+Jo36O7pNlAKfzgFX0DJn4Tl4vjx5m9zcXmQs3mk
jk82Nq7cmcfuLrAV4VBwAYS5u97z1gBAE5hFHoMYc0mpd8qpfEHkjdDGlJn2z5s6
O7xiBBDNANGoRUVWQDPBBkhuwAThDkpBs08JLUpaJIDXEqTW5Smli6YXp1cE3E9s
qfxwVvKQkeO0z2dsmLxj3IW625EAMam32TIiP+IRKzgNMHWlyN6Y+MHVeC7AAyjh
y5w5u1HL9CxLMM1aKjzgFyMmhY+hp/8vc6YWMVY9H/I5ZVT7kMqQfHwq9Kyoskfl
R4PZ0UzzooPHM7eXnktDC9zXm5BpT8eInr2L0Bjira+cjqeqSG/YwDebhoSjNyi0
dgc8CISEpIxCvtCh0iyZwU5Rg/oQwdgPIT6Uo2GvVls4a9932HggnmBZVth6xEYI
OQNIOyE0O1mgDetzWIpyoRnC40uYp7Qnfj82N0wnM+KtaP2aZvIvjiwimarY7f+r
hf+gNHdWxMHo/V448IsKxLLe7ryTzM+BEbNFw5QgLN3ZjoGFb8tgWwt6JsBL21ef
6docF6laYLJ1hFfZvK7gEHeUgjMF6IDbE1IOe0da/Z0VrzBTtkgXvWAGMkAn4XQL
OUDuyfrV1eF9xHq6S/zVC5WkLGUrkFIqOEU/yzvj3tu6lqweATCWVX2tJFMMtpko
oIJb/wlaxbNCPgSPSNhQJ9LuzE2e0U+TnvFtLuOzr4oh6z8bibLbrYRK+Z7yCtBU
JNvVKYWZcvnWwUSax8IT1mHO0+ZiQjSdvip/GmxMjkYhhXfI9xcGkRf5ynA34RZR
2bQZjS42W/ThWJa+j6ZBbCgI+Qce6y9a1hpFnNPhBJrpaX/9AmNknofdm8ypKgK1
TT0kaFf4Mpjzc+O272uZ5FKTH+Uv9XUqaA83/SET0AGYxuY8paBmjBkg02w+0tuM
ek4gR2dU9zS61ARH4J1FGGBlvnPUkTV1z3Sc7j7eyq9hsLGA4K8UEyUM1uecQO1k
v5lzat/wfPLHAlTqN348efFc/FD2hawAoTxlyxWsG1mBhjVLtlunD6P1j2gZMyuE
S3cqFyMEiADA06fQIdU/x2gbrqzx9IBgzzOvKC3Do01D+XVs8Gi9Tc+XQoQkblN2
M3hf+eYuiyp+9egT2VNByPPHW/+Y36wAqlP8GDfkJbjJn0F4EshvWsPTk8sA6GOB
4mWM3qcFyljXUbVJdrOY+VslMHH1VDSeOrBW0U/6B12hpcmzx9XD0hurG7S5inFo
KaEJxJE/q4nZswVfUJ8HdVTXpguwo5RB7MuUEd7zI/drs9gmlLV/GaJIOSlmsTW/
Z/5gmqcn/tkxENOB/7sVLgvaU0cncUtPCAIN/yRiKF2nlzxssqZsl9sctny3Kzxs
74xzjdhEBlu7U9q9/NT/Kmvc/QjY4aBD9WAK7PTrg+/M9xLO4fQRSOFEvyh3XFG9
aQciEnfs89skxaxKOnJ2wXkBQuOgSPa/Q0iFxd8X+T1pxTkKGEhfTYtO/ASBNyJT
k7CEM1B9u0AmLKuEKa1onj8cXG3AnSv7L8p1zDof+sVq5953ucdG+EbDdGrF3MbM
T00U/tTMO+pZalwHJd5pDNTvoRpdXxzrLm4OHslAAGBbciDEOtoDsZg53sGxRGVC
rV05RAng1iy5WUZ6j6N7mZfv/ZIv7P4clJ3c4Tce56wfagpSiJWX6sxk7/av40OD
riciZK/e5VihZAo7gTvkJ1C4BC+n8kfG8Ag6mGzfBcn8agIe7Fc+8Da6arVhIk6o
dXOHpLgSL1jnbVyXRG9nwlb3xUpKRQR/saL/z/VppZ3INUVfv0+xC89qEMszYuPs
vdktXbDQdH2g6UuqjFn+POGUjTLtxiWMfoIzaMTn8BbenilFZQmWyeijbmld+c/W
Z1XqyV+jiu7df0+XfFaOGhd+GOjNAm05qcS0gjDxHuC4Ymg/NovCFM6N7qhR1UDX
cCXiwb+mePUaQUgJCO/HPnUKtoQ+Oy56i9fI0qYR5RnBWWHcEr29JvsR6dCrQBWA
VId+8ljgzjZ+u2cYcOJBIbJdbZzW486xXsZ3HcMBYCc16I1XYGKD4floaLR5bLIo
ypz8HLyDjuZwzuhhkGPW99syR36mlTKF58wiSUW8ngpPAru0Iu4Zy5fDst8G2dez
DwoQfU6ynNGNx/ktvUYcikUiBgemq4cVU0E7ufKw36b0kUfl4RqJWWS0lfl6v2kU
AhehJlz2LmIZQvhC/jv+VY2FCfnx+oPJ2aPwMMvYQjBvJSVS6HHfkgSZ32+YRGov
dV3JIMDMTLFnMkjF0JRcxUkP0b7Ya4xm3tq0+rm2TVmUEK7k1jz5IDy1OtOzmqFY
bG9AnqIuQuNDF1i4b0OkaHl7n8XJqwD4A87m0xySs5i6x4O4UTDUtXnjxRwgUDGv
rRW5SIAxrLfgmlekDBFAy7ZZf+kpqu8hvTtVUhRnCgXLmhDoOAqvDMB5ERvWJ1qo
BVhJuM+i9w/aMNcVeKD1wUQlJle72Ra0fdXAMAlcT1WWALwMjIuG6mN/hScyAx6/
oJFXo7T1zlXMLfFgji7D0OErDZsHYHhr6bB5E6BWx8sPS9DUDcgL2mQlhHU7Angb
dG2ZEFwG32VCNpuEeJrLCnXevAfSJfODiJN0F0gXW4YjsL5hD5YsoiYJlfIxgBrF
F6vyxudxZb8/n1Sy+UnMyNNBvGR4xfaou2TfaSqCYH2TOZ9GtH7IBc5ZuzNcGQqB
DRYiyHTzpfz6cZpbNXYVvQ3KcRWhuxcw/0Ru9XIo4IUg5naDT51GYTsuZPAy3pwY
3JsCYAjakKKIy79o26YAB7IzF1uocyAOEMIONHBAG9NwiWRwhAPxIjChE41pdC7i
0Em9mMVKh23FlMsVzF4TmKsBiM/QcTZQ45YAL5lkofjXl/NpvLJxsg6UiGuc4gtA
shthoRu4W2ItpAsZEArMTiko+qOSK1HfwU6tfIhF1ieFB3t8Zb38sG2ad51X7Noz
Ebps7W+MZGrH6DXlNnQgpuqDXqIub82IlRbsoznqmPG8ZSIp6NZ3IOy0FiSLulfb
NQFsSgf7lIJi2bkSwUx2sSGdD4TC5xAK+OMZpCBp0u4Qci8R2Ucm3CyXk4WRICsP
s6nrmAZdadbmdXzedMAfx8lS//Ze7So1RQbyix4MAsgfGJVp4oVuOLz252+o6dWK
NiA9R1k/hPWNnTg0d9E+kiqnmpYLdoWJ/7TQcYoMb+0QV//JufCNbhmpnsHmkN2z
ISfwCzheDjLEBrVXzXXfwUhoT7adqmjWALqdiTbeoRcf0T3vWRBPnNOJXXzazAv/
XcZakiclWgQxVT3ZD55qSnAAzjzOCL3vaykdJBrp23b9orDTHieNll9cx7t1f0CK
68FRgI6PYbVs2VTxOw1jhFR6HIYfuITdcZA3P4bNzQhXEOW5TQjmJQc4fHYChHQS
8Fj/2l3J5plNDqvqoEJUHbta4Ndz7K92udxYGCC7rNfCxl1KTBWUE0IXcvRE9peH
IGoZ2c4k6/9S62ayerwrl/wBGbpUtC2fathh6o3YQevxsscMDeoC6iZhHB8Be2S1
hQlOI+Sm2LsbrWxrsovHqLiNapPEOmB/Dy0lfI5zRXv2gZJGXHQJscNeuY8a3MOw
bYl3LtKuOoqsEh8Xblg22RGoEFPD+3kFMJOdrVpcoDACkpqLB4ZM+aesFLRcLGEL
QaZD54xpx6qwbhSh92l2pV0t/ELpiOwESxoBcP3VcTQJW6hRDXsfza9G0R7s1l9w
FIg0UWdpbu3LKY7ELa/ps0rZBnp9lInufc+na74744AU1J8MzUfVK1aVEV7JB7bT
NVFcpUP+nbipcbogzr6IijyNAaKax8qPk40jiVNZx5hwk/sBtKJrnqzKC7i520xT
4w9QiKgkdMvYIa3lWja66afTCP2cWDd/dzCVstUgaMvBtWYHjfaacLmfOzq6w7Wn
9SsV1CIPto49urCEyY5yIu9TVWZp/ldf71uvwxbAFIVemNa4Kfp9eoY31tegokH+
d6kw8Xc4cHehZTEWY45NX0lTGlsCETxPIdz452MrJvZwW1fW4fu8oSYO8Z6A+0nE
6lU27P+PBE/X2JGaQM4UEtBF7Pw4tqf72PEVou4nW6h84MmncJ5KMwIiepMOAaJr
GTx9F+Ay23HrHHzj4vlcJ0qOkN4Vxv2YX2LiCHHVO/wijc2BdoxO2xqAgHOdz4bP
9XKyTZ2DMmtTgjRjd45FNjzP8acg75OYR5q2fBF0QJ1f4Lf82DNkhZeyVAE7+lUs
Obpt9p2Zy3KkvaWo9KR7W/a+B3nG/bqIGWGqodMg33qRQo/nVPbSUELIOF3rSxEy
wzIYkgfLvjCmw4o3KhwtYycozn4Y7ysWH26ZhRgCn15bQCNrI1e2DDR3rvkWItuw
YKBCC8JZzb7A5+4v3EwKuRlUuCPwPSnoeImJOKy6kqmB4uEhheY7UsfDmN53wSHv
Mhp1NLEnCq5w5DvTHioBPOdGUwZC19NWAh9IQ5jVIa5DE5L/9wN8Gu0FbA5BG94j
qYBNkxVSQBBnVN5i2ZrsDlzGspxaNkqBGLT8cq49QbfuZI6A/wBgxq1VrM3VnqtP
hVWmrplBz8/sj6xWrRv5898idYE7budR7o2BYxSgg4ocSOjMYzzYtoy9aqgajdHn
QS9CtVlsFFLIW2xS/vINlumLlOcECroKjGiYDaBIn2SrA6HwFfSHBQqX1lYZQPK2
iGUeV7SXyqs/bWKl5jYtdFjuyelVA9Ts4pDt+WlOa4dH+4xrB8TW3WfHJqyFyvrR
2+f0flYCeCSuTnmoCxBGRYyI2Zx4I4dikA9EZH44DQMXcJPhEHOmPhvnUP+O1k2z
fK2ZCeXm3i2Z3Hd1L89edgYV5AnoGw8ZZhH9v9Qxyq07Z57wEB3X4vbNDHX/BFk0
ZdDVi2P0KOzKCtcalIaON+WZHwYyizEl7oOTtDrNtQQNN+b6dUZAdvlK2oi50S+F
6EKhPRPNdKrr0w7nFkAL/7bsFn3rUMRJF4v8Sn3vgAHlyukfifNrhRXpcyL58fZF
CoHbjbcG6a1zuSan3ypwtlW+lyXyjnth/za4cXJqWQ9ShvxypsZcVcSQ1lqJIWfF
PFK7Xi9okAuvcXn0lAhq4OG865FZhkmP81cPQRor1ll6c8sP8OCtL4gy2L75qZoz
ogoFnhYZipevULrlFGtmRO4FsDSqezWon/1Mq8DJtRgh/DJ39xxr+KPjTPwWoV4d
c6mX1uk8IclLhVNnZyTlYE5/4JLIjuW/BD3/d0dDe1K/wCvx8BXGqGD2AcpSWSMN
DV3Ye5gEK2otcv7dp7nUoxjNL81kpCCrhwUldD+asej2rNpWhXh7IUNjMuwq5ePZ
5HVlV3puN7ABkEImHVPgG5Fifc01ObA85jeeX4Q3myFLRzBsHEjtBXijhruqb3vZ
4blJVIwenzzJZdLpEZusny4qB1Ve3tcqameuDVQ87qLo9rpBKpaNZDbkeglfDRtM
lXDvjzyqiaZS6R2iJN9ElvhizeXa/Ol+C/R1NHlEM8+A4/1WFeKS8Dn8NpNSgATi
trgDH/A+xlgGfmz46GQufpmrSZI0yEFCDUblrAA1PwQg6M66FtpXb8Ki1LeexWTb
3nCMokck363Ry7MylGU/oh8duJnHqoYdY/zSpvb8cRX6NiD6jXXEIggshwFbwURz
Lzy0ywSTJSzcLBxG0Q0pl8uV7rxJAs3X0tEwdKk7klBrGZKeaS1vWQ1rSFGJcMyl
kTbH3bbVEibwYEAeR4I8yVPiJJR5IAw7QVGgSwUXnuO10msdCfxDp0UvSQeX0zgA
aCh5a3sTLhjYpNm8pm/UQZ9S5E0NTbqMZxDcwiSxaHWmsxvC+tep90tkCX7Bnaf7
PhArgKzn/PrKUWBsbAhe/klPX3ft+Rk0vKoiIvfLmwjniRqvTeNqaJ6hiF12wrHR
1Go+fjvpjkmfDwty6QTX8J7N1LS5MbBCRs9eikauG4vMXWsGCe+VgStiOSRWDrGV
dvJROSftHU64pcxbuiEQm+gETsAVITunjBtp+Tzg2tO0QpgA0F04zlOaAz6n1m5E
KIeuRdQ5aTshS/B3YLN2LriBZSr7hQVJbR81bicihXY216++zjkJs9onllNCq4Y0
KT4pluxk0fQBDaIxRbelF8CWbdGaIRYjMqSgiaFX6rUEF2Ah1xkOdLFh3Xx9XExl
rWl0ByfMFJblUWM5BUa4GG2Vr/QoobE+DHE4vgO/n/6Ljwi1Kdm9hLpWLDAhSFhs
4pHfeQdXFIknwW+ZoC8lJoLztI2g2wD7amoD0/rqfzXs6bWxgdHRrv5tLTLJyAzT
DNmkeue8j4ERfYbSyoEKCusE1F0lnwAEHddboFVQEIQpkXl5u55pTAqXzSKGjg9e
q/WHWXYSWyYOn22h/MOAkwj1hTpA9Yu+DO+wxG7UTPQKdKVH9Flq4+aDppM3rpZU
fptMDB963DgyT6Ytn+Bewtq6JmqZLhhZ8C0jRumE3ZDm5JG5Hom2Vgkk0ouldS9x
dUWWIbAMFtv8J9OhE6+CHXOkPQUan+WdKLlco6vVpPrv5AFL2Ku9EFbshqR9WjUO
0A8+H25QjXV8bGMjmAvClH6iSbdNcbph3erJlStEGico6biXwSulUezsEp8z2r/M
myd329NORJeYBMHtqrycusBfNWzKwxHSW5alzHjWm3+Fi2Fa4E7zrPGOM1TSBPNn
GLDlz55ibAr6vHjd8QwWCiWY6cPwrtofUw6OYHqgHhKeXJP0ou+Rh+BWYzU/krzM
cmdKG/qfIkXyitaCP96tlYk83dp9tKEKWgTo0bYmoHvvLgmFrfqs4+/liBk1Y6+b
UgeovZx7cSK5nJKjARKlH6mBhppH7BsM1x/BkrqVG1lgXa57YjawXdOzOr/pMH8e
Q4KyckatngMInn390GmTW+neB+3sC6+d2rswaX7sq/azz7eUNdpWLMlJKE9X7uxp
WAKf0bpBemNRR8sALvWuHRDPhOjDKXH8UTUj3nq/TloAF1oz8vewX+oMTZc6urpj
S5UL82ojuHDndswkorhNLYCWDQWRsFW6yLF/tmA7NNXc9BJuFbFaB04nnBeRBNgp
F7w+R+iPNFZhxrjbamRGBdDYFliPz7s34fxYgvtGZHUbSY41Rh99CNv1hlDbCCOT
1nrHOm/2c3qE8O5YsCJ8f1PkzviTMrK5eKG+oKfLqEihMqLktPVRMQFLxPKv79zR
BVGup5CPtjblVxFtekdWNssvcJxYP8mYtLygoWg1CFtdnjLKXqA129PV9nXtTxt0
nuYS3foiJ0540GwM0i2D9v35RxLp8JcAARye2tQmm35JJ04yr5avMhRyZqGhuBNa
qC3ATXe57MYGt/7Q9/s0+u+rkbBpAKIM3vA5ifoErbGLFPt4zdu2kE7UUagb1Qn4
2iq0BFcjqyRSQgMVDmGigI7FYoN0CdrPigNERlYRa/pZAIvCiMOlDQn5scwJ12i6
6NjJRhaKCm8Vrl8/2CSsA8V4vcduv85YjvXJ6tWv8Fy5QKHx9BjeoZseifxXfe9S
hCEegeW8FZXJjTI3O/+1Po2bnMZjqi/geo0H0Aa1UaTXBFqLcGUkIlnfhJxIv2tf
d1JGTvpmYxpi1JIiv4V9ZEFKyQpJewA4tzlkrJQ9P6rShcZgg9DwQKRRzAFXc5Px
qPidjK1HaniTKcgo/WcTVzcO0+hdunKBAJJv4QoEKFBRzp4ZQccszZMLrvzuqYm/
UCS4tVIeWBGVkXfQVNG9/wTKx5QpJXrROCb5tZFQwpBQGRhNkSVIbMeepTIKP0gQ
wYzAioRMZh1OhlmCXRnNyXztGTPi/gvBMkkyQlKKuWGTUq8OItIFjO27eXcYEj4p
U6Plvqj68QqRFUJqKeTb1117wWTYZ8XGI0ImGpjBRLQYS3XqTVff4LhXpLSRee76
55MTgd+wrfLNNYyxUdt9sUkb2mjkvCXDxX0rYnZBfFXf9ih/UIfmLBVcUeckufbK
iPBRNS1eFFkS4asrkeVjQHjg6gj4Q0/bQgEGi7mJuxTQf9wfCqAqTh2xZLdnmZuD
P3A1wBn4Hl5bt917uaNBhPWhflqeKRwvf7DRMRRr63hEZt15hHwE3FUzIzVmkGc9
mmfUPwumfmSoipDxOD/ZdA8Fd07mCQSOEH6l6HnKklDSlI/i2UpNUOBrzk5rIX4Y
/0QjsEzV3udhOu2tt4Zm2aGjmyrU+ccPit5yVoGyd6l1Hb5IGfk1it2+Gnx767zf
/VpgHT/O7m6ZrQSzJSg1X69iJ2KWBnakm8xOlpiFEUWPrvL+0RilfD3viz7sf3Rh
t2a6hIPIW9W8CawZ9SKv37ZgYGe5rkodZcLh4Q4qL40iOZ1Y4BSw042mHzP9v5nN
KpfEK+D99o+uL8fLl/sRv08i/En6HN5ll9uRFtXVkXWnNEOnDWA1ognFenqRy795
z52GYb1Mu+F0/bVgsTBW8nRsL2Tm58w4zOTjF0vwHnVw7axO7PsVEdnVX04BHH9G
sEBVgrVcGKfyktEF9SO0kYcJVaNUd0IcYtbCJtKgOhmhK5ZBNBpYLeSz0VCwBPmD
Iyq1Sj4rhxcvABaBNoqq3392QQk30CnN/BF0icFr/1Zk4iLRMKfyotv2BPSDXJ5h
E18gvNxs76+vAiYaJMTo4255/XJN814nKrnkibsq+bHatuuMVBAvRSwZnKKYCgDR
54Lddu3/B0nMO3YpIeTjrjEEfpTnfSBxee6K6dW5k99+et2eteClDbEVt9DkfS8M
t9mNThjDqkapGPPSoa+eqP23ZGA09trIdpWHKhHXiMXGGkLk614LnqkeBLwqYWr9
2RUYADTDS+gnH7KbK5C/bqFJFrWLd0VFZ6n+U2r4QJXgEe+M70zQVCoqTQ8Cqsvv
54+6Gcv9oc0H79mNX9W7n0xiHncWAnXL4JQXLd6tzXwkL3xHxp/I9VtV9KgZez0p
PdtNh19aaf7yce7UI8iG0sFMfuZNFjwC/fpc2KhRyqFSQgZTbyt2FtRij4tCdKsQ
j9vRwBYzchoKJJFTjy+ZUtt3WpiZXxP9gsOQV0XQKf3VkxmvSMqua0DoD6NJrNKB
67KTakSCW+O9chRvtcsSiGckCPvW08E6c8BkdmDiRRuJxA9UY+qYXiWDYAciLfjz
5pakO9iVppdWHKvglFWRQIrSLD1NegaDIx7PtUw2VJ8d7d+9G9yIOKdPGHP6yNME
lSV7viKVEvszT7WOOYgz6poyl35TpI2VU4iTyJmZFJCdA9LyelR/X8A+EMXpcL65
7KdqTDg/L+0hLrmdqeodW93h+4C5dKkCSyJpjgPhXTXw+acmIk0zx8mQclQl3bK7
+FzJEEkoB9KEUBudZ+/eBpdOUMg38Bcsj9NcJdghrBcSlny87WGb9d8aCHzLGXYm
uLG7ZLzEBtrJBANPvBzauF3rqlU1d/5IaccMALwh0ovFqMP228txgUCjkUY+I9TN
WZRVOW4Z+XgAODPRyqIqO/Ltg8XNdW2yz4ulveHYl10ZQYqwiB5oTehdtcY3Aj9D
RHnF+HPubaLN73ujk4kMKvaPhSgXrmKzLCx2LDjaqUz5AbUHwwjZqJH4AKrx9mQt
zL+TpXffjP7XcIaL/TutxZCQjEYD0n0JpGNz0BwEid3BctUAHkSOM04PP/45AF/q
wK+JaHfgQDTmG3ao9JaUVYqJstyVpNoGMnTcxB08CW2u0odTlq59iohBcOSBgPPA
rgeWRhTYnW3CbMsKhgzN1bmUxouQQgSNKDpZLqbgg1u6qHulc7P0db1KE4Md77eq
j3sa6GOv1vhl6y24ZKTr1rhDxB25Q8bpKt5qumauoWijeh+1wIN6N5EhWBnqnEbB
C8lri0sDHqbnEN8CtnX1IHxjbMcHPg0uQTz/fuUIsRi5+MLQvTM+zL0w3qqolzL1
OFNJNQOsqCddo6dDVdYx9K3K2HJe9XNT0N14qm8Zusw3dS0D1vzRTfStBcGllXkO
uJC6teSixGprgv6pixwQV5VayseiQF3zgALdVQ/A/7qkYeObrHIQ8BlYo9nWLEhv
lyaL+aiZc1F6bGHzL436+E538GHp3i2gboikFGFEu+PfP6AuQjeANQY39n9CS9xj
Jxp6LkAQljabCeNHMVJjXD6tRmX0oOriUVicsq409ELHK3ryXfOHSaHjjywVZb9k
u9mq1xnJY716XxGRRbpYNflsVGc35pdTSHisVX5erDnhLPDjNJ9JFeGzYhYlB00t
bWHNCuk28SFIFfUOBFeexBoHMfbP4FBzC1h6nF2vyUqQDIHIQJaNm+Mx+vNJpqCI
G1mQ5Fru85FCbYBRtaNdk1M9HC8QzdW5UPBUR5Kn3uKfMvI5xlFMN0BSBSOvpkKI
hd68zGUVuHpQOZnSGOZSPlRSRFkurSYvv7Fqi122JpfPa21m/VhOdp40j6Q8dbBd
Tk53rI0/yeE3p1kt4WoMhZ4kn9xZ9StzDE87yalK9UYZ5z58bBOR3K9S/LCEVIH+
KM1LfXy1UvJZ4EZJka9mllVVTR1QaoCpZUfSSYR8HJ61pSqcvRadVc50bHfnnWto
PORCzLaqEhJOwweeRouseTt3aZVC2ZUyf2yEbjoxTagysuqisfWwl+GpSlWQHFAa
JvP9Iwp8Fdri68AnFRXF9tBli3fwzcJqDKfpMi+xHydTMa19MLvbUGpUBqW8Dw/C
60Oj02CONtBz4wCC+VkmGw==
`pragma protect end_protected
