// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b9a8jWjY4Fn4VZ7UFC4kWzJ8eZs7GaOM2Dpgy48y4kpaP3X3wAUDwXHI8IV4wMgx
6PPdg2z1qZl+hLyw+5WIj3jNCY6zMjAjXhn/nm2BsEPNdlDIo0pGBHPnHrTZqSyd
uozxgitQLwLfWap0BZrkXP6kSpiMoQ+5M5Lq2JHBu3A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7536)
PoZyYa9YdtmIpD5PltzLRAaxKoI4EX1D085WPAMAnQEWMduQaGia8TzKay+nLu44
v1VNVdSSJ3mG6V9ED6HEWudkzn8OCkl5QHO7lczQeV1YeIgP6OERLvarYVf7iQtU
JiP0rJHhF7+lagj9xX6n5vgZ/bYTPvgVDK6CJDoiQe2VXdOSMAjkDDMC0uIwx2o/
BVXWbI9ni5SVHQ6xg1RET/rCL0226Slt7KEd73Cp51mppm9U5XXW0acpehv1p+FE
G/Z2aFHstoWuUBpyG4GXFwAjnDjthYfXVueNAMhdsdTvrSWkFGtr10gQ7vcFI975
wfiGbc4t+0NuW5i8YGjHj4pQ/3gA5yEw5o5StkIujyq3CNkYKhM59Nkf0X2zgnOC
YbPiiL4wIPnLIcQeGRe/J5LSgBkMgr4DkixfBScCJLQWFVpjh3pLWW3Pn9rHG/fJ
MrdA4MNEbHhyMC/n2XutdEXUUL5L+DgnduBuMlvMncIkf10kAPiPT3RgLpDKjDX5
3fNwpeOJFOHMGCRW0MUkFY/xokJiv7J0UkDw6hq6eGMftkkQqtSB9h7GM2hX/DCw
BF/MoHyOrjttV+tr+fiLHBwHKKe0zUUwXFbQcUFePrDymWZyOycbVETPBGwsihAQ
CBpCqZqlNqQa0wXMXOJTVVzuKQwu2Pbbnoq3ywyssKgsZoXav+NJiEB0Bqvk6CZZ
t78MvcgU8IhI7XRYaj6Npvmxn2NFigCRMs35xP5fIVUi11UTCejVsvDYh+zYhRm9
ZIkXtv+Hk/XWSwtcO07uOIBq/8vSE+F0mGrm27qHeGRCi2ot9UBJFPLm63I9iLXH
jmzG8SyJVWM8zd2JsXR8JeOdTyuK6P6hXG66e7MGKWOrJs9LuevgnClS9ovkIJG5
n1W3t1cJ/AAKeyg9XX+SMzUD7k7TJyK7hT3xA1Fa+DjV37eIt32ZO/nXFtIW05rZ
cJqcm6jLqt7Wqx73pLidbC6Mk2bKJcdBjMgSKC9S8l8AjJPcCsTPtO5Fs88u+Snb
Jd7LMq5a6aHVGBFK1ZmxRaFtCo5REUAXR/X9H1awE5wZ7nxdKjwJkMxhISy3cs3Z
litiqz/+iKkTH/PdF3KGIfuI0EzVWlqaaMKNshCjrRcwOPJbMAQ0bVYQDXbxMjzf
zeztqDAOgT6hHqdMAzAZgfWhPUM/UDtZ5wUVZuVMTMlG0eDycQSbXf+mJVMulOPc
ij8x+GuAkzGSoS5l8rHsLKkSrAtas8yUAJXCYHxu2jPfGTbuWweh9++Ye59Zxg31
/VhRjvmyzkCL25BCLBMefxvwMSxWr6PCpZq/RT8Gsv1o/GVEhWtIxCBbyDe3KgZU
HF+9A0rZS1Vw0qcqaRjtfdWEe8VOPkCwQif6qzCzYkb+qbOBHD0mvnHcottvo9eR
W3QWsqGziuZXtHfVoJf+cOO9USVsm/+kUgbqcrqSWSG8lMftcJB7KgRQ6RFKABVt
qAxbF+TFd9K0xNyzwJc2IppVTclns6Y7PNd8xLsnpAQGMnQ5WH/1sTJa9PGOJkA2
sTUzA3Crna0ZGnFE45m8UsF5LNJbnd2mTlwDS0vdRaB/SX7T5UH8yzeTUm2QhwtB
yeWqpn+Xm9PagqHFrpv1/N6ssgHm6oR5UFEEsIDdi3Ud5C/iswS6+GDB81+xCT7f
8idQYY2tKQtvxaAyQvXS6jicu4Q6WR9XN9sFzVK0NwgkS7HlqeHqwoCSPewJ5J+g
XEABrOdmqF6hyFyxsUeRpNjokW+v5foY3bQvFVOdpxMiyDpYYyEQvYhBnlKy3wfw
Ze4J2nBN5j2fDIdlt/EEhtWIiGDLwSXwnje1BixcUBKjXb+mvuxl3S3kn+0mbUgF
6V1+lZq7OTeW8XqZxOwAcxMN8kZPdBRnr1lxkerhgeEac5bFuwijlf0721PpTBzI
hLezD3+PbLM98k+z3oG3Y8RpmxvlClJXQYzH0qdf7io1itTTZevGAP4f86Fl/dXm
G5+JAffb6Tm6NVxY7aL1iHL6BCgackBQqNrM5WvrbY+JhsaPtDNuecOHXlsNqz4h
i7K9k6csI9Uy0gqtsKsLjLeuI1xtHTclHsSN79QpsppQHWt77RTYlqkdKmf/9X/r
w1sDQ4gbDva8/IUayFiWbBs1tXn9yZzFDDC/e3aYcuzHCMEcmes6xTmaskqbOSMV
Gw7yRDR3lp0bcoigAMzEJsLJyip5tjoxWtwPypE/LrBO3dlj0UPR3QxtBZkT48pg
maAuDmp9emnbeH79ow4HH0OSzoQLsRC6It7fxVnvRF0yePajVJ8VNqCOYDBER0jf
1+GMdAJ6lQf1uFIaU8tcz4xd2G4ZSR9SUeke2ZqtE5uZdtkiDqYpE2BW8YGVgtQ8
MqCLdTfupmYVX7F2o/N7jBsuiLSVGLjMbge+uqj0NQp7ICUdWIptZ8Yo3aMXLJEX
U85IHYVN7vl+ek6n0mtGaP3+wXSd2KFsDBJtsGHXZcG6ftOdWnIQ6lt3DuZOPgUl
0H72gvpfAXzLQk3RjQ8oRnel09DzTdNXLuSIzeGucBitaHq1ltzLUBt428jfg8Lw
L7HPIKh1vSa7z4yDNQUfuwLWu3FRs3tITjRYWk+maYd+TySopqkgeZOPtu2MKb12
gHWrJu2wgUbu4IYaaDqR32SkF4YFKfFd2rpuN/zAiJMn/1ep4pihFhalceg8PDUQ
AHNTjfvnVtP/DVBXh0vkULusBbGvHkNsg3jdBaN3k1EeZy469xvpGQhd3VM2lnH8
h6oTxBhPHCC8pxV+Vdfo7cWRUF3H4stwqEL57mNkagYcbBM6pdETvLxa0uC3/mg2
WLBjTbvwNUstJb6dPyt5pbRnKgM1K8NRTv9uiOwqmdPNi2dlbIiKbSQQPE7TkMVr
ahl72lpS9vQqvqzXvvA/wqekzdaxOo1yuQgRWS/1z9lpFLHvvzTQeNzXtrx8T9H4
P+C8i87yOp46SC9mfNUf7jzcYgU1outeBXgy93XS230HXknUSuicqDsVvqi+ya1i
X90QHy/z3vrN0vLXZasmmOQEuo3CYaKZMhP6pnYhDpT9bUU8kU47KyIvAL6iwqRE
V52O3qP1xTBuTO3hFa2w5Vxm3ozVHGjLBN3FSt34PfdSxgyuo/nC2cH+Zixhf3qw
wqIaiZHczn5ohUDCC6NjNC+cGIp4wQvmRBf4R9q18y5Sv7vJaAC84Nntcm9oaGYe
EUOF5gdjIzALudzEVyDQ+kRa1Uv6/ZBtrSXWdV6SNi2HdO7eJY32Rl+zuhOBsK9o
5EKrWVMrVQdjP1sjj81cFLtXgeR1R2U+fFptmV42HrfMD7ZeNmfnxsRwkjRzj6XC
WF5/l9Ic5CENqNeVk0B4tuVvCw+HL3NcZOuEKMZNEOwmtwbzTvPJew9VLMbtBWrV
dKfxYEaKNIwmQua69RxjS5RTIQTynLBkzeAGsHccAaiCh6zqViKSZ86m1EspjwVL
jHiT7B6sjf49W99mnpojBwEPjUixhHIl0wzY8/3dStt2knc5UV0xb8tK5KhudOwa
s6xiiE+SV2BJx53+TUNPq5lgH99oifxFmYxtNdci/7kcW+8anXydZeI4uWDXbuC1
fsprxKefVlTY8Vb7ueg1yYsdA0S6IiTx+9fVltAezYpJTQaftkY3TvJYCWvqFj+/
YmW3K7SFSfRvqQguNW/u1ONIF9BolsKcqBHYyjxvOEb2DaMST0272LSfI/PLFcG7
U+Neb5FLvp81H3iR8tQD7JyraaUVjRQxDVKA8nWXjeQoXGLho7Dfne4uSXuoQ1m7
wypECPeZsQSgip2/68IW99QqW1gUuTlfT7ZSK1bdMpS8gDFBmKO75mI/Kq6KjmUZ
g0c6jSCXkhUVCZgM9oCukkwYLiC/FQ6XPPV2LmU4Fi+zYF2PD97BtAiktPBrN2tk
apLP6ZlCL+BbQrOpLczNfmxXxBqNSWEYX4JpsulQqcoS5ZkdUtjclnZQ3gncIA70
MHshfVLw/BulHeLd6W4PQ+eFibdaxcUZa5/2MeiwiN5LMWL352vRyB30/8l23Pd4
Ozg/0soY1usAL1IU8d9RQGcq0E+9CNuYVJiRmaf0jaB54SX6Or72E8K6l2niwzrJ
fQi7EyugyB+ddE7QZQkeCb55zIHJKAgmEJDl4URQE+R5wXqKfiBISPv4hdCHb5YW
CI+Mjto+wDb+GZZ/QUY1YVYT0DbgVmT4ydBMTdyBvE78JtfvhRvp8nWizpyIemEc
JdYx9qjq52iRWp/lBo3QAXH4bAQfPHL8gzR6j6c/bURTsFOXpfdsLeSnJo4JfbaB
jVdU/MfLMpengCzNAqA/Nudt5TVDCuCZhwu27+KK5DWRZDEY8BWvMX6Fo2G9xQmJ
GCiPjLvn6YYS9IwjudUU5dH06eSxXhcNBhnLsloq1AnVJE1C9MKskeJ7ahkNOpew
oOjMc7RSZPSOd2sgtYBRzKbndWOrEVce8J1QRLo5ar1A+sZp6LjCVQRDieZgiBz0
KL6rpgVxBIbNbKcIHn9gouxBPwqzdrGSnXFz05fd+LLuFPYvnLJAnCSAcnkstj80
s61ZIcrWAoWpXBenOnAe6+DUjtiEPPmizBZWAiFZmtQr1DnWXEFYBoxVxQcFki1G
8YkgkvYphOBjZiw4JAHv+pP0MS/QUIiJNrc1b4I3O6plVEr6dkvqjFQtszgnPp1V
OXBCPe6yh14rjo86r1HNseDgQZixwv66mX7LNlhbhVWR41u1X04sIOVuTM2xyPFg
E++nlbiFQPZV4KVxyt80q0R9mbd5SxvrLGOdB7KVHyRn3sbaYXunnCn0YOv6iE13
tJ6Ka8RVkkrNFbaL2w5PhihI4w9mUBlh35BvJSfrsJ66cIUmPgqxODDx0ZL02lck
GwY4SM5sR8T8SR1JrCfHNbsZNZ5ueOPItZJ03IMmCV5XUM2SReKTAdZhHfC5K2vV
ZqD7r8GWiRvNvqrAiWy7aEPdRKRO3VtmEDfj1LJeKaiSxIgv4zDbPcZU/Hj1Ez2Q
wcvkTsCkcEHgV3NNUN77I5abSaMpGQjIyvuOhn8ATkwlobCo/EoJsRAHDM97ECYo
AgtX8EV3AWsR+wcJv6QXv0xkeAkkoVHxOJe/UrcTTfRSmy8+dyNnLxTIIEF0/fDv
RMc1mRa1kQcFgWKfyA5QNOvLJUc29f+3JUUWIQiohmWIuLTMWJe69pp1m8ocdolP
jlsLbKg2d47X/bJgVqorZrQ/THs/BR3rcHDaZ7LmR1QuRBR4c1Ajkf7Z531BwukO
iuY7Jy4ntJ3fJeck7cnbXeWJPb2nrofeSYWKykjBoV7k23jhq27I3ug6q/8/EwdG
1bZsj+xxE7RrG05BHFClXG7Ckg9Ehdtsqx2OqBu9JTba52k6o4AR16J/pahwTowK
6wU536ENbNdbm1Lx+QU/exW3HHx2KUlP8r3IKJHuBABiB805pxFt1NWkFiEF3+6W
RGqZW5SEu3zggsVg7mMfaEbeXOswdfpqJU4RjRYNlxKBHmf3FKUaVodUu+5946Qc
rSwzmLsahSi6reHvZkwDFnGSTvICo/KIMI4iKw2fZ1e+M9Cl/Z4UN9H7RvPYNZlE
F57gttmADz+scOn5vObtiuIQ+QAS39fxyvE9FKgu88jt9w6VkzyzYKc511UU2hPN
fOurNvZ/ybgbZcyrI5TJ0m9LUuL+wVKbLiJs916glXcLMOuGWv1vZPqKUenwNAsb
lvXhIIZDa5HiW0GLU0fwmZ99k0sHTM2eBTSlc44JNye8+gkCERq/RlGawlk5qyof
QGGCl3BunSRnuu5Xn3uywtdfS0gNLvhY0kP7YHcYvJSggbd8Tl/r+9/tmY1D6Rox
PiYFpSQA/sMHeXG/ayR1bONWRpsPcdKUAB5Asfp9t7tIR51ovPnByAJGhdVudnfa
IBovIYiBFNYxakLbz2xBXvZWjd5d+ugichrvRBHmiEO/u++jB2FWkNJRg7kxvnLz
vwg15t6OJbBoA6DSPuEyxWr/Cj3m6oDMTirKvJ+e++G5Jz3e26StfjGzchzdS42v
/EoGfkQLBkdaJbFlc4ywd5aM540WlIuJbcHyULIFlTgvnKTPBx5Fx2I05dlgfoLg
540mT82nIPSFcktOI4UoY0zjG82eiZ364TamHqJt073ecQhcABOE3q+qXMyllzAy
lrpqtt7+6TUgtTdeWXK6uQrh7wTqeLo4Q1ntruNgDSi1m6UTRgPCnm5hROnPjjUx
1JSHOeX5aytQyVIv3wVLsxnanYCGqqrLSihbK+pew26Gku3sdbSZFqV6hsk9WP8c
vxLs0Lo7KTDJSN69ND1NuFrDhelsJgF9Kw/Si+STE61tfrC4CGfKfTnq9Fh2b1UJ
LFu+MivWUBVifMkEBjtm9y64hXTL1NEGj0fw2p2Nd/CcZv1gQFddC1zRHqCi2WiB
IdRcQiPxpF9NcsqL3/NfQ6Ht5HAnUyFRFSqW5+8mNeIKLBbzGmVKxDqNpberc5Z5
7antZeWjVNCLJWCOuKUrTyJq716HHFWR3ApFpv0gx+xVSFStZOBcmM8ibGeEzlvb
UpaNBn6bWVd6m5H7O7HgbXa/IeFP0iJjne1YGKYI6TnqmBtGfbxZXptZnTf7blZW
9OFQW4Rt82NvdQfqBHLuayt5cecEE8duqA5H44xtxKGwgK1+qUxLAK72KADs3pFD
XHv1pNIzelUj6CYTdESoD35eWqZ7bKeEFjrKXeLchRcoU3q1PDddafsaIknYYJyR
0GLD3wcDM3ESQygvgqAKV8+yr3pDG5+GbfoqL7YJEA8Fcpzu866u0qq2VICZU/1j
0p2t2QChq85doOtsYajS8Ob9Ml4Jc3MN2qtjm/nUCTwWbnRg6YhTANQvaU2WfC38
+WDCt6lqoQeJ2VugdEPhobHf4qucrUMM7viNRDkc4kQVnc0kYraKEWnF7Mdunm8d
rgbo53+y2AWGMaAa6XDitcgt6a47/qlxlInMw87M8mx59IbZuEV3XGTfYui9tLMP
lK18Za/GkQ8sWgcyeYYOn8hUenVjUTZua/7W2Gyz3OGjbePVEZlFfpRIkq+W2IP2
dNwwB/kN8cGVRNcfpCRXzgEy7U7HOefgzbnC8LF/8rehuC5zLFzza12rGVaBjnfB
PQnRiYWApd6k1gAIfr86SxpnTGVzTmsJBJFp0LgI5Udl7ToTFMlRFIa8Pq2HCaKK
ounfkEqMtXWk6RvIDK58FDS/jUJkOGjdPHtJGuOr7nCQ+Stj69itFjqv8GCSuRTo
FaVstvagxHxQGNXi9cQponPLReybD4J3BZQ0jy/Yv6ahfI5a3Y+aB+SJWflaOeh1
jHowTAhObtMCOAK+D7pRIybZAdRKRbjX0XcqWr9f10XdhKdw08Jpsh7mEklr0SBy
bcnlbyDkaoD0fRdi3E/5VfzVncTgGTbPjaQKuQ3/ij4kSwCblpKPpVxn9WjRWcWL
CkmMdMPYpOX7QYlywP5Y62KK8FVZKemR918tdgj/maBcwXm5+UfoWSfNw/dLT0P/
yZfphbAuiK7jWoa8YMXjDOx36KLc35ovyFos3JQMscVyUYcjs/GTWTMxqXmaeTV5
1CAp7SLzIQAfs2+VuPdp5mAFNNSozlxa3CTsT54K1ERnHq9fBF9OSNxAt6kM34ly
YC+nhOKF3b/xc4GMc7uDWvOAgHjHMuAvFvs6Y5sTDmuCS0p3wCzBRreH7+8PBb+/
i0bs/RfQmzGrBwzAbxqdhDei+nDbFA8JCxWSoey69r5AnDLXRm1zejFyu9N/3x/K
zM0bL88ZgKQLMm8iDXVOqOOpDExtPFsMzbQH9yoeSJu3yhpxq4SKico1R2Vnunkw
XPpi53ZiMO6/IBI2duaT2ihmFHgxv/BLpbVSr/3fqOA1fBgNZ+UzzM41pcQx0Vce
j4uDPILeGamA/y3vS3iE6JxHyet/cGQXdsJ0wxaYsjQ9B0YdkGDZEgL0m8hfwTGe
JfQFSf6WMglcaoI+pkLD7llaSqjCkW73+/lJCng5eX3E//hDwyIxO3oiCIeJR1GA
WjSyg3Zpd+LBkGfSJDOJpM8q9ZilflwYa9ljKpor+IPoEPj0U6idP66zDdDH2vO3
ctrDQc0MEKOCihXkvfz/6HXbVfNeomti9/RWXSmX1/0rKxq+B75KEwwvhf7b5gdN
h9mEjsW24XTLUMnxpZEh0q20kA9kIOvFY9K+Vp/kb+ABMJq1QeIUeQt2Oe+sKLJP
e9HMCKrmu31ByRP4txhQWKDYZ6IHK4MQ9n2LaSAheSows4bX8YDFODyvQGIvme/M
0FIgqtxzZSGmwtWYfMnS7rMby0GG+DbVHmH2cMRYRtSHV+3SlIVj27pmzid93Ijy
gBInTVBHbzVIQBT/BaTHQmwyxBO9pmLnG4LdUe8mZBxu+Q1KJBHcuCH6BrXNRy7v
R5qX3spg+ETxgeLLAMHZwsZ4bZaLG7BPDdO/ddGb0ozwtzpQuxrFP9NDep9EhCwO
7JYS0ljx1sX1o87TLhLiAjqe3MyBTwXkaLzbBSZSSbHXywK/7zqW+2uLU/ezz0oa
ocTTDtXbYQ1G8POVevLCP72CvYijZeLLpZSjWVZU4hOplzvP2LLyrgUkoy90HwRJ
DzldOQT//fwVV4RELE543oSuSOLbETc3iJqBKV8Xa+V5NRGitZNAM2DOfwRqT4kz
v1qeaI3B/AnMvs8cgdleswUkpzI7kiyrBk8xwLkwPguHTV6ruc4CuVYCTUV9g7Jz
FSAzet9EgwuSRQLVxLSJt3dYWfRGO6nbPHTnn65jMWLEz6RQTjgswGshrU1kz8dU
1+4DGUtbg6gMGmHAJ/oTtggn8QgQvEUL/WukRifSH3NxO315/Jxbzbqgx1asUXAH
OOrupVR1SvV6/+WBo6Pf9rA03s7Z1lS40vwsj4zepeC2uPOHWF7nNOVpXV/fXCnr
nldT/ZqHv5k2x/1+wDxKMmfBQhmHI2gVjqsRGtYaJBdo6HubL7PjvefMIBnAXwPZ
fW7Aw45ubkf7AIpbCopgWEQNqJpy2xrwy2xLWzQIDJqUXcQz598KRfUq3tSV0zzv
c1BIchMVLSsA/8TPvU5lGFxbZp78h5gMUzHzaRMpFbctMMdF47nquLvQER01H0ey
NJKfYMTlqpvUhMMjqdO5jcgdT0MMT4NapgOvOxe/Hi/2LuCjjgagGn8e6zdqHTbe
vYor98FBkdRH1KUA5n/TurDcBzpxZ7vJzyroPc2Uy2uxEEawDKr3T/W1z4WqeHhD
9qshBcPkbMuP51j9g+yDzQE3x1/X3lcVNyDVhgaVw4ujWNBhZjkMltgkVvp709zn
1Zxs8UHVDEB06YRU0UlWzsY1iGIu0i44pn/Ygql98FCPRH0IS7K761LsZELx17qb
wiHt/92TXbsx/OlAzZZjVqlwGp9t7dVxX8wTIbbzM6on6286TPYrLWcr9iwIRf3D
G3EVtUYVdnK/ZP7vEHeeDSJWY2apWuiHUzG1cR96d5M0pnAHKoh2rxzXxLGfgG9U
2EV5H34HaLb7C/cbuA/ku2AiMl7LRIeGLfNi4IUihBkyKBwpJyBNDhTt1ZBEWMmY
XyWIwnvgqU/0cYxhEdjNMggL1Z7AZus9Df4Aq9UWgzJAWm5COy8wc7WndWJIoRxP
EOdFCpbA9CaJXH8G1MdjqpVEmcyvQlUb7GeYvGBQtxNv7wcmALkciBlGURr/esWh
gblwvbZPv6zkS10J0txqg9kqR6sx8JGdoVj3gPf9qihlX5fMZB/n0GCzIUXvUSMQ
aETkwocz+nU6rciNTJhXBcub8DkcPy02tsAQLNxSAOvPBhSh1/WW0ggsZFHsQyHn
BU2XPeY5i29192RxWV0+3uZ0d8Mu4B0LCqsAN+Azmxj8D27tXpfC6+d4gS8n5LnY
Tuo3OPdyZxFUB91sqb5RzujGWvcozCwAU8l1J3SkwYQ6MvElpFtwtv4iBb8xBI5j
2GfBryKoGuzamw4cy1H4uQ6mfANyPAri2d3quGWVp0BT2dA0fkrO/9OYJnSaHHoD
MYZg4d4nEVrDATMqiUNHrPaD3sPmSHfmJzCsMite+PoP9a2I7xcdoYOxYl/PJ+T1
`pragma protect end_protected
