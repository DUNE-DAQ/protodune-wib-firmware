// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oK0K5jknNTQwVNtfXkapncUMVBWKyU3iDmsYme4RaI9ekCWaZwq1n+mZuLxjVYAB
vV9W3Ku1qaanfBfamRFM776LTM0p0kWr7tbrYuNr/DB3+WxI4Wcqgws2xu0pwAph
mDRBam4lmyQKPzXTxDJ2mcGtEgv8KKXuekRgm7J5gAc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57008)
DAj3MG5RaxUQlln3xGJY7dVMqauwlUYankN1AvbnlHzGerniL1boG8rS37Zd0eps
d+a5mRrTrmnYw/UCshL2MnT3MKDxt3KGS8h+mVJ0FfLkU3bGEFB1LVG6rjg9VLD+
su6+9YvnckSYJHxZ37pjgHC2VLJmCct4yXb1WMAS3rW+KgiakZHLI0Ckmxo6Q9ZY
eTXzJIpPDwqWhKAUNhkZBkgIwTbX5iCN9Xxex1sgYYBomxgtxsGq/2U26VMMo/4o
VQKE+wCyXidCyWP9aG27KKvYxbvdOACq6ysQuY5lEA5mRQ5T4rvXiYBe2/GOhZoS
m9mOp7FNz+AdxALAPxiHO902XUJsrcYQKrfnck/d5rpwM7kiYHd0VkpQJt5SWAKz
bXSmKrS3oW94FZFljcPO4QpnMsTFIs2McS88MEsxXv9nmVP78C4QW1lN6hj39iy6
u9YPwlWLijhrECyii3e+mOpe351s0J+b0UmQr2PYlswLfsyvNbKY+JcJv+5q0xyW
4ia0BXT3nZtwmUYmpFixmW2aA6y6NkxuAf0GC/xWUcuXIt4ecITq+qr4duMLFYAI
SM+wDWOiKu/7grMhv2v6WHHZ4XAxLWGQn7e0TkKEnzAw1md14GoN83FHrAD1kr4Q
jfVUmmzw4lp2EUF41CrYcV8Cdh9IPgKRbGP6q6PF5GKKr30+Ckp3OHcKE+PPB0m0
hc1U+0/Y08797bt6FCS2+n15SOICpH+KMSfXRDm4qEple8oCj/VhZYnVJaWLc57u
C+y5uJlkYncmogPZF6GSrvxQqyDaaHGWN/MSLFuVlys/cGknU0sHcjoWLSrPY7kn
azWExQ3BP7C0P9y0o/UQpBgsYn3MSREkXMKUUQSAICCYUsIkn3kXC5QeEM1pz5Ao
0wVhklNOYFQLAokt2vfKkpWY76yLWScNZzmgToCCww/afU2UsbRVcCQ/t8L74IuD
pDNE1Bvzt1TnZFU4Ud5g0aX7ptyHiw85ZuKoth9c0XY3b0sKHhynTFRAEswoW4N2
aDNAqtyMOy9piWWFh2ZAzhKauBfT2QQ+TDQCbaiFeJMGpy4gCyhFZ4vchyVr4O19
cIGTTOMUsoVqYONgrwYi+uBMhskFr136UAppGOlCos3J7MJKOPUJdF6sCsrOb9ua
q5nhTLIaU4xAKRi/s8Jd31cqgE51gJ9hpCS3CGLOAeBRqxBh9vB2l0TQlXKmRUq+
liWauPwtmSVrNzoT4xCXpnxxiWmgM4cgtZQW59YhdppKVrdmZrJyQHlCOyzsVa0b
ox5CCd7TtKMBgLayQO8aZySwkWk0ocLcyA6ebOrvmoasr1aOymcyvL1yWObB0PoZ
4UiI7owyawvs7z1uYIQoKCoKoJXG9Togp8ms+lVZL5CBV9Xi9/Ui8uOTkA9Ccqtv
f/3BhDIR1KkxK9tuTFgnib6dtPevNisAHQtIY8RTATGPl1JHY/I9y/YbsOsBt4we
wiOie5bdSf5SL4hzELTTqABDh/UDh3VgjZK16mpP5ASLAgyJClOsr44Ed+qeqmC2
icIlMDC6n/IIiW2hbLzHjxh8rS8GGjlhyh5Zz4Bdoq/M1l2ongEoQkhubfzp8hTb
JWh7eAHHdeXw1uwRrGKhrGzHFdVNDkxNuN7yNXPauLa9Mi2PkSHD/18hZ+1JXj7Z
IEZ43vZIV7SRb8OqFnTf/d/QENWasjfKogtOEihPQDbEnGTwKGW95IlKYNazSOMB
YC72E46o2s4twQhaXw84DDxL6LymY+lahCcDNX0IdgDMLfFjEJulk3m56Fwsn8cN
pb9v/w0gNZtnnxDKrE9/AaQS4FWWub84unM8p29jNlZXiL865/Rz2WbzeTO9Fui9
L4G0uLFCCkZRBRu5oAwKVgtSlSyRyzZXhYMc2MF/RuV+yWoDQNu+miv0Xn7TXdNP
JmWhPEtmfQm4kann/V8yd8LgJI3JJJ6qWnbLFIGa76t4DMUacFTszAzyBXbuU5WE
UDnFBngBURvsN//h1Eawpuje5d8jQWdUxAZZm1YZF77oD1103H41TMnjXVAGmlaG
jm+trfc1spbS1ybHqYk2qegQG8w8vchESBAPe1pMfHk9TpK0iw4xOIRwxqGh8FfK
fSMJOnk5yDM3Es3KB7HvInXZtn1j9ecp/Q+Lv78eqKJVleUKj6um5N08v0//tzXN
xIDG40r4iaCdpukrhHHCb3FtX4a8l6HNcuqHalyVFfztQc7J71S5adiA5Qyvde48
rN5WA8lzerYFSc2WMDSKbmZNBnBbumDGqKVoFQe2eg3N2LXzPpOuzdvR3t19UM3i
85yDPcelezy7C7kphq9iGCqpR49nMu94/+pkasqTozyVY0lCoT/nVkwU/9RXD0Qa
mNGxIgLftUzOum7IqMmdVuajhtBoLJMBbqmg7y+8JkD14kNqxDrJbMxO6CS7dDHY
SmgNzcqhPVhBjWigxvumBz/P77b0PiBEqO0dXGTIU67gJ85jW5g/mQEC+MVOYC1n
k5PuNH/xtgt2q6nslSRNgLk6CJxBQOLCb5X/3aeLLfvHAEGSLzJ14Zw1yJvnr2Bf
Gh5i+kvQ1WaypZRmGTuHQ9PQkgJkU+kDbEzw2siZ/4Su/ldnqty7DT6k9SRFKvYn
n2Ws1Ypy5aSXC15Vpk4uxlua2ae7k3nhz7TK0Stzv3OEznfFan84TCJuh1A2PXNw
kryDjL+PHw27gW5hAJ6GtO++6ntypxby+fR6s5HRWwk4H7XlpdvGhykliym91g9S
Twp6R9JUn5K+uNvsvUkFM6lfS0/2d1bAqZv1v2Q0fivE+yAjlgOL702YiuzdtKpN
g1fVtGO8pk4b+khJJc9mmDu6dWbOrJKPM0uLWsGTadX43C/N9LA+QS0bf9wSSit6
qYDr0LOl2BCrk9oaV7dDqjP9oR6njTCmv82DFP+GJ+rU/ao5v4UGNiDQdwC3tw5N
4Tetw4h/j98Mg4Sk7NxtJFSWYri+tjfszqyPf1PWiUVcREH8JCHT4MhzyfxTqH/6
nQMlnrVEXHiCO6H5OGxIaXpOCYqCrVTvt8NZOnDmdSVhbqf2o6lD1KaMJR/V9mAv
eYtEmICYUNGpxPRVrREbeWw1LIPAMRIuMHc6KcCJlQHRHrFtKAxLQzgCrTrGolsS
imC/Ps8QkC/+BvqD8RfEf8ZN6nUm87dyhlarRgR2LV5S+tUSfFl/m+OYdKJRUB2V
T4TKVYGK4WZnlbCYBXThbWdI2WrKuCDCNdtS7F/ZwKCdlA26an9HvDgtbJUPW4wr
pj+JZ31oQ0wLZL8dvef9d0w3sdQJD99e95EzA18oNCZ9ADL1hDaYRD4U8InNZqZ6
H3+0D+nPM6RbJC+ON6+U6hHVD758tLbiQxBfnGbQBUIT2kZnxKpIF3KOUbz8bnjN
PWwblKpsEkN5BVbD9JJOg9f2WldzUjNMkJIa1zUXbLxsxSlLnPGpGw2JNOmONX0E
Kivb22gUzxOnqky7YRdYyC94H/vdBjjYw4Hb5268YB9zP97M2aDtpsTtndXfKZ1O
pq3YFzfYMS8rsT6B9AUtVrB2emmd/nTps9Gyrg1vsIoAy2cn3RZC6dCxZFgnEmUy
fE3/gx8R+XMHIF6vXRxELVqGeo3weX4IKoeh9VB0lcXtR46+6Gg+jvOeiGR3HxfB
4lEwpRZPf1Ih+mOUnTz0cRkMXONXuujsZAISOiNE1oADEFxnVhAMePa06PwgHFOt
a1PQeJZgJUsLGJZ5xf2y/XGMUY71TzZrUP30GgVoEaTj0a5r773mxJurQhYLwPpD
XwwDDICJKcUioTlgJ/t54kbds/FvxaokviElF7JEUXeQlBzSTOjIMeTViSmmxP6Y
gDfxctoYsMkBmt6bSFoIZxNAcpesaU8o2fpnoIX3AzQpI4CfJw4UiwKzSWiWHtkC
zhf8R5HuQJF/Ecoen1YJsdAXA52slEZbf9N+gG3uz4vAlZRehGiiCzfiAK16yipI
+W4xLPJUHN084CGJuckkOr0kE2ssCTbmiUX++zbS+VM9x+9m+dsEz2wjFkP1vJDB
go+PZd6E06Nl3It1xfaqo3dAxWWX7bnGKKHJNYLQcKSAVRnVS27/fkbA0OmhMiRU
CMHgYAqVBa0C5mKViRXMGfe5oa0Ft0j7Zy8vECFZbRnXW1Kw2oxyYvqDoBXc9sOM
umOsdMPZSqCucjmWKdSbgvv3w/k779bjdYvSqJ6qyRw9nKYxBjd4vGwO3AfnuXur
utwGmRFM0d01zOnC41luvfGupWX1Odk9gNUCHKGEDnpRAAMNiIA8Ojv3i0FWth9G
h0PPGwgMz6Gitw25+kpyWBpBh/ahWUD6sTIBMHt0aWuf2soW8609Yj9fDdt6ARo8
g+Dmqwuph5rvKD4PUOnODDnQWgzGQEhxTObzUYED3PmzaG9vP+l7g9oAEEkcVkXD
cUqfPSFrdrxLTT2o2+FNneutw0bEAGDqrWN6l0XVhMUN6AC2q4llSS0CxybRTdws
5K3TY8fHWKdNZYrHQouftwGoEi+936eVV19fohuJD6gCPKaJeSPwDtvlgmyHi5mz
5sLw3dL0a0QCsn/jDgBQM2dM3+OIT1hMBUSdoQMmXupfqqCRuP01JhDEM6V7gK2l
or5Hl6fqN3B4M+oeKFeFQQBCSBAtQqjfhHb1IeX7yji6P7x20a2NQ8S1TqB4PHvw
P/X8ZY1kHTvggqGASg09QJxifxUs0w79Yebyc3ONGdwXuxpqwyEruxfeZoS9JKL+
47mYNiOQICdhhodNkQmEEqmy4A1QVu/E12DXXQyNiGe3RJqg+e2j/iqBg0PIXQng
vjjwkBGY4uR8y/SDtOtaGhWZN2UEKCTU4JG5OpmBF9DKbxPt3Muf3aIfLRCpQCWQ
Qn0moMK7Ed/XtBUyyfn/qF0/QpHSVBf86jhB7bW0BJrTwoKSDSlUIKR3Rv7ViV7K
v3pOyNcTVBIz+ylRD9pswWAqEzk1guf79v8QCoHrhMJUSKODRyoqQXIP6JX7ffHe
Q0wfbSDfdos1LBaJrvtcK5xZaJZXF9Hy9nOT7Q5rT1CSwuXSVp4kmliSLsJ4/KQM
31WnzPkaq1Cwm/yK/5yTX2an1/x61pXw4wy/2pc8d8I1Ftp0f9mZyFniKbga6yqK
JWy84rp1cLlRXY7LgtckD+FjTUTw9K2XpQaSl3IGgdaubDHLMya9HQZGSTZF0YCK
Pz59LF/4IcOQ8iXQ1f/4e8yVkNd5173zsNeT3tPE6zhyDaGiuzW/pFUGcN4oShH+
3t8WTh2IKKRHAlmTDN+hoSTGVJMy3DaIbMtKkeudfgMJbrcoqfjKkaCG4dT3WEh2
G3128GjnTLf2t3YGQkkL3TyB/mWG2Pp5VjjjOE36QbW5XW6PY6RN3ooQkZENfaUO
9h6mSBdK39DLlLM05FPjkqmpw88sHXPQ3paHZqwlKKZsUL9RIsSDml9lrbvjoaYf
eL2qhChdBN9h/HMg2mZCZBtfyPXcWAVJt2VGd7KacrwoAN2SFBhYdZ/MzAeUNB5k
EXywOYbRJ69JN3+cfBSXN63JsJpJRz/t93jhaEiE91FgbC+Rf9S804CbtehNWdYR
B9RKzqUtZTrpszeyrx6LllbnrsAq36flZtW6ynDBGvODUm6ew59yajExI6ZxO4H7
+Y3kfqXntcPqtzzCMp/fvoYBtLmfdiml95yKkZe0pmYZt7uECpsVtjagqlVBxe2T
KJUzmoHj3koG5Gt67bh9sGaDmTlCCFR9gzH+sRTRaeyZGtxlLCRgOQ36bdIUXwiN
iW85sXxyk1Ps6SN7JjhxoucdbON9nWGY0wozxELUilqJXqPBhrlUmZejb/AgM7Ly
+Z8fGxHUjZjhcZK4PB3L5JyKvD2RG7ojk4txMFmbGcMI8krSOwBk6EnbF801YyEx
/7C2y7jObsLD/jps4OIK6vCBspmOhcVHGyvERBg+uduolStLVNJht6hX/iPNCXEQ
4an5o/GadL8x5g4ab2l0Xn5+2fNl7WiYGWqr7rrT8GFF9npmjVrVpM436cJKJrQu
LZUJ5sLWHPkX2Q8bPU2CYVxIiy08JEpTrPhbu+e1WG1CKofCCI95mq+Ki1VWgmgQ
WfBSFKm3aN4WF6DWBa/hFn0WuQx9mvvhogJgJDyd7PHZitGrV1P2XzBousRl7Sx2
O9SPfwsOw7WQsd3FS1Lb3JMIROeqmmUusnIYKJ7pXjySmUHIS1PtniEZ8DTn8wUb
+mmr6FTPS21Mna74cevnq0+pQkRpvlXdGzdXhgD7DeEGXFHADwWk7nkTMLtQaeWk
9HqONOpbts9MLhK2ML3519cxh3pl5q0DafYXA8JhpZnpN12F0TIwDlnVoPrhpo0a
nL6XkNBHrHTyUuPsyMQXhkLjnuguErfrSNJ4E5le097FALH4BMA2J/ztQlOO3FWF
8+Kkp7ieY0yeRX3gNBBvmeC+vim5sWCN0SERntOxDVLlv2wmUKUshtwwZIf8UjfK
NREgfRYIcGurHCpPrXTY9Rg8UEnbyGBirBirsOUgiho7bOwrmUqrbNeU6A34lR+l
T6DqnxxB7IL6rZgF2KF5BNbcwkYR0QnghOtXnUpnMPsE1dkeA/Rj+ELDlUkPzlrb
9fXLfu5Z45H4z4bGN7hAvz8NjfkZ9AAxMyzk1nuPt5Ak2vKj7JVyn9ll1mkmad/M
4wewdUUWPyqtJmOW4AePNhM0hap8D0wEsHRB8S4zhVn4kcrZK1mW5lQPiN7ecf2G
fs6ugI7a+bHK7HobMBa41fGEwrB8/lHOnJbsjgI8Xqnmkgq8pk75aqzbDWLYLvs2
pq1h2/HdJ61yUzgn5vZwDoUDH46dWRFWWoJafAI2fKULMaXn6C7YTqBGMYAZiiTQ
c803Fdukf08m/Qu9QMzTCinqB+WoP+HyUhi8ByW945ylTMf6xBUMb3HK3yER7aI1
eG/WvtreipeFR/7fCymlY8Dya5Fv+ZEqN5IwTpzh9WN6drEwjM4YVobMdbOInB87
w/pmkj68SJ2BTESAxLqFzCPLvbmA9s7uB9opjnmIyN9QTHHdNqgQqYRh2MMV2KaR
Zn8W7lfWt9gcArbDmdr+wmWVFT/C0tesBFo4bHUtWaBzqg9LimgpAgIoGOZRMHG2
tPYSTG3f4LMVoJST77+WH7d7hkSsdnUYKtuZrWrFNZWNnxsRZ6u7hzWifqH2ktUU
88f3Jy90Q0fuNEKE/YEwECwzXoZjFz7DAM6k83914yC1iDZ/O8XnzOqUw4DFPhk4
PzwZqGGAXNL1PNzXhcbl6G9+aiatOb6Dy/kQdjz5aGaM4hjNT5yyjXru5Iqpu/27
ZA7q90UfwQoju8hv86HEaQBLJmP20rMsmAjDbdZ5cQ+rGwyj8O0ZePWa2ksxqh9S
PGD9SDr6eeayuq5BssUiHoNqyAGZSeH0UWqhLwrd0wQpMHOM9/Rn4YGbbtm5kYaC
VZJ8bCDTPBzouctwYkrhY4b+9z6jhHOp65qb8JU5fkR3IpYtb60/gRSpXO23s1zp
NotRa/BDufhSZpesWbXl/tGI8J9sacXpLfFIHME4bATFm1w/14nb8lPqS+jEUJHa
77Q6g5rUMQFOuNoGDV0Ocvt2FQianTy4YHJUSZ2z7PLRO3lAXup7CkHRHvyzQKal
a1UoJ1ZOjy8x8gxz27gr8GgFu2+e+hNNa/CO2xgQewXDHJbBxt2L/ilvMxuOWW6k
xKIlGg3uU0paBM3Mm8MN/55n+94IjrekvhneVSsUP//Xuh+JPymP0NDJ7LBJaXwj
1/wiiVEJs60LFOLXjRnQSmVbFYibrcVyPZm9JLaNNtgTj6mfGz7kadqAisXHObhZ
fk59cs8INmSLzPtT8AaYs4nnvjMgV4Hr+V5QtswAPAzybzQYplKE8ftYGqIdLgUq
zFWSQGCJ7/8PFe6dx4/aX7ace/tRpDE9tyPeyY3DFXoDpjtBrFQzE1697kTzkfOV
wcTbLcZ6TgTtsyiUJXn/HDXjLOO97kUMeC8H18iddgUhn4KtQ2wtS/3vSfmYQgGh
UUfz+ZO+Vz/KDtRrINW8tmG1+DE6QzwfoEStEN7kF1+mDyCVC4FIiPhKvi6ex8lc
rGMuo3SQQhzqiKcVZ/oaDVuHgQayO+fRC7zMipKPpNqmcS3HErJ1pot0CvPknFqP
Qhg1ZEp4ZV2oX54z3a4sXQp0n+tSwaZwUd7PHHZ4GbO1MrY4fJUOxMDr6od0oeXV
58LJGfXadmn1UGCUyzgjOxbLlFDX338Q0Jh15HnQbBoyLDFymaWnsGkdynQ1rUp+
3PC2RJViQ7mmXfo2p7Fg1GkobuZm/l4fL+Tptlu9riBMaJqJ7iXe3kEWNy/Zi8nG
rGfFWdUaCm9DKjXBpAGvQ/tuf1NOF0/g+3TuBqaUGiHIVUjfVzi8sOYIW8qV1avW
Zzn7vY9kezSjlyWEPZYvunQrYQrlAo75sERT0nS7U0IyIABcwB4LMGNyArCP5DCO
49ei9ARDHLTRowvFEpxun6EdcO+/SW5lM8svJgWTODG6MdNRIhtxmhMLAOmEPgAf
r0tu4i8CA5DpL6qeCbWdGxA8m3OqaoOPvq43Nrty2r7DOLyiHTkw0xZRdaJjFm45
gAlTDSOhiisV9alJ5AScOXUlJ0jHYxHBwk+1n0AtSTbttHK9QdGDA9ktTbEw/uFd
ze4XaGV9z0pMVtVt5Hznucl9Zf6y6Z/0viVKv8ZYn4mirif3Q5WWBPIlK8nMnzis
QiZ84+rLrlhD6Ov5faq4jvQmqpsMibRz3juLk3tp8D8w3jIu3XfabOOaKyN+W7NP
YeTo4PCTFwJ+wEsU6rqJg2mW97MU6WPRXgOZ513UmwjtMRjgACVEXROfFHr3znvg
sY4V/dBMdbS1dRHgMktTKBKioxJ4oIV3OTcG5mwPv4Gz9tuHkx8VVvy5LiTslLC1
GsnDRwG5wzLNcwAsJ3llRQHexuuVdtlxzN8EsXqFODqMXeH1Y3R732ewYk+UWD8j
oFeH5TbOJ+v1qstwvcnAjVQONBbg7gEVwoguhOc3qQjlODUoednXa67EiYg9VpvV
Y6l8PpfXcmo4bGOEZi+ewYfFPlvtQYEq4tehyZuILFdCSxE0TeI7ML94ecxgHgIQ
tyqvm3lK7civzjdtrLwP4upTAeMdUvV3WFtyV6E0h9+oJ37tsHKvvCUykH2vMYWe
D1/IPCjpBfJ295OZD2GhnOyAx8LJo/QgKHNTRx7yatlPGQAlCcYuQ714lU7l1En8
wnEDJaYaQVp78uylsZGjnQOi7oLnGQlY4p6TFnESNdM0/I7di4U3lUqdk7hBXXGQ
RsaWAf5w/Y3slTpGSjXJ8YqksKZkxgaeCfEhQUSn54bpYBNOlmNddvB2mD6BnPE0
qD/aFa7zP+ifd2S04+96NOfOHLG6ngdnd8Oyp7ldvDRNM8MkmbDH8TajvKM/ch7H
y3pW/KJaZgKbvMek5VS0Gk9WRK/gSxOaGo8eMSguy50ZoQ+ygAmimPWStsx+qjnv
XFl1haGcu6uFpn45lrHZfdCh+9qHIbXbbPta6q6J3yDaO0lsRO8eFsC8DaYNSyik
4qNouX3P8soYyoXbF13aOpUIOh7IDKAeqwvR+JRPV1jC3y7Q0beF2wQuCNa2BGbX
B+vtObEqXTPEMcpnKh0IhmRPv/eAT7zxDuogs01tp977Go+JRZidiILo5Uxijuir
E8FQ6EoVPkbKEdHyUxIa4n3yyIq2AQEzNDvqOhX2gFr9rQ6eaNSxq0UWK0/lm9oT
ZAm46Tf8xJEdhEU/dX1Ernbt4kfb3tbyhCOAO4ak+FYLUbWK0z9NvraII5Igdt8G
wV9a8EyoA0ivUmmJs8VFWi4H62/eHOhX543W24HJVMZ2isuWegjU67oK8w0gS03b
4K/7zx26MBZmJ6WzXRrn4TNv+DbvJOHutqlxmyR5hLWPpP7jCQFyLuBJAK6r+EIO
0sdq0jax53x8Ts/cS/BrHJ+bE/RG9JgPXRjBZJblpp64Uq1AjXMG7Q1PG/5pu3TY
+pPDpiak21DvqwdbTRjyT8FoGIviEg9ZawpzVVIixsIDOONvSFVII3cLT6Wf/s9b
DxT9p69cEYHI4OUGrp+STXCRbNG86NSG7Gws2pRI79zTXdzFSPcD8WxNo98EWU4s
ce259VcfsfbN8tQzrTyV5fAUiNuXcFtiRh+yLbQx+vf+DSQpRWvjX4ZHAX4toOlT
9r+rkQlXG4E+bqOaaFiRJ1Ap8VPNRghcMQFxv7ZMCzYWAAK7TWQBfjFaOx45hIyH
DXQU5KdLqU1kQJTzB9qIZBd1FWUkTjuGs8s1QLbREgrl2ronAjbAB2+YUOjTArRM
LAES0lJ3HCAi0ZudGs2OgNS1+Qpl24DGaIvW/UBJgrlUgfY3EjY9M6Z7ItknIXjx
Z0n3WnpV//aFRNm0C74Bv7MfxtCMlyxgmJ9cy4iAAQlA2QAHip0w9whXDBtRu/3q
0D1QZzmH/3v6kYqqbngqxTW7Pp5h3fNnUE5Mw79tdW/JFRumUqVPfNVTY+qCcL63
98KSylbzm4lUMi3dYu7hf38CiNHEWfOM3TyFEX5Gd6zLjbw3TwJhEm/I3spXdHmb
inR1z0vvqNlbXF3RoIg1W5Q/GyqR47APW/qOQ4CN37EB6UWqP2adykIveseThLaP
xsycFXEIbfLUtYwCYZlolFFTbikmyUG7s5USOTbHfmgWVzXZ3J+YNpTl+A24yF3S
uU1tW468qVkuMuPpDlKMWYQpsXJnvHtIWER7SxQAEYd+aqUN/JpFEaY/K1qGnz7G
ZYPm8eV0egHFh39f0jt4PESlGaxWiu4TxsWGBJZGuhXBxrlB6EGh4ByiwsfF4lgs
J0H5+O3z61f20uiLtJGZmHWJwEWbVOteBBoHWMDDTHkQBTV9I0stHZ9AjyLi3Lj5
s71drhoghWBp/ZURODUGt0Fq+xEg/jd/38wgpyaXPw5rpngQBULP91Ex9SXeh4Dl
pc8h/EbzxWg1Vy1se41H3PypeH3UFWcM/UJ417Q+7nJcLGiYanEcM+PzR+4ipcuC
e5J+XuBx107d8W2u2AKjQQFRSoeX1/jtmNErELYteJs3rcZpJG/qa5tm9RRCE148
nuVYt7wNrKiybwD6L/PM9iuOgtfrnmKn/d0VwjrOqRVZYPNjNNaqVNRKX/qC4TJN
DrtKeiHqqWmntHM6LlNh9dspIy5acBrHdyZ4nS2Yc/WvmhnsGNcewKAHgUkTwzhN
kzU2ezPlM23VdzMGOZVE5q5RRl4siD2pe6UPzNplLZhLT9cSFumDR9fdSURGUYVj
CrdCH7dB3Dyn2k4EvkqcOFX4yUTH6mkQIvzyDfCUh4Nrp0EVhG4WFDwvW+Dolj/U
XCxDmbJ1tpkzHyzxQrZC4o2WUcFJ9qz7wHwrYo2PDsLUpjw/H0TghGyRDUFju4PF
aj3qWTHO29wZCv7+wRc9xOSSehP3ZxeHGjLQTGvsLVB06lmBa9iPypw4MNBbcdTE
jZmodr6zVoZy/kQOzouIEI0LyOnhK71E/A85hhJNa+ATnHNS8lHcTH6aeiS7GDko
4CQZAhxFLxy4bwkNtD3JzkpquaC3Ti8qCA78bvfwtHdwJqOrYCMneyktxRkhpcYA
LnKueFRJGR9zuzW12l81ueXToeO9a1KxKIK0sISqMIIqFkk0eE4fiZmnOYjJlvxz
GlN4e9WAhck/eenqXZDyRvrdoaV3XCp5pl9+KLmI9OzAjvwLsIT54RSK3dkSGB7O
UQDMOClEkJneLXP/fw3YTtLRGEXOBrAsV7MULC/VucYwlU3SwyWIOnryAYbeeX/G
svh9FS16hCoe6bR3aTfViBO1dO3VEiiy2YHpHm0jKPYAowiw87hfesLDLbA4KkSm
SurYK/d8jTOGJEot+NPINL+oZbl3M+LuVGZWA4nFI8gJKqiQWlbVi4EOUPCF+UQN
iBIvM9EO9G9VFctV60I5KB0sk2sG7laRbihR4jKzL1WH0ojP/6xGJU5PMS+9PvxO
0XKusCtLG+Dpx4dLGXlNdFjvjzK0ODVq9WfJxyYVW7xccSxhmOFgbezyduefeCgZ
S88mr4IvhFH7J3+CUCQrasVMJK0R6SUHPYJp9/wH40V6QuQbrNheiLC2maGVc2Rc
bqlbODW1ofx8GbxixmRZFZgy1k23nF9KP6aOfeRGjsclAx+YZrrk95+7dVPGhtgi
jrA88mB7IoPZkwilqV2pQVcTDHQnhpTL9e0JSVqUku6QYskidjYAzLn6nLx4eApP
BkCB3SpwBb3m6hZ7KkJqI578YlP08RRmqK0Yl/FgqStC9WKTzXJUCaVlmc6aDBZq
ajeIYcIv5KOTxUMLiktAB8gy4VvG7VoRhyERdBiQfWqjOqQfuLXWXPOQ1sdE58pp
HQU/DSvjp3x2U5p854e/iy1+Wymphx6EKcAboxZoy1cKz5zVUGY4MU0nJ2xOsRrK
WlZL7k4xHfX5VS1O6unrHVUr6pCfbbLOUDftQi0O9rG5n0/wyual2dYsWt2brMcv
HKHtJnzPRdXiX5fkiipzHQbX8qpaYLDdS0dD8IjE8sdKglnA1RcG+SUqk9Q9obUE
m+2qSJR1Yk4H8sz4C2PhLSOBiOX0Jc2tnIU4fuAn+xJEKkUygU0T6L7jt+t6YxAq
3l7Gar4MohpGj7W8809KWY3zsLnbF2jz1uXU3wqajAWSf42yyxz/E6N286PqaHQT
a0c+CGbFhZ5JESb7bFZYHersHjhJU1l987ObemYB1WSHjxJxj/M/10M3Au3WPCj/
lgmv6KReSe86cCqX/k9kqcDxAeFFHrnqV5JNNH5pSGqhNSaMCtv5LX00+8/0KhMh
QRjV+KMMpairnaqPD5PxFV1Y82JoscdDSLyd3WggG7rBoaE/UcVBxd+RYGO6R5aL
5AawPhKSNzm9yr3aXDtXlLFoenBO/ao3sPpbol5oEEBhcZHJdpaeJEcRRTmrnrzy
EsspmAgE471xgiUIgx8O//kyFbIp7Wkz5qStxH9nrQnLEJWk0aWsovFwcmdwT6lq
aiz1OUfpMu1xfwL5D80NMxS/Dhdbb2pZBjB90K88c2v/+yl2ZQiw+LxMmeJcVtSm
U7tuQT+3Dg78qRUQE6xMyKzOOAeYLJKAfktZunQoifUiPrgySDtqRyoG4+G7+9SZ
d+Ny23zUDXQgdcY83o1/hOzYPVoviRE4qxb3f90hhnCXptsW6M7ZfvuMZAxdMr0I
HwSxMLR22cAjtsvKcoy1mHdThH78vdphJQ1HWZHjVxkQfWrPGOSWFIOLGWtEVCsX
d6FCEX6FerpzdqIjRPJyEtFMpaXOPWSJHDC3UAwNoftAKyUA7rQM54CaCrrOlvKW
negE0T8yyQpo6aXg+wOiXocjAXasnAQANRzs1y17zqIuwFg1kT9wTtU3GLeXhF5N
o0jv8fBl59uBE6tIOdB6NiqZdPCNlGv5qaFs/XvOu3aMa2lf73JyN+/E0+Ak3KsG
RRDxyiHfNr29GIBaAjQfHmN410H1c3AhA88Dar72TM90LkrK7L01zGyHgTHGtClM
hpKQ3D5h5q5/Xqej8yS9FLoOxhwVyfHPKuzPDpX8hgzWpeP4ArYC9L6gy/7pPdO9
lt5/5X1TvS5P/4pAPEb8NjzaVKUgauQp0122XD+n2o/YwvO/HaWi5QrOy6II3kxG
jcJWoKC/q6I49NgAaOMnOkTAA9PdpkfLMhQ32AbKj+IsK1JlZNOlh3yvmnDYHeBP
T4+IXeHjrt4R7cIGQ6bYU2ViYkdjut/HNLcAbPj5LHOE7jHzF2y26uZE7j69kwxF
AfX/sKWf4ijoYgqPhzCHcdrs3x2iYbabnfsPoLs3WeW1dcY3Ybr4OgkOwCcniOoj
Z/XzE3zLWAyUQK+MLHXC6niWTB7QGt4IzphttQEdiCTsHFthwAm0YDqASFXTyly1
Si/DCwZQztqHeW2GWLOjPPWTw3hKKV/yGLZkvwDobVnwyJfceiERagTIyex2x/yE
QgDGT0AuYyQkyKLn7ti2qa6hrK3f8ibKuDqqq8pVxiBF5IoyAbYmDU6AxHYyPV5a
844rEMGUpAwIFSlo03Z9qG5QvvgiHnnPZ3IXWwFpvf4A85FkNlb1Gfq2syKxHD44
f9UtOwPUKALDi9q2BtQaZMSdnbFjFv9IvmGCHi0vyBIyJ7GrPhJOOr9N5rmmeXLS
6l0nSVc79xpWOH2nbha5oVwzyWMOpD2MyYyBDKnnXVmYwZUwVm36fxofx13sfFQ2
X1ar1DoJwCAMO47M+djG4WUey8r6L7ByJKrO5G8P3m4s67QWfyFFeun4jpbQVpt6
Q9PCwMyEDnAFsQRsWpymLtrO+gLHxrOIfNCDIeJtjdaX1KKNFa5Ofx36gsQpjYc9
sD4dhNpSuyEGhoTzG1Sy9td3lgzaeEzgoeIR+U78VLZz1LNGlpo4HaRtUGZAv1ui
zr0xTqPiIdAHi/eXee+WpwSpplkigYg0nJvgzIUiEFQzG11HWO+zRKpspF9rA5X5
a4YBSkh7Mw2iGtZvGQBVnBhcsQlYH86ZaNpkhGCF1AfNSfrZz86199SO0QfBBNpN
1949TUyKZDhRc+uZzs0P7iDtaVQwFwM3z+/SHj0Zn3gyMH2uM1m7VDJHNhmbhH6k
X29cY4rDEadJFlcBOn171yYPGE65VZSO+nOKxQIcx9spM8Qqku3ZrbqON+IVoEA7
D2Hd7ucpP0m02RupepCZV91nmHj4fBCThtWdd88iODwsQ5RTFuE5QIWQxJ0Oz92a
KYA2nCSYxi01f/RpGY42E99Pxk0FI3vnP/OGdM65J+E3p6e4Hit+WIVUoc/j1BLi
ysaA6WTDMWR7KMwf93gAF44MIWxOCMfjEkZQWNL49YxXFYSWsNXi6Lz0oImBS3mh
JEv2q+vZ1WTAWijgmWvHCXUqYKv/iJcmb6PXql1ZmrYMsCuvQUvT/F/BK0Z8N2up
zpY6qvyqNvMQ9FWQovuQfq+Yr6IYcnHcDQHPZLKU81P37jCaiUt6FDuvWwiUqg4l
OJ+/1mEtVRpRTQykXKahdXxalaSFQQ8cjpc9syaEqkMVno7P9uA4bs03aUMlM2T9
67LAHQxuwkTIsXmSIOTT7wUXcDcEw3fhuf5M4jDJbQuwAm+806GLmP6MUzHYdoeq
m3hkJoYjdrVngKmfP69IH/mmu3z5zYYMRjqb4j3baGG+VIc5sx7BWarkaP5VkapU
Qf3xONK+/e4FMS9GqZ9J2BuHvQpHoolkdUHbGCBC1YrzNYkS2fqYMP5rnWnBjyAm
ta+87SeiaO/caimeF/FdccfP5idvqON+gZ4SflXGYejKqrS4ADOqFWAhRYPeAgdK
7iQ3WRc62oMMq4R6zWhg6MKXf09DljMpGYLfsG+JjrkPL5pHmUSiKsKSqwfnZY20
0Aa/t+7GPHpDmJZxDxrm7CmjJ/CIozWewA37IXBON0h2egcVQ+vSqiz8UeozWpVS
JLwMKHiJynrb4ExP9hydg88nXFH67KfDip/q2A7CmF/Eecz1oovUmCTFg8OD9tLv
RapUPGVaHeShj6wjIfz6vvMXNMcJeZlylDmuqt5f018ERGCJlm6w6urlw3m4z40S
ky9jTjyfvR/5NcrcVUY2HBibInyLARwlb9yE76Gzj35oirZ3suRMDJkjZBIaLue1
9sTsyye0M7JqwLWAKaXbyYa462vP2PxcI3kTHKdEC5ekKG/uVykTwG2maTxX7MCI
FJhI22BnzgBxO8r2Vhx3hcKeX+yZHJOuYPci39bO4A7pW2OeDNKIo/r0TYIkZQUn
rtGoiwa7/adZi9Ezi9JgSjXcmyUtOLoq363PBaCMO1Jvc4DqVD3GCz4q0BYSHtla
LHiB3tQ4/apz7ou9G5aHx6mn0ihmffu58h6Wvf9nUcuRrsaov3tCkexTU5GIzoP+
N7K7o/TLpx12ompdEMeUBfArGF5cUaHz3er93yJ2f/QeJCBHa5MB6sIKXtdPpl0V
4sGe0YCjfnrV2trkPRy5oT32U8/0/ZpGLNTQ+TDn+YQk47HWdmXmVd3kV5rmxCf6
4Vz7G8W2Kunu/ech24JME+ME5cFIsERKJ8K0olg6yzG1pqx6iRK8IF60iDHDQAp/
8pllnDbFIJiZRIvzczKVI5C/oM4lPoDHwktzRIWJgSM3YdDF4naOtxvCt+DVrroI
SHjsXmKAnbeceg4RgTODJv3AZoLWlnV4UoRiW/XB+k7d6RuGS6dqyHVvAt01+vKT
lv9a3GFwAanfg6eRa3PSi5m7D7+vXdDHn0uGHzENxq+pAYMFyvxmGv7eDLouETkP
RhDkPZdMYCz0IyN71e9UgZJR17EsOh4o/TiopRo6OQJjczzKKNr7Ybt7nrwhgbt5
T0LDCpsCbpg4v/CqZ9wjtNy2DHyxMGXa8/jwShgXiriX7rju7LUbiK+gYZA1c05G
M6QcOQsrQ9nI3msV8kab1wjOmpWYCh8SqLrh5F0YrNdfKzvpQ8e+5EIoeAhBS0Wr
n0zK0YX6x1JEMbR6INWzqTEZ+ciLkGs1gpWSRmsjGXu7v8gp9ZzcPnluJC/MLzmF
Pitr3dFWTsuJLXUDh9c450oFXhozAcGBB0k+pfNAtkKDqb0dEXzmJcUEeKVa9Bwl
mcK+EwN2SIzqiiU1qQBO983/+B4CzDnonXDhK2Gnl58D/CMS7d/tDzw1mFcYcTuP
9wwcRUYcxKn6Wn0r0/3TBIXR3iTg2eNPaMgpqmvnA7sN4Bkm4TVInQPXae+//e41
iNmt3/1quGT4Edpbue1RnglX+ib/46iNVYoOnO3EoBmrQuoQPXqVKG84ysnbRGAu
CCvlCrCbDVeX8spyx+Qdt48raW24WoFGpzicm4Ax/t5uv5zsfA8bnLzEht7nQf/z
2wznLo2rUNWg2BZ1apAWIuUM90L397kzPF/VECWccacFv8NO1HROwijoaMiMyGxM
75Rkq3xIbFTn/tfbWgadeAQvC7R0jZgPOengWx3nSlk0Fp5LE7rHf6CDj0JYH0tb
6OjLFdZffU0h+swRcLTHD5WAkwVkT1YHzKM1eFLh3i4/ggamxPGAZiyKZapTLNZ5
bt5WoSL54Oz75XRTzZTEyguwFoQ575zsVsj0Xdvf+UQH81+Q6+ZJEVVR1CIgR2zn
lmn1Pg5D6k1KyWRkiEEObE0Hll5T03m9BNmJs+K9/RYiZyfpAG9j0kLa1ZvmTKPc
lTRLebWFH9G7U4A0pmT64PNjvvjS/rp1k2TgYUwmRhJxXZ8Rvy1xfbz0Y83VlQe4
fDJACSC4pd7x70btCaiZAqorz4BQIFCwNBheNI5EA5pTG0JzWIMrtsOYbT5BCJ0D
QIoOP7YlkwzFaSC5LhubzdH1tOq6dM8P430oAKe0zz+dP9uZAdEXUInn4fzbhks6
vX7LH01013HbJBU7/O/WSsebjfok8jAWYOmVryb7+NdkV1E4dqr9M9/A6Cqd64jP
JQkAmWixK0vYhLskRP7YalPSc/2tDUikbkUh+gN0QLwhNrZ8+xLPQl060m0nJ+n2
xHlzuwQKbBU/Lmfi71CeIO04KMnDsr89FJRXTvxWiT8UgRwkJ6tWX2ontY8SneqD
aP5NFsTMZxyPJD8L+nHr9c57/pklXwcgIbarqzXNyeNIu66hhT7tgooiGbgI9h+o
Vw9CGP9+B2UJyXmrMI9XvL0hxesBFhs6Q0Ltjh86pIwt7bfRrntK+TDpSgEL9EJB
aBDYm7wwREQma2QuzhntbIGubvgIaps6TMgH6Bi+oYKNuXt0aFDomknICQIpI671
cDWCjQyJd8yocPkpVulwsyo6CI8yCm8vCt5OtYyzIabGT+GBDzN+yKFzQu8xf7T0
wtJPVavlYAJsp5UtZntQ59OvKpBjTo1saQHOUFJiyplJveFR9l7kvSFN96N+esSh
RM5JM2rfRl/8hRLbQBCcU/zgV5/KPKvgGXTe2W26/SRDupjuR+5luSKt6PK14iXd
5zDPt1Qjg4Shi+J9sW9iEzexwu6Ik5WtHI/6wDvA0v4NI3sdbuGqD0ieu5GMg4Xl
Q3eYNwoF71BedBiBqI12QOFYeeHbssZzZNeMWWdODWOv7NT4BQ42sRhTW180b5H3
SqTWjSnXeWuA7SsuTxQhEwrrD+jonNdiFSSUY29rXB98QE2Y8eKdEnu8SAaUa8XT
3zo2q1JhJnn3Xx/pQ25KPQbXJM9Qwk4CCqi0JF8Ik6wcTnh2C2xZ33MBQQj4t2dc
nAthuWQQVJ+n1yM7KF6Qx//kbbBBD2BesGd78JhypM5uwAR1WtEi3iO30E/423ta
Wu6xOkWMwrfXZxY7luiNPDYDQqPCmpOy3wcp5BKg7c5W1jIz9StlumZwsZAh3eFN
cXUfYzC4YhfHq5gbEH3jhGgKhgL7kwx0Op6F+wOJ6QMwvkxoNWR0oSZXFpGsbOi7
2HwLmnVrgrDp42d/jKXr6Azh6euh0ItKBPBItu+3WSYfPqz9cU4WCYdDHgWJZtij
6xahjwxTD/pE4cu/fy0XSkqtOU6TsRnCAfefqOnL90VXiLsXjLR773gUEENI/OEZ
s5zILr4uu1H6tP87UY2o83SzB+dkwtIFwWMetNPrzxBhQl2vCBmssbaXmcUAVHAK
cnNiGePDYfbLcC1V6jwMr/K9rY+s1VgQVj2/ZI0KeLPBUNzClPuQ+NuMizG7ao1H
xC5ukYUxJd+0F/lWmiBR9i/Cxn1i5ktjbVr1GqBmJNAbxlNRqMN8w0HS6SS4Fy0p
ipKJS1lPuvBBsKYFyMQidOet6b+rtawt7WL8LFjHXKxLcqIFtqMRpAeOChvHWnH6
AcfgCS9IlZeXxkt+A7UYbZ1jF6HWz7gNg0pi8oE7OTjnIBKhbNf/YS2LnYLZpCrV
XVQPC3wHWF30Dtb/PpwXYjfnL+f99Z2cigdwBT7WvovN6oMIXZ1J3Vl4v4mrL5JD
lrX2e8ADkLHyoDyULowSlV1932uyfb5KuBkK3QhO3FVr/7obaxvuPPNvnehCNO7c
598eB4CRdN2y6X2ORmpln5YoF3VG05NaKpOXhE86lziiPZvGBGF65ahjBC+vdEcV
szieMAaQlmejZIf29GGYpiOQ8ZXUO5b9qsRkUXzCAU+XfNklXZCZqG9+hCfzSJko
3Av7DhQCPh/M3c26A1zK3HAWe4siBiCzWcbvfzSitx3QVQXFqo97rpSQySp19UFQ
gsT9cyYg8+hDGhTQ0bYOnqTDEKURAYQUtKdctPJYDi/QLJNPz/iraIEAPxn6Di4X
L+AgDit731wnt8CaTyg4Afv3MiJTzTMrtqtsOir6hDK6ZI0i2Hba9YuJn3YDiQel
fwJI2lTD1VhT3OvEg40BzW3+gYj4pQ3to7fZtOObyP4EOgWK1qjt1V6zdPjzOCCI
0aWLchOaAUBDrjBtjfRZxZigSJHEitIRgHFbj7pTypUBoARNFXNkFOyN1diJ9uEd
ihjbRTaYenliiaRmFmi8hgNA6fg8LHc2/fEV4z5/FYP34Tp4BqhUvbu+eQICoefO
S7XrEyXEfIXpmvWzC6QQ3HMd3Su0rPw5jRpe4pdYoSzq0Z/9iYrPwWY8kzkc6f58
uhaPvQJZRJuVuqcdZIWmihFOJzJRNQQgoc5s9jtyn7Ph3AUzyvjM1eG0VWWxZE6l
dYoIdVvoaWBXNys+otpEfncfGYmD+bSTZL6YSgkVGRQsn5JUlTsRmJ38exkupfJz
vgqi0rDberv0Js6vgkDEpgTVP41InYhcKTB+c2cBWDbDal+ZD40FWza3DGnLObwc
al6bHGU6G+k2V5pdW6HPQbKRYk19O//faw/JEeZMmg8TvbCCnyFp7qNyi+zXULS9
FI44GrjvSqWD8V2ZwQZQl43MguGd2uVN+GKBmsLtOsh0ovuwuXlWriGIhgKStrfA
849pnZ+zmElNQ4gPCajweqov28GilekoMlI62osUZWz3OxuqPU4Dsr2mvwbvXtxk
n9CkyWmuRKXO8IJ71RuppvbQawe7mMw1ymzlBweFZI+fxUNLFsOvsFJiIxNEIUij
lUhjMPtz3ilCQmU0PF9PolHMQtvLTtcEj/Q2GJrX4b363D6h8kczT9fwToI052+4
IiIUDVjdRUeN+KQVtjGDpSRVpzvUGNP704bJuanGsGKpCZO0OVy2ac/JssjTRRO+
RJF7RF8D6z1Jd407Tw4YPaXLTUP22xZkdNrpmrrFuuO0+Gia01C2oxGteYLL8s8W
Ix2noS5F66BId0vbOJ5uCM7MXUZwX8ZAatCABQEYaC4k8ZxnJzE0Uy5fp1UpdIuC
4Hoc9t79KGV2DLuaqtso6IoJeWWHC6Xud13fHBkYQE/i16tMb7WG+2C6IbMidSw9
d6r2dhCkUj+hPGB79/O9/KiD5Xn05nkyKxDCwrTz8YQqGtlxVhV2Ph12DHKTm/M+
4kCnpVUhokBvweFdIUxwSbrw0tuZvnJ4qw5T4b2ui6rMd38pEHyTg1g1dXa3JABP
5py6XGzay0FJzhilf2SATQu1W/q/ZsgGM1sJ4kIZoqUHuTcjWC4DSKlfxYDNd+Mu
FYoovlCfzpChhdTB6ibAcGduK+gQPdUDk8V8+0GqUUn6nj/kRZHvhj+lIaILjexT
MUi7ztVMShLJPXzVlfMLsX7lCiVlRXfFpjZLIZF0nw9AKvw18nnvYcv/QIsYU8/v
lRWQ2tMEh+EETqIQO2JxVusfE9DjJgdiaL6n1Dg1fox1cvBcXNkpqllwg+IlZD4y
UX15DaXJLP8vZukvJuPqiN4o7xKMj23S/Th+SVKjIuityj7fxxcSqJ805RJGNi0p
e4bZJu+ntDfkV61Nwkvr5Ojg/XnFu/rhlthESXGfvoGWjnGWryd8f1gGW60vkhVM
gubXyocd8+vUoC3kvVJnLPj9fP8/ea389cEH8tzgSJiYjMxqKydrzRFiVmbCWTrZ
oCeIGwdFiVzbUZo0dGUniYZO6r5QoWfPmHuMdeZenxmp0+ekVlTsVKf353Xz/7Da
x6mOXSKXVw2hrcD/LCcS1ZoukVYK3vEfe9Nl2C8wvUexJqI6msgLwgtx6KNr3jy1
dq3Tg1A6YCTwZuBnpzpKj1v+OBct9mjyr9h8nASeGmMZoOYgjQ+8xufrmRS2RMv2
+60lnKJDnGWBDatksPPqvibOiqiIK3wMLyYkuzKOE9XDfWDKY6io5Svu7xPzTF+j
uosGbe+o4mm2KHix13Vq1R765iROAISiagQNCtn6ixoNcOJ7C87beqd/1W2t0Nwg
c1SWCV9KijPLndCelwfmSqxDir3f8hJJVNif66qiib1wITQrVvB2TdZZf+ql7gjx
WTfIiH+tWNTGA9D1GhFDPzs6+R/LFEMbozQxVQpyiYKA18Vv/eTBQDUTADFFvWEd
gfMhzsdtK9aWFJsKA+FrdRBvzVG/FqdTUmI/2lhCShaWzxDKufT7MDx6LFzElsg0
Kv+M7J7cT6ioEmd9JUk4Ca/V2Go2oZeRYvADkXTsB98w+auXpaNW2aH1ywAsTdQg
TZf0cSADD5qtX+aSFRtb4szovJk4ydCS9AQFaYXN9fstiy/OPqBj3CtFnVOiQMq6
MGnTca/q6g0Tw3k3Z661MW/ywtJXQoAeJedCiWJMqX62bDrz7ER7gKMvNgCAUE8I
IzxsbFH4rkId2itf+DQSSakVn8FbX4Qr6e9sBKubHVhmt+lVfENGQtRoJTLJtbcM
19yrfn/s2Pv0iWQjvxJ+rry6Mkd0yXxWSn/Q1aI4F9VJyzAfoy4yJcxeVMWaSEjH
dexiejHl55h2uGWKzzEmH7XGK0YvBbDQ0iEgmIcK82fj6yGkepr9hI8zf6odszix
6EnspNYSP/ozoIJf6VB+NGObL9KXwikPVxF4b3oDsjHvieXVY9EgoN0GJnLq35pa
rErsW06HXUhldVbzopgYR0UHdEn8fcMdDj/sjc+JCRdKN3kuprONvAMncnJ2VtwJ
LfD6EZD4c9HqznK3QLHFAMqyWl8NYGWcPbVMkXTkIfx+l5D74t1ILbrNEe7Tjtqf
VjGi1C5rGiGQRfDF5uKUMXR77QuzmscPhJQIzgTGN4XRFAjJA0UdHjd35T68hST0
bvQ1FOFa3luQkUkanSHTD3iCGXPGaJr1IZN2aaRNR8CY0poSnlJ6UYmIdHfKp1kt
6eyzeSdVvT2Cgx2220gircoS/I2YRfXnL7gM8AQ/5dJMyVppSxtq9JxBFUaQR/Wz
1bjgWgrxOlu5tARmFsmZZgMN7bh1xq/sbt9LCtLhYw0btuzxpA9wX0u2qINf+Jgy
8YBs6QDwn2upqtMjIz80QnzX2QyY84jOZzIIXDd1R3KtT2BUFrMfAUCH3h4DbeEn
ezUaSI96edQGrDncAXfGh46wGrK5qzWY2HTV9peRkLfm4w945MAEufez+qCmoe9g
5vl1BXX2yx3p62vWdS1Bp4gHIZUxU5X5v43nGM9NEogF6Tl9d8Q60vllPUD0AF5h
GiL/g165zHwnN3qbUCTpODLM/7xKFbKymzozBYyGV7t3pTiNGfeo7Z3xgHbcSmpK
y+r8uAM6Xv0mfc4m9c90MPIzPQdr+CaGl79gPch+pTm14XWin5/Ckd18dNmsOdph
xhVje1Br7GMAH5slqlyDEc5h2n1BC2wjQxiD/BKtAHoNK3b6fcFsGqHJ4D3xjDBG
ucWA2X0TqhJXzeU3eLTfXj6D9vJ4YaNrf/K5q9ohgm9IYTt46xwl3PFBhXEFa4x5
ZZPU61m3Mf9NyxHjKKbMP6waWGSznLk/579zSYryPVfazRavFa/18PbfHLz0PZiM
ESEZ+tt7/QpGD6ChHH1Rw2iwSFWFKHv3X7XCX0fXT1T9uzX23/BqE9Lh3vyNNiNy
1v247rHGfBhdOPphWzPaFehVhEnqTHz+fM1di6oUY3O0Y7B7KMUyn0GBodrrxCM2
Bo8m/lqZIZhQLinLynjE+YQo9sZ4iXUzTlniTS8WJFzQGndgaVJasY+5nx06Ok5o
hjDG1V3HatnlAG4DItKcsTwduajPJxlr3MRzvCAM3ak0n+/RP5YQAlR2MoRKEm8x
xuBhqc3l/2anMi/Un5zjMlCZa3atsHceWxj/ut4oqQ7mdmyAzXy6uDuiUtgDfWyx
byfvNRtym23Gx4nbf9AVbWuaAm1g4ODofRVwONm7vsQZN73/kVBqpnxuEvi52gcH
uCmzAJ7FryAWuyQFpTtmFuDWrC/VJ2TwdB1VNeYgQtSN+DlMs4JJEh4HnP5X13NJ
gPhfAXcwA3RYNjg2rrQka20n6r7V2RQ4DOmXDLpwpVRuzVWCsnzuluuPbeLVq8DW
KuFdtOd2rFSH6KRdqmvZRutIduUkwm3WRpn4fI1B1bWa6z1PvTHYd7qjpjvG+OJ3
Np68n5rMFUyeT0HkgcLoJ/GiJ7qMuimettEtsxt8KytMCnMrGwcKLsBmZn22vtsr
nELOJHSyomcaFHM9ZKaTyn9S/mo7HM82oCZaAmk+yqbRJylxPB5iEeONzxwC0nSo
QpKS1rV3kX+1y8ji1YQdgDmovQRJZ9DCr9kRF5B5JjTtdCEtUKfsiX87v3Pr7A4U
QSHWNeXfD36Q5j7QZy9oK0y5688O6uoLTrQN9ov/DufQExrRZEosbGus3MNb2bQa
m581SprgHAPPTNpM6utszJ8osxe14fkyG+GhBbxZLDT0FxkvdWvNFKX5GulxMzNU
YTURgRzrHeh0sXD1tDassHtLMc/XPkRVrmr4FMrnii5NaRupP6SDH7mArJmZDXAk
A1MCcDbjM7lsnJo4y5glhgfxUtvACw0pjclPH+aOGUtUfCxcsLTH7szh5gNBC4v8
Hjt8TYQS3KmeRU/yg0MaplvmFNJS+ke081xSLU+E/YR6ZRT4mm2Gc0T0V2bPDJ03
//QuNxQbTNmLM1O+WVtvim83a+OcK5IRqz8GS9Y62oqQJl0TSzw3apSfysR1bwyB
un5rylhUThYDWrIbbJqgajxDGAX38UVKvDzMg9LZNe4yfBzmYrIpXyuQi6Jw6Ks2
j1PC+1giHTnOGhduGUFcIBHw2XA8RVjBo23NdqnrY8DPo1eSNwzetGhxM8xMGtOD
XoUXLMy2p8TP7kc+KypYfobEkuunoSiZ5X9JACBz6y/HQR7rmaK5rsWPvJM7Dmah
tE4kPAo1kS0/wIq6VVe3ypznUUvBm8/XLGWgadjH8+/Vh4NPfdnpku/NNzbke1Qu
Q7/8ybHi4XrEupDiooOq56WMD/xUd3CqPVzuNw32kXQoxy7mXcottzl6SZCbKvCQ
CkiBL56nGmuejMEFQJkUMoG7Crt3KqCxXFgQvE0h+MBdip62tSRsKdtkvFYgK3vm
WvVG/iYgjLwe6QobOU4agZwsr0Eu74SIW4QQ1YfSjWkvhi5B2kMdQg/0qlS9V5K+
QYhyqXEdq6XlPApLgT0/nX2MdtDFSCm0+G5vP6Thc1s85GymsFb40CaXYCTpwl5n
gOQI1JYPOtdsuDwGhObypyK+EtBOTJinjCKLj2UYu9lSLSE53HTy2gUl6p7d1kJs
FMmmSy2TNkXpqgQABimdKMCuO9SCThr+4Qz1Sq/HgD+VHsYphLj9LnN4DiFokUfj
+vrA4+fpUepAq5XWpbBM59iETDq+BoeLZaCEjHBbP3r+S9ya5w/4gwBhRi7n8jlo
LY5u/HoU7UjkXKXI2lBw7OEJW+rhVPUcx2FI8Gspm6d9PVDu6+syyDErxCpl6SFc
9lSD/KkaEgnHpIblf3LPMgiP2SB6ILyli+LCtYZvjuKtEg8PwoXMNk2uyg/m1UBJ
oynCDuH2Y6Y7zp5BnbRvs2ekpPLsxA6IG+W6Oh4/34WvLVjVF2yrLl3aCrUD3Jju
BQmUTkTCyw5i+t/XwPXWqsLFe9m+7NCkvTensKOTFm0xAv0nIiEhaZiBTjVMUt/A
vF8rlpzti7O3bIIATxgzgbGNqnewBhlI5HecFoh5x5V0BbvMCvbIIszVyOJnqFhf
g5vWMNZ0BMKLBvLrgmH52CthGhdwvp2zYl+DieXINEXtRr1V6XtDQV5taxnaX0yK
5ZDsuipsOXpVrnwQPIz/OkK6FLUlRcR6/k4voh/NVy1rqH0xRDHkqxMFY2BnHwwY
wj09W7LeKkLAc1nQsCkzYyhivgBpmUNhl0MPDB1pm0mKen6FFc40uvU1SL0tz0RG
Q3Z3GpZLIlWiz0GQtPYW7exWbXHq6y9rJBnJTzJ2PRUQqac7R1TY/UUUbVz+73/j
sccGF6RilJBWKXdJkuftrsAHp7SvLa9/Cqzx6F1H1AcDT7erJKbwMmqaugXJfKv8
IP/BIu2nxTG8kuv2dsKt38fv8iQbZKlL7YcauLrKfOGHR0igCO/y6C6tNyd5eA6m
BwoKxRPuwT3iKi4ntLhv6gt5nNqwc/MwoiedvGtTyddvZf6T0TD0oolhPre8sGl9
roFnVvuJuYIDx+AvZFUq7b+qMhDhVK3xoFvpwUacyhvUqbHjl93psFV1q0rOMc85
TT63sRTr9Cn5NpMXG0gcbFA8rhXJAvmznKgjHjjAVGw0RMCMpHSwLCl1jCT0eIUq
N/BILu8V/WfvULL+RPJBZV0jiClZXfN5a3ZjCD3G2Zoh7BhlPenUySquzMVe1pqd
gH+1KdOd4oLsqhXcfwcLx3eQIcKS+rQ7k+Z9DwCR0TpwojjpRShcpsBBLImMqfM8
v5EKIWTWR6+ahZSXVwxjOS3RISWeDlO8UAn7/iFLB1h4PQdlShSYW3ySCT+UBplw
lwm37kxFDBYFQYM+lcEbrxx4YfTdG4P5zHRbT8iPth+uav7k6q9mQLlXDKL0m88E
JhMDx+xYDZXBc/PKQC3Rjpjq2SlAHpzCM6mb4lmxzZE03OnQATr2VSYA7lh7kHKl
glDxTxL7oEAxgW8aCkveThyXVU/5uC1Rs1sFfZLPKTD/yo1j6KztbomujNUJ2jPf
HjYrqmDskIAyCl9Wsreqo9OQ3yZ+64G+XbmP6/QMK5H+Zh/v7oO3LLJIzXpnF6w1
6E9AFarbWaBwJuLCfVhMGX4lscSdsPRwLX6HpXIQ3CVhFXO2ON3GLgttF5XPak4c
iRxnTxzncdWMqkpoh4GveirRWlb984cE3Y0r9apqISmm5F2IzGIuufGxkSwKQhkw
xciK07gv2JKJigtKXF061T0BySp7swLBgh8opXPEi928i6GQXljQcigizg1QU7Qy
3TBODxINNlVaVXSOs+06ZfeMgGnYvi4L3BcJmHOVTgzj2594QdtIGd2FHnNIMjYg
8gwoYMDUreoTF5uQEVjY8/uTj6sXrsrUSMqjdxZxYmS+73t3qL24taUagnZZP79P
E8P+pptJ5wXqeUl2+58I2O0PbQGm3V7GUJoDaDrX9Z7eGzL4VKAG2LSV6t4ds1lU
eapAAIP7ppjoZgfifdpkdy7tbcvW4kKuLHRbaw2BKBkHewex9nmr33bWaH0LWGKt
ObMjf4XniP//uGsWSXh/SHrYucYDEXnXE9AfOhzEjqJSar1+5yJ0dEzH+XwlF5yB
0zKTbqvfnQSdZig3N1y81ENb/uW3HiKvyqA5ydvKYMBqbPFnjkaBpdpQjlAnhbp/
lvHxeGbKyQ5BNNkTxl63L3W9AW9N7+Mga/xZu319vxRw22LB8AOWpKUzkswbJy/G
A1KFpCnD04lpxQNXQi11gx9UL0ISWZEaGu6p2bK2Uas8pkP005gKgoq7w1/i2tOO
mK7iobfaRsGKkiaFO6CQfDW4+Fv43Gy31OQRPaVB1IRxLQ2L6GdLJRNB5OAM5e4E
b+gh192dVE3QpCeEi8hU0cBqXKk/bnpjyyAFDL49brRskAEGNdMy/9Tsx71BXo3Q
VnDSBywRHtNqTfkVYvYWy6vUjP6YdMgaVChjgOYlI0TH6QQe+LaXdBkn9gozpCT/
Y7vUYFhl53eMSYkRcsvAfRDiHls0aRyWwBprm7XSfKpS28khgaTIxXVicyTpRdc1
GY8YT9iBAmMAarj4zJs1oeStZt5+t//ECwHY6vH/uqo/aQ69XdJ/QrHmEWGfgaNe
Z4tIAU3yK0QhjDn2BfZt5JzPZ1ao/UsA5ItiB8RJ82igSxmKLEFFKIeRPuSRXMP1
hLaEVB8r318gPPaCou/3t80iQJtESkbo13MddlZ0khc7VDcvB5PaZar1bobUzVje
mi1p+Em4gDjOqvVXkbu0p7qWLUf/VF8xuZWFrwO1ilpGju1jt81Eqd/ogcNAH/4K
QlZN+pz+95IKvC5N3MIvOaV9l39IDbNduI01XfLPzDzisfzibrmz3uvnWoljBFI8
OV0qn+yAjTXFFt3mkywzt5MbnyRzhl4+ZQZtMphkW1gccbmpvJy4brEImEqXkOX2
GP9zW1qV+W2EaHI0R/tj8NCg6v8NHr9Yp5oHSB2mQPoUJGJZXjlSxgKuiBWEI2wZ
j/tUjC9MHxx6POzP4I1hBri2+Buivvj85LPzl8I2OBLf1L2ALeCv7Fb/1yJNxLf1
BWPqTu7rqnyzZ64fAIXFANba53s/rXPGEWf5vmW8O1si38gwQULzy0Tqi854Y4Qj
ZPZw9wurffrJYBFsiKbA9AEjcXqqhIm4W2xwteMxxRmTHJngXaWxdCqNXdhxwxmz
oHg1kGl975rVTgdcM/YlVbKblevY7dImU+wTQmYcA/S2ShYYcQw5KYZKx48peBQL
McpQcl0qEVCHu6WTtlrjZDdhFEGZv31obm1UBwvvbrZL5ydPXiiAKR1vRXtlCivu
71Ji0lC8cG3hMJCfVUoSTe8+UVdaDJyr2Hr03lfVdvafJdxTXNTUMg9031L9Ffp+
jZYF2dlXx03+kZhJB/34WWb4Jw0a31AM4hlMBgG6bucK/U/WP6VxwfjkfqpFfnMW
O3Kl79vaUXM/Mv1KtZkVx0h+ZzHPn1nMWvXQoariXoEUJrgmEocNJ3Se5OkJhr8A
xRqBYsWwA/b7MV1sa7tu4RcKohhbC5HJ80Km68/kmd61p8D57FovUhOGBRrlxK2b
KP05Ak53/jDOtFmlAMJzKDfvd5ZMlmy6tVqLaYWD/AbHetu+SuT1IYJXjjHwvr9/
BFj50sq8O3wsApPXWZNdt0WqPXpHv8im2QG9OUhiRQxpmfCi6xgmYcGk+UsXNHIr
yZz5BGpfSVTfm/Xb9UY8qYZZv5THgTm/kL2uED+TCl1uhIdKYuToreGxqTDSEKBa
N/ORq7HCCUJWllEdBMsPfvvqLLhy4RI3uJxkijujOYfED8MuRcWjcgthvT+xAqsl
Y1x6KFoNrYwutF/LompohhRHppMNweytaauCTMsFuP+EwgF5VrcTqa9SpQ8mJ9/A
KuT9SOntkl0x4+YHgHPKeMbadColmf9wfhMlmVbnVu966Ro4A7aMVRWkI+9iPz0Q
+gBhBfnETzdJfu1ORMjNjBGx5bDLTpjbz8TvdXv686O9osczcUuLQBa/FAonCJcg
enn6CPe5swwisZ2gkKL0X+3W/7926j25IRYFhyUGlzoUGeaunx3jA13B7nWKXC01
BqiEpOCbbKpSFgZTtc4bZPPtfLT4Coe+Gly/6VDKMk0mAw/+/mxTcDIu4ZChxMCd
ERCgBS6ffO7SvN1yAOJC6Vw3Zsc9tkAaeMbu0phqLayZcF8Iwj3iUlO7Uujhzamu
a7KtycPSWFOuSZgfWQtYA8bZdumhqqgmmtiSYmGK4ztT7giUX1YoBER5v1HAxjFi
bvcBTYjRF+OoghCHmHWTi4Sjsv+WdT+pIWA7jyCRbgez0UwmGP8tHB/bmZBG6V21
YpWSn3e64Bg3qndeONVa3gLYmr1tA1f/cp7kzkgTqmV40sl3C01EVY9l4obdGTU7
FltqAORikSnNmiGDcX16sKw46KUQczIJnYSEKBCn1lZwavTh/HCBwGMB1bygz3OQ
3kiULl+xCRORjGijwZbyuk79x2svYplAqxSbfBzpAsxmuKtlnXT4QQwXlEFqcjgm
XUs8zKlXue+JJt3rVAN2B5lXN6w7vERjKccKegLRnYWuHk3scYQaf0fnkdpFdiwW
NLHlw3FJi659R2XQPG8JQlyFqzf89hD0oXMDOPmLMcShrQNuT1+n5DE3OEvA96m/
eFsrNw2s3nICrU2Buj18esfJYahPGaOMUViGgyOYZzMxfwjgqE/8oYC1Wfup0eyh
Ssp85CLIZCMCHzhIQBb7GN2zYMBhKklB34Z77hAZgvDbbJxf23JEq92NRYS4iB4P
nnThA74AWDWrwZqGsVhVUmz3152iLehTRezUkzMxdKQ7/ait1ALANNPYDYU4d1Lt
ATD78Pg/an+1lrv9Ewz0wuEIOmMNXlJRWa60YJ7P/h+T23kEEydJTfpc74RlmM7u
coc+Qz1UzcEYHwIZErfRVf4G3yDRHMZdfz2Yuc/2+pUTt64baiEMsksIbomMSoGQ
3cmVPrKwn4MZC9dRbjkqrVvnL4WDkrD+stm+XK4KKsf+EYMljIzsTYzEQn8vHOqy
Lqr6ASP7irPqpkq0qlxB+UP2oUzfVlKuGKhthRKjIsJaAWhvM1DhIshCaholsA9D
dmbEcADY4NF1CmOXsHK62D46OzsySERGgxAc7wnrYlohAuehgUDLCFiSANc9f2Oa
73dF5ZCXf1CAdzMGtGDYQ0GKd8RLMyX77vDRIg/wPxGKf7D7LZQH9XP48vUCBaJH
uVsb/6udnTNwJXED6B+kkaqePpsy6TpVuK5uEgaHL43mrStb7k3Qe7ZI8VXHISl2
HqGQq0btJ2aDlChmt/XzR1zboE5C1ixWylbIaKa3pUafoJGSWp7qDa4N4O5TDlS0
UHvYr05HJ3uQUq19Gngt5gXo1ENx+x6H38VBVRdjnx8JrMteb5oBMDVvH42Yf1pR
DMR7iKE0sfKH5ULTqlMYpDwsYPt4buY86pEH1j/Yn/ndZ8rwuW2qTpnWhm1ttgjR
yu/tJVaidBWZivBTt7Uz2QumUHOdhORVToKCy8wEEp/rMrXGfhIExNjyzSxpEcE8
tEW21ki8yxITpGaVDm4ELkNoKRkT1PVJae7MWnKQrDNDXe/s+UoYuo8dNo/MXhjw
mpvMPWtgeSRSRVd8pt5mM3tfVRjweHV4csP9buUy2WmsQb9i9WsUhX9II0r2wtZq
6ewelburP7FmgzFcBjmg+AutAiAdqR1alDxXA8wpHovHAxeq8qoNu9KbYewThhuR
Zk7tGxxRGtAeoKog4N7DxNARWKBc/ovQxUFIU8Tw3ESSqW20zJfd/Y0mZ/XYBTjS
prghC3BwZx1gsc0j5SzIRwcsd9nn+nPToXED9G32DI5j0QbW5kAQ/lcPufO6kWN9
xnAK0BdAbk/3e5tBOZ6Tbg1+iFf+wEE2Rv5IeNkLkWqLIPXDRGXFrkKJXrN4WCC8
bdqDGF6WY6XJYCHE7wc44IaA3fg1keXoOWPhYnrx+eRsO7cFjnnwsFn+lLaq00OX
ltT7q2ldespm36r0omhy7+c6mUcGUt0PxNGuXFPsDWL29obcQHlj3SQq4ABw9oRn
ejZX/+iCb+flLYZLVZiEiLZsvvX8vDm6Eh+dSHAQQrQupxLQ2OMyIXKgp8fl5Q+G
LUDyE5Zyy4i+4BCfA22M+ninkjn+8vZj2FnPRtsOS72GpTtg9LMUIVp50gNn6/83
PodcB4wHGgIlyy+7OyZmcSPbFGWgbtcWUzOx3j9HF8j1du8LGSty433fbHmbLP0e
bN6+JS7f0KJSK1KrJo1qVWxqZSxZDcoccyAfbkXk4zE/e2s7PBqOE1bZnAuBsham
Si/E0xMeARX+l+ndLFbGwxcyGOVsUEtv8//fcURH0gAhrNMwZYUd69ts0nCfrfQi
jLrM67cUKAb/YHxMobkSJstP8khIkQ73/1q0NibCyWESzDvbIQPDxjuMVFUsquQZ
dovM7d66b+WXc20krtstdhsmsZcUvVLByN45oYgL9RyBwIlV8ZB7NtS8eO7kOvm9
B8TMvEZGsM80EzcnQkmZPa7U6VFfxH8SiWNWqspN8ty62tSF1D0FMo7qBFAyuEKm
LpzQsay3nqZfLNn1t0SvnKUTkNBNtTPlw+exGk2h2C8WlZSY9e/4tTRfdjR8Y/6G
LSJQLpEStmwKht26ohx/cTUZubA8/F8lpTeKHXph/EdxDqER9Ii0tTd3wBPPOkJb
w0to+cF8luRGdhiO6OaEBpbgQYlVBK76XZ3ZtFA/Zxg6suYhwcO0YJK1yKfagTX7
1KtfYjuwriZkQKnUy3UMph4jM7PDIxqa8a6OZwEqBw6pFPO4hUG6Nl7IeskaHkkB
upI9alchI39Xy+hDLU0jhz/8SvVvlFi/GLjBc5XBHbsFyoTmNbKcnp4Wm5XVgkvy
bJmnq0QF0b0Aez6cVF/sm4NDvNoTqZi8Bt8GmV5uOjS6nk4K5XwBQ/sm7RmM/29d
BeHo7+AxYnVpP7yCJDXFoguu+2Pp5e0aFC8ElkSahKYkFdOZ21W+qFtrEkkAsd12
7fZfFqxt4E4S38ZY0sy7zzvOdRblKMZFvY4Y+spYg4DsNbBDpGIMdCu0VW+Vwi6U
jBnPDmOKIvPf4g8Z8CJDQKcDR13izqqM5CbCpdL4JAjHBOQSirbWTttje7QTVREI
kai3oQHfpA6bmMhqjnHfRU4m1I/ORf1lwA7vT7unWha58L+M9PEiwIixV0UUdmeh
fn8JVFsNgr8yHnl3I/FoAeJGbFUUelumCvfP6T0/sl10JOSP7gFVcxh9qPKK++bF
1ZSfask3uH0wTzURJ+yXjHLs8o9+C04W+AEpTZai/B0PlRtToIuBL7/gP0I6lZND
+q/sKtjKeMlhltrVT61otwUoWgUWYPcxvQHwMGGod3n3pEhpG9gdrpDRiouNr7Yf
GGJC+RJRPKf+Zj5dXj/Ua7yWgY6PZihal/WYzE+GB6RvhK5l86ROCt7HSzd2KdiJ
8ctG1Rgs7b28IaGERgKdPjs7mr+EUxULLw7Ya2povGLUsm6hMh6Im2Z+IHUazLBc
SCJ+KJkshfASox2J9vHOys7B5g5/pqwzWajzkK+UPefZZv8Man0rJLrsHLwfx8fX
lvdIJgk8r8oy/nK6cu4bCPimnxvRPx8dgBM2PHLu6HPRjrerYPCisM//lfRrNtIJ
pciTdqLqw5kCzQwld5YfqXmkHSVqIzgIWW1CuUhZ7gtaiiJK0gMZ01iMcpyang35
LPmctaqAqc/mAwmQEujCtBylhyj/GSyrqDM1FLeofMVF4T0H9XHTJmd1aozVly1o
pp/Gqq6gRWJxiEZuWvU7TgycEv6nqDe9VzLaF0xYhptznt0L5654FlTZQl1C+vAo
USzuKYtYO8iNIwf+zEgXyRY5F3wGstttiwtqKMAmZCv4hxIz0G8d7vYQzlve76DQ
s+LT4XSzWBoP0IPB3/OtBCHAuidJzVpg+Fl24FkSdmQFMjDgghgWvyK3FJwOOz+o
n43OR3H0Axcf9HXRLvmbBDkAnt8O2fKVIc1k0aDE+gHuTEqBxfzostKw9QVig8JE
h/pqfecnd7cGxkQ7DEr8CfXJiOzMHfGZdWvk6pAtDOoxWXRNGuGI0IjSPQbzhI9+
lebM4PRFBsRfX3pTO9M3DxmnFhHVPCtMNMGTUIoj9lUe3kAJumGS/Eu5rjQcPZRF
Yuq5Wp0kdnXPYKXqdpWK2PHn7sh0STyCr7fXbFSM8+O4QB9ZmG0CYT10NdghSVgQ
0lWlG0tKMh5EvkRVRzKYhJscBm4VCXkdhQHKlnj2JVGaDHsqQo7NLrPVviDT3FdQ
zSeHOMS+E7jR1+7tS9EWqFcvzfqOMCe9KE+YLb7xi0LKHQu7LUiB3dSsCjATavsq
6U686jdd6/aEmIzXN32Fej/neaCBBIApgP1eNqPA/uBl4tnNvIO9zxlgIWU5ruen
xDfKjCsgUfJ78vwy6Hi4+R4fAe5FmMGKBJxo+GnLH4yffD+bvMjmYpDR3Gs+sfeB
q008TO1OtzYSmRXK7g/v+4F7CzA/BLmrMQ05BLLGPgeenHK2oUrfRMLGb4Dk9JTU
iiLeTVYWA9wvUyrHAr5SnozmmDEBG202iUPLkAWW3L02S4/l24h4HhyZ0dBTZWog
XjgyS/LCKHeI/xwrP4Fpum4Xc4h9onB0wq/jzKBhICAzs8Sai/XIV3DaXjlYe7iA
eURkvgYclb+sMsxf7Wm7BDinRC+Sjhxvc/j1EWrak2kpWycoKrFJ4SnOQCHvRYc5
Ul0Pd+1NmXPEZcfv+L15H130CtDG6QTYGBo3Z0PbfByP3K6mD3zW73wteeyYY5X1
nFsuEzyf+yRrpz8M/CUsPFqSm3DWEhRqID00Iy4+bwCI60DHNuVuG89Lu3plTG42
O2hs79F9u57Opr2Gcb6ifDOE3E9Z+aZG5bCKgcu+U0i7YsSpys/n7+yN8uXH0Y+4
Vp03nzOsjiRiKS2RVkchUrs8X5d+pSGGYphHpeAmMjShVvt7V9X2CxdmaEv/9vtk
c0VlF8YyvIn6TxZgZ/BuZPlv7YIp2jGQ5iSDg6bC+6RkjlvHt1X4EuV7+PbPRRXF
AaI1YwuCcGCur5MzViIoMJocGv14/oNbpLlA62qMrS3OZdWh+urrogMv2AwsZSY0
hiuhbXjK3eLPoBg1IWvqP3kIH8b5IjoN9tIr/08Oymk0rSKxWH8SZc9JYVsWOBsa
CPbhnFFaY1EmZA1yGx+LGQPz8jyUG8JDR0gjG2PMdugdcNybKbWWuNcJEP7FpA8E
Mgdp/xF1GZ1e79WmREye+ogkDUYWx/NU6oEGlcDkEUpTnPvFlJrwYuAfQt8mhun1
GMwFCY2vRkbUya/8XsxRKOYAaZGuAhf9iAuTBhB2mjZNieB4p08YD83s8g9QkXuH
FvFNzI0Ge7RBwqsL0XonIjoSbGuHtqeqqA5t81a/LHflsdYiFZeZy8m9VcETXE1B
El9uaJZ2Hak1abISGopgCxVEEX11+iqfbw0mgvOjA7YT2P8G6YwhKshHCrkxQWct
1561a/Zwf5WQOpEsUbLIAeycY1BY/yP6sliFm9w2/POlx3poErDhikntXPa1flCw
xgqonAh1wwsPzEjFR8ttIja8FpUKbLLVAGrE2YHbDFyJVWLywORB4u6wgI0VcrhX
d/IaYK6ztGOvBV0ldrDI6kGWyrbpMsyn1oy7UzWHo71GoiNgILu40Kdqg8hBIl4j
dxonTVK0+N7OFiDx5BWQ+I7IK2OCLxrtL11ZvxljKvCqOoCzrXRY8lH/khGg4nel
OgajKnigcD5rZ0cSiL8Y5Hv4XJVDCCGasAdvx8eXr8mUuLoofT24Ko9Y3McLY16D
LM/6fzqDVj2gARKrExqbJPhuDUYHblV+DgLQrOPtFJLzZXIfhQSpk8hyLSWFNavA
jjFdNolYxjKdGEWC2ybUaX1jgCHUmz3q5YTl0wf5z03AD6IrZYK593mFoZX1FREW
bUc3Ul35bpYKLL7SdWZQ+/6dh8xw/Oh/OfKnQGXwmuL8mec+2lF7QZyTbPHNwF9Q
3rX3MxLPUqe/vpgpRpPKRTJVm+Vg1bXeomi1GBgvCQWfW8iV2HDc5NM0GxypvRoe
kEninKMksX483oEtxddFAXS+tpKNY06/IS8Z9jooj+9TW9pfRAdsOAzmsF9kFNtX
S8cZeeU8j1qfgH5f969jWkRXJSunot1tZAVmA70WaRVA6n+7vfMWxtzKF/6I9DJj
EGD3/lKtitVB0Xmjc1XSCOEX7hOcrlwWdbqNMpmFQPW++Pk5145T/9VFH0lbIYZu
ZszfNqoUxG8USibFNdbAc8J4FbEC+RbdaC7ZdmzSGzL5EGbYuriytNg/ZZLmKYwD
ct7oVBXonDsjNv9GBQ/t5xKkNEu4ZE/DU8nhtSN6ogkFCTTe8/2rIPDzChS4+Dst
dcFb82I+5cIvIcTRtsQEcuUbx0VfHJwfXw529nH47k1uNKdVMktxFPLWX5RdESUu
tpmzP+zSp3UoJx/OTr4Rnx5o64z0K5Wy8S716wuXCIc4mc4vdlpHuez5Cx+wF/as
z/rxC34jhYYzV1FsnCn8ZbgbUNaX7zdT5ijHjthakC071l4DPmQsxpP4ghd1jISA
egW8a4O1ezKxAd0VrqXdLdqFjIsyqjun69e1ZkPzPvqfSiQLSl4tFCuf0JWPkDUL
Hb5kcF97YDaievG1R0L+qELAgS1gubYNGghXvSwePCvDrrW+qyOUWVM+NByCjqJj
HyNpGaDYleRS+d9OzZMHYOlzyIBdmKwlP1mHnUrNeINqbMJS3KhGONDFxcIZq17F
4OF+oHeFw8sVBPQ6j9aF3+UkDFfLktxu7vHlwAweQA2V6llsnn4+xQyYFbB24HWm
i5spmCHJDU8zR2z0oFHp2OBirjCP6k+vZ127Fxx93pFMj8B2R6aqqH9j/CKDbuqe
U4c366Jt992eeUhk4jVyAdloO+61qrAKPuudwV4pAlKix8LJRyMsDUt62l41XaRX
1jygWfsLp8+zGrbDSWiQBKZEllc2qIb+fihcLqezNtZxgsSFhSMSSkx4+qBQcCNQ
quOZ59fyR7qAibl06CZ3RJ9bE/Ab2BeMdVSnO2BZt6XCXY7dmpAZnAXc8yMRJNUt
akbw2spCi86lSd4EIcT1T497mkwuVyM+eNU6GCH3J8uNqFhEU/9/zWnxXUy5DpBF
BXxxsIY9dVb8UUNriPipHLS4CZuuXY58ZrZnMKQTXoJfRdGSJaCGSFJhrhvalBqq
e9TUn7TKQTA5gOQXGfT6wL9xpmAghtB+YQntOJ2zHLUgyw29rpPcdZD51OO/7FaT
5O9cjzPNFzZIvo5Hb6NYyHT5FxYwQ+9fASaQVeSRedFGNUPtcaeLZQSqb88StsAQ
IbFOJCrzIzcn3wx8nCXk0dM20wWyXkTpJDuKfUs9qvrNqtJI58ZBXWZeu+Ft5WRv
F2+CkyuiQweEEdvtFHeQTV/FZymkEoMNcuUtwbIXq0GU8LjX7DK1aaT+mB/RZe0t
Md6IbUMCmFu+q1pKr5eknxxOV0Rbmcc9yl6Rs0H/9/uOTH+9hkOVmyc4SByVP0mO
cEnTPl6e4IAtiGNagz0VPgdSR2oHtUd4Xdyjj7eDKrmCHmUqvYPxJL5gWdARfmgk
9CP9Y+dGK4XqU8nyXEKZHQn/hvJ7ktZ0K3FOu4E1ulP/zdZYBOd4Dany//J8Vlci
P9klg9Ma5y1aJqb7deL4iXvVCB+YgeE8wzn14X1OSNdhNtd43WpFtX7PlDymob/T
aUtTGkiIargwqr59MfSARIntoWAVMmEJG+VoyQ49mf0TlijguwXmadNu3l4Vio7y
LOPleGSl2mKaCZsh3g0gFg2rfvBpDShY7rCchgzqsgWdh4HbyY2y02MVHCcleb4C
icvNsmX2HDUvbDlRh6x+PxLP8+bvGVjywxTx8Re2mvbEdQfPVHklOq2C7ZfMETnF
xGR5JVFw2vDokZS8DIel1eBi7WUCLQwh5bEC/aTOvjj4tQbrBSkc4ikxiX9yAWwg
KSzVKUJ2vPIXDxWtQSix6r2oPNmzIMP4CxNKNCu8NGxqUhlSsSLD9lJ8jgOLwF/A
YQMFKKPDFyOnC+GXRJOTwNQtVwcRn86xs2ET8fOg04ax28lSkkiOFiO4gJUncp83
h2TXtoGG2zgC3jStzpU3iV6RUJvjkYX/iTY94stckYw5W4r3NFKbUZZj2sMdg988
MSBAugJEd0f+JA4B6zhZvyNB0YoGO1QyX0N/Kdr4EI3xVGTLCeQyfxnHY8kr/ZEv
3vkH4LqI2bN3eg5CpqsxsV4dVzaD89ZZfP2EaMxXWvK9Eeys7AERfoU06ucAgVYL
PJyHl4GmG63Bqzxhg9X3kehV+CnFgb0liAobMo/W8co7PqDtF5OIfNapQbjE7m/q
5dODkh9ClkgVjKZ0hU17qs0l5+9dCcAuK2HADQgNPUOIh7C6OVrKAf66xDpZBjsY
oRtke6wnbgPCouswjNYT+QSvryN2+raGmTxIzuTIJEEKs9voRQ/sFBu4YE3ZFZFb
tn+6WNB1bXIxhrlG+1v9fdCUdWOaE/YiUUKR9P18VPxrhYmY5KovZdj13WohGWJl
nulMGAwo44W18yGfnlQGv1csqX12gFJ9G8hyeGHzB/xWKb3t3lixE1E9gMxmy8RL
VcAPdCGdgKq0rfOodDW3ArsrJvWY+iNGfFtc4s/fmsKbtKtzQJzjvo59qQja4GkZ
5h1ORPNQgZJeFzLwScg6LnWnu7xX09wy8lPPi/jNz+aAwTIIvW93irJcbkkpfptE
X/qAOkvqD+Edm7CzsY88xeRfWn1YH72ex1x4CHYnnf1FPhhrn+862AypjshDcfC5
T/QgBmd8QOwZa068gb91imPk74qhq2CwVPC4jvGg7+mTNmSgLnkLYUs9KOenb296
jJA6tuDxOw/jyaVF7uFk/6tpybiilX1xBWFFKvQepgKCZrs4BBesQnwnl9Ovi9MS
H9BFc9uZn8azvdmXEM/9XbjNT+2JeGm0wu+EUYLrOHBIQ/xw+jVwQAIQoZHY38bw
keazJ887ornaNYfGNkoCvrYeXeOpAOhmvrL4wWZFt9/QQwiqU+onsrHM4RQi1fmF
Oyfei0MZfuX2BjJe/47Ai6NJj3YLvd5wrLU13wBjZ4UN5Ti1acJwj/sCHHqpyBsN
tyfk5VZvp8nJiB7L5J7hksPg9mtjcNhzRkhS9ttIfJ7z5ERPGWYxwt4Xhgp/H9et
2owoubiVTlsnhE7poG6LpP0s3b3WZ1rHLYtFFai9ZzahtxDkvEmwEH/PvU1NPBjI
uGRFSawb5QmOLKBhtTmiN0omR0u1Ms2j8+97HPfPhleoMqWxIzIldfutk4OCu6LM
T0ZaF8xP7u3DYkt4yEltog9qFqRv3hXqim9ZrJLvsaSg1iobo8qhbcESFhCSd1g2
166SyT88ScODNJEeqse0q7w9csHUdjUCcSylaVXF0EmNrCnnGNYylZ3GEdGtUWYr
BiayKTZ73XtOvxCvDjWzgMM+aJYkvE9miC6V+t0s5IKN0YQDGy5prml3bi5qJ1u8
R4RMvK8nnUexf11QKAWCbxBEkJyypixUWig5j2dH8sg5J8DqCa4PDebP9N9FfbFk
9fqCF05AsOXtO9YPkObf6qEird6kQnkkPoWgYz7UvS6zBWO1BYwMjjpK81Jtf3W/
CBAIPDHGw1MnDwkC8N7ENmnWViFDfjJRoC0u/O0HmhdJBgmBisnlcL9dilLxLCgK
m+dY36nT08mTJirFqSzRlY0ocMFD9zEABKhlDR6jg63krd790vCVEygiylN3GEqR
bMRIejl0ZTyOaLs2lWLall/3k1DxR4L4CEhZKigyo3uNZY+QGkK6R1vb0YdALr1A
k4tmW8mq9Frhece+2HkQ9ZnBihmFcxwPeDkdxyFG12Y+3nd5QnZMc92agIGBVGs2
G9+TUXGtmrmKnzR57RK42EirLle93nKjCHYjSM8LYpCVVlA5eTB0u1bXmy4IZ+2N
sQmC+HiqdzbD0Ol06Z1ZykJe1iOHneXUR3uzUFwJ2fqdnYpmtoCl96WjHaiI8eYP
mjtBjTGplIurvGdhObs2KmVgzyRWkcoRqiR45CXxQ6LJ5lAq4SlrxXmYZhyXHOEO
AQtaeSnsoCd3BJqkjYPD/whcZKPiyAb6PwRTxxAg1wiWwEx3M8FBLHMb6rpoMJ6N
b6LqgAHZIgRNelqc1etaxc4XVRTiQpQmzxevYAhSLzeLYmHy1OhI6zZO7nuhYXgM
5c/EtAuLgExY6kjyNPJyJ+GoUd4BIrgfg+8lqiQAH/S74oObWYXRbxkd0aiecSmh
Ef75ipy+j8tdBSsykMYDMiNfK3ZRyqi1INCa7uWCx+2D23zu1C33zf+wepNTTogE
Ctjw6EN5AJSrMex5LauqOPHeOqpFLHnkNCy4pYmnMOLVb1Xl9BC3qfvAROQd1bPC
C38tipdxZiwwD55uRjGn7QOic6AtK2DKFdiIbGl4Lqo1WWhi+/t6s+OH0Zs413sw
jy34XedipJNDHgxLwiECprUoh1NJd85+yr4gfSRrNVmCNsG5P14aLcPUY2/f09cx
OAp8SSbDNIMMixUjuxf2zR9TtRShLWSHv0mEK2Cd9r80GvYt34GfB7Y5PjmKMhYI
i9ONphsJtUhgpgU2RTengggautNPw28SqL2fJQ6oCwHiHtw0lFYqcDvAE99qI9vX
e/5T/k0zBYaqp4wdEL/bvvg5QKUz4b7nI2Wo0OMxWAmPhE/SE7ixRjEzJNVV13mY
rlFVRYd83BVmu5SU4Arvlaxe3uJ9yyK0q2M8EAF8tuZbX32Mt7Jc3P/IZUZJhRKj
RdZPBXl1fFmPHKVtI4cQ8oClx904xMhK/J6myK/ysxZBRlb22WtZQtqev52Imk1b
wByV2Br6CviwCVi6bI/6lNOVaefz7GezZ8VSHLcEZoFcsWjxU71PYSiQ/OuFzHGm
mQ6LwsbJPanEaJHHJIzYpGjA/rC7XsztsxYprT4Pw3iDYNRHsMblluvZArS5JibD
vaTz1SNh9A+TkvatnczYD0mylaZ+AOL0SgcT6eJ1ZrGKf/KGmMVLfnu9fR/CK85U
QHrUn7zMRn3JxjD/bDwVlXnZGAsxr5Q7J16HJtiYEXXPMKbyTdU0G+8MrPMtm0R4
G/dZvBskf5A/ywQE6u6WfCjcZh49Je8/3VY+pZ1gnpC6/vJIA40Hu+rSEBChU/tu
m8Q5WVh17YVJ38fY+mnLyWpV9X2P6uIRtBSTRp3Geq7tLL0xfn1jzq+sv9PaZ9GB
t7HcrIe0IYxn2t86jRVdNAia3+jAteRyDJXeAcKi+3AywlsOKDAq3PNRX59ofEeR
MlNYCiy9VQruovjT6tyJSDCTr9zu//p2eQYEnIF75fWXD5gCw/6Kq20GvbOyGY5Q
sckDrw96xc7c3GDBn8fgL5KP26u4WJ7gogmC1gFGHV40b4AbQ5lBzInl3d/8k0Uq
dH2mPzwtk07T54nm+xEzam6RxD9fy6SADqRzQiOcOF+TUkRwJBlsrvRVzu2s8+w5
HZWsWoIvZ+eXJf34fhiFKGqrqYWYH0RWIDHriXJOOdSsuUD4nWaG2vAoXJaOTC7F
SCNPBF1N1Tw850CCxKcRF8hTr1aabs0K+a97qaZs3/LPZ5zDysBqLiWzoe7L21Yg
ffMnTbuVxb1PEZZ9gtqK3Jel6CtPErcGpn+/Om1WC9xOhjTKTP/EJoR1WTt6vwl8
hdBKrJny573IbdN83h7qhojKauYHr4qfpXkxIedeNZbp2B9xYKnEI43a0N4P/1jT
yz/XzSYNWozg7PPu9d1ek6kM8WmMwUo3VdKwxvosROd8/zMVIGj/ioEUbtJrp7I4
sehDx8rs2/QEMNT0vraAzwxjAiP/4kJPhwsQ5SGWwlvHVoOVrwQZe3gFlpMlL6Zh
LEXPxWfYTbTPdEAwJWLu5J9qHY9lejC+03LBP6LVgxhXhzcTDPJKXK92kQWPcyPf
Ec5NUkj7PsjfqQgBAHZpnwRgWFcvWwR+jOCrdx81qjUStll8psiinnyNK/DRQmOj
jjRzLRZvEQFyztgSDeZ+rgaViyrXeEH2O7EA54+cXUfCFiCtAqJXhFQoLWm4LwgS
7ibAS3b+GzVdwSC1SLY4HNufeiBUD6W9S4VoXSmhLtD65EP+FkpPq9udz2/ddxeJ
j7elKVWvZVzWfykjdzR6fZgTV/zFn3Ak9EJZ47/SSJuSLwrR9Crdp0FVyPxbrvBc
/jCj/VNfy4ZvdCXzpN+uVbAqgLF3vmSfh9kLpjxLb0mMW0kQnEd2bVX1crUZYOcW
U0Dtlg1i0kYx27cVJcfXjEa8UvgbiyOcl3R5tcr3bYXLafCtVCh1fZLtXWuZucu5
k6wWPwiYG76dFTiyNCXpZJbe00HrWVK3yGsBxkQYTJT5478GsMeLbv4ZB3iDB/vU
aFzbqy5ssQoarjHcFldavGdFQTUcJ3o4TYswDyOQXGwlazR22dpKyPAlX5Pk+Tlq
i51kbu3xb580FVMR5DI6KjM9OVc0eN/AVo7XG+cFFse/yijpc6eJcFaAKJIsCYtC
51ZHYXZmjNP88PERNw4g0cup9zraX3QF7hyuK7KCiH2V2VPUu60LOeLXSND7OIgm
jF4ba0DtuOpaJSfknNgO/FkYTIT/z/Ce9+lpkIxwEwgLRUXlhIB50F6N9qCaJqta
6mh1eNNnIRT9YHIBIH16u6Vih7/rOU2dhGULp258Ve7nHQ2E8ET3IZlVjRAoHq4q
twZo44fD46p7DYGZ5oKuXdG5woyHrkOaexztcHGVS+q/7ClEnsSIqSnXWbMGH3UB
o688yYIf0URpApejDMT41eM2D+lVgquA9lxu+Nmi8jJMR+IDPVj00dTGDXrJEh0M
Oz+kQfieZPnoUsFfPtUMFEEBMGvtcZW7Px23pCK1qDE0Zrbm+Dx/E9T+XSAn/zii
9pa8JeeUuBaJXHfCm5zvHaisKKkw0XIYMfyzpwQPH7l6y/RpoAMmCICu03DePfvM
udnkkvOfYKrCT26Q9v2d3CUN0mlHpZS2slHRxKzwscCs1Ptm1YQmd5lqBxch3SXM
RJihNYdoLKqMV4khOH9PXN0Eniy1vu14YKGdHbJWuOxFJzdoEBgxxWhF5/VkL+G7
8Y5ocHg7VBz2kk7stB2fILIsfrWdk0rgN5uCIdLszkuVk6of0dNsuQ1/vBfmnzk2
Wi7tdInXSmaAozcbd9e6uOs/5e0623tBozfcJScHO5xj04tppHSulh9H/7PJ148k
LKrSm5s7+g6sJUnYl2ylWySkRREmxGCcqKKms9I2WDxUmhRvihwJxHd8G+Okuzj5
mBji2UXi1jqIKTtmXQk6+cEYFScN73867Uhwnn5oIK2KDa7nH1Fpj7qSpjErBivS
9Ch1uxJo63y7Lhs8XXAhV/zwNCmxmfUovuZfhXn6ZijojaDNO1Mq6iFKKgnNQlTm
u7S5byohLqiOZBK/NNUaYusT9iZUqg4GHB1rAJ4tSexb6i13jOJ2BiUZCK+8pLV3
AiR3og3roijR25jJF0pIh12x5iYUdkkPh02Hb06dXzfbzWVxnSdpaQTXFex8JGr4
8lZsDg+9UV4qmXKRE7ZNoy78pm/bLms3QavRK8bN8w1cUkon2OkZ1iULQK6ApuS3
7sp4itbvPQHBtFuiDkyLzH91JO5sRBQURYQx0RHgUelAhgheo8kaSk34KeeJ3bMn
2ecfGGJC36cqokzVrzxRnLhG8rJ6pkWXkborNFoBU0nrKBuBCxlx6e1HtwL232Tr
8Hp1YVUlqxdiHOKyPfz5lvZDWOIdicmT7AjpNwqABQzGZ+h8I+lEsJRnnoUkCjwM
JRedunXv1zXAO/ebUdiezBOFKdG0HnEKgKydso/A5gxrXuEK1bzB88e/J0YcbLBG
bkg3p5hzemgHQ+9j+ZNXWAVpw+kNggtg78OMwqtai3swKKQx06pjQw6KLTHJSDod
Hwfvoq3MVGskU0LXdjEHXGO28JyqpLN8j300YoYrApLmTq0P0Fa7iRiN/9888BeZ
EKGaSIVA8FeGWeFJInIcgqGBuiOcNrlOa2gGvRuHA4oxuSeFITil71/AiODXZVQG
VtgEGVBH7bv5cHTz0nY8lqpsczsf/Fgty6Hk9/V45tN1dBd88lvLCANYK6WoDO58
9qIN3UwGa7ZsH0IO6mfZ7xVisny7JT2sp5BpzpzYyQP3cPe0GjYrmHKs3gDKn+td
TlmgivNehl4NJpzbhg7zBPC2hFXzTv9W4CsKqAUdvPasmD5t1Ctgznu+Ng46J0dD
7p5WEmxU/ciYTzZYH9PsLzClnlflnYwe9pPznMWnadDtYt8s3UR4fFZHYxVpPrjv
Q42PLdwyJEny3iCfYjjEyo7zf/nZGhLVSW+LrzmZF+RTb9UfnvFS89i3uefu1ouR
YWxhIW58UGgaXfBjcWsHIBUs/zyaYT2zsIe0Va+N2uaqX6UGUAxjz8R4t21Jh7MU
d53VNuh6hg57MmsFOW474CnbQebIY009cvWNvLaR6jDDqhmn0S+eZuQfV+2mceq5
EGGi2dgqFM4M6BUSFKWYEiDXV8plNcBRG7S8QWVrvQghFMsnDDKuIa7bYNDWVN7J
x5SBCxfEuXTa9vmRWNbznAROU3Hk+yTMnHE7TprfvqbFBNmGZKwai5yzMgwlTjjx
ykyPSrRMdoV1Do9it7JS9AfzGBt+kCwVXyNKZn3s1GZIFDcIoreJdEbNdXw1NC/e
lsn+3sReap709DwRKLdzqTlP5DmmHvvxV3Tp2pi4/jIRMhsRdGwtQo1DTmD/gVEi
ZF7HXHAqGy2+V4qJFRfOoKRMN0fQVuodD7WAxOxTgCcYt7aN2YTDSvFyqAhnbl55
68HChK1USniXwu5gP2lzIgDD9oYDS1nFJ/p8PjQvNfHuUHD6jJj97fewWxBV+/Hg
0wLu0BTxjWdHvaUCbS5E1wcZ54p4toCy36I7TDUIrsV/Z8RJguZ6rsHl+QWomtoq
gt1EGuOdHXY92g/2f4dzA8jzbAgu77fzYEI6uyvinY22OwX54j6Z1wZm+3CGJhUl
h00UaDOMaX2po3syk8QcXfmQHKIkG2pvUw+jx8KCNgQ9+OJcfu3eejql1cbsvVLW
3gnjNvslHODIc+x0KetrbXwzNet0dO9DaLd9WhY/JjWF5aYSidldUwB9k73agR1a
raPy0Nvv5NutnON+lwVDsHz+O5g0LrcMso66scux3iM13SrqiSG6pmglR71IKX0d
cyzFN4kzLLTOUS2lVOospV28dZl6D+eVW8Zzk62/3VaxraVPwPGu1v+6BIz5hN0T
IcL6ivJhIitcW7mx3reWKFBunjcXfiDHAWolkuRSeelPinZfE5m7l5iZBAVDkbsJ
iaEB67N1LczCCHmOdDhlq0FjifSm2NiLbCMKFTRQabhAY+/cdY+WuWJXxtxVpqeu
08eSGy3C9xdYqyF99Cx9UmkhXvI1wOYw0GPBevBMOul61phw/RHb/UdnJYTWGzEX
tv7loimUtqkFDXkWeCHU1p63OgrZkSiMf5YHGHgwso5eVLBTdvkWC3Ua8HuaGL5A
dRQ/WfQqweabbQ20qg9XHhtX74Qma7W+zlhG9zHHzvqQxBXkbZcp96BNq+hOPa1+
SBKOpwi3qRn5QypaG/ogIXokQcqEJ/kLGaIhTj8F6uBXN5G6MtyUtSwo+rmaW+SS
tHQ/kZi11gmFG28ONARjSJNkGqsdcqyFoYVLh1u057rtE8xLU2J06zwJMq8mj4OA
WCJZqmRjqT7nTeGrr+qmN+qYKn1eYGmMeGJy5W1074I+V91Jk6loSn6IxcMoOXGR
jUhMHPWrl+WYKsjMOa5MaPZll8Vy6djJSeydIY1817IS0sfQdsqLQc2pm56O3h2g
Bxzq10YDc0RS7lYthPewFvwqOApTahdGM8Rmc6sXXLPNuP/4A7lAA+4TalbQvBue
wUK6bKtPa/nKoTAmlz5uMgvL5iorUx3SPQCkuyOi8s64bYq0oQkPge83wOUUQP9u
fShMvZ4uWfn0835Bbo1ARyScObDruVDG4ZggSOzignyPx0fdVBbwVO/oT6uWI0Rs
C3gxl/bNaTEGRRKvIS9HOWidpFXvebVxgnx8OCl7rjM2079OAxwPaZTstlSeMmHz
e5HlB5BtKMLsBHk7+aZtJ1RiL23VJfckI1b3gGnCGUeE0QovtZIwfZYhzFzKQLJC
2O+bVpX2qA4DrEZta3uioXjzNO4EScZm4q8WBdBnKhVQQozoN/Ayj7wNWQdY5shI
/xfx3WTVHnUgQbUr3VFAOiJ2BAnyHt1V6XBGyBqUOqaORn+wiMumsc5V68WRI0fJ
QjLRYwKdGLPSelaywgWtnw8WD8cjXOqgT+FMv0iHRBqbtdJtLuO59opxQQcix/Oj
CiX7MOYvSaxwDAtvBcBpHH65M0bmRvZSQczaKmWng0NeDCpG8pnPRKtFUEwfjWyj
AG9RX6yEHBqRODI+IZ+v6tYjurzJ8rojJchPyT/vA7io1Z1SCfuZqZAg69cSvFbu
7ijwxmpoT/DwW6Vry3PPxkPuXJDpoHvFnnfjhtI7q+DBJD48dTR6Hpoph8EzCSsC
8HHpCNyj+VhuchYHVYPjoqCV3TnBrIpNx8EYuJsFUs18Tx6g5XnKMoRBOLuFnXgX
yrCw0gNooQmVevYcUng3NoomNvFJrChLb/3TB25arNdwTvIueA5lPWVsCE4SC7pZ
NLpbsvVpp9mxlqzEIvWgGeenpXchK5z95/B8wNWz2sdaDGIsXkz2r0r5THQ0i2pJ
XP+p8MPC9q+4ocjg1CYttcVo9igfmp4tacTkn4I40QlE7pmxhqkZCi+JnBkjyXA4
hw/Vddoiiv0x5SgtPP/bGRQZC6EQuFb2yTSttnmoAJLxt9JbyYXI1HlMEzLNYNKG
T2XMWNpXkJ+Vgk4jksnQDgxbljeLLhEw4nstGXuIMfo95c1MZFEs+FJ/8b5B7f32
wvuO6/8afWQPo0ztTR4yQ5FM6J/g+IHR2ArdGuMqTXbPfBRauqMwGsgGO23vRK14
R2TJZaOrWoZwtiz79sEXxAvalVrXxPMS29a7UK7SYYURcxUS9OmktyfgFYXftQma
ktzynYM6930pHfCKIamnF+GOfUs7JZtVZyOfZnw6n/8OIHXJ8DCFnAuc7WbAy/qV
04NAvdXks0+FC30xZt57jR3qIntWW6dFYJ7vN42nJ9dk/oC3hfQCONNvHTzvEBC0
/2VFKhBBR72944HvY8N81926JK1j+eayh4fgNPlxJs/dBpqGfegswNnhsEM2pWXf
VpvBwhUQYGx/3YTOMxYZRlkb/9BAL3ADwTWyZOEI6j89U3s182rP9NIAmfwjOLMp
/uk6sQDrWLEcELUM8uK4tpZvUoHDV012h1E235Sr88Onm1DoEfdxIiX+guqugbu0
hVT6Af/uQoSr6KrtE01HRdqArNVKrmTXm4HJJ02WfiNOZdf0Aga8eTsFD22P24z5
oPjd+2o2XdCZEuO4SbKh+xKV/MmR28PlSEym27BG3vTkLnK0r1OH9JIOfeGLm2KK
44MZAUca78FPm1SolVfh9Vky8TU5G5E8PIBwH8+KSe4NP7CRoUOIrvRHeVJglLys
xBy/U1GZ2HXF2hAER/3wq/++KQgl6bJg7PwAd77Ifoq5Yg149li6F7K+mflEdpcc
lvDD2uW0tAYXtV4dHHDWvPcmyhpaCtiQZTteQQIDKawVFij418jODlPEO6d2dSK8
BBqILeiddeiYfMVHYJXUXJTwPjJ3k31HWdNCUSFVrQx3Dv5lpyuoUZbi5/hQqi0M
LzP9iU4w9COlG+amTV+NjvGQJPgasUANKplAwA236BBQ6RqkiSTCAJz9cC+1iXTQ
n+gpM5taCYvOrFFZSGxOZQ2wGo8KYXA0W5NGGXCLM+BoybIwiZbjg8KqPxADKvBV
6iOuVU2FNFImmIWw76Hyy/CgmPiPd7uml+xrnG/l3q12Bh+ktFf69PKPndMxHfRw
0jMhTb1RK6hHliEmH6kYI+Hbj0VmsyUwzvST68L+Voq4REXFC9uZZHJoSJxTzwfA
13fbfZrGJHBP9kdFbPLHDY+SPEDZ/LV7if3qf3qwl/lAtFGHl9WlewvkV+jPk52R
e6hbYKDDUHvD2luBVe0Ni0Q/pg/w6rAEuqm3uiTDNIUTLvF4OawU+0jYGTaJfEZp
IBP15I3XVA+iX8tji6ioE1NzUs5kMJvnATJCn/qd8cuQXM4CJ2F9Y+JVmBxr+4Vf
AOOVVpXOTcdI8jUZn49GYb9+7/OPfw+mwclJa0aLN1ykOzFNWMeNUYcsl6TeS5PU
Z1kkZjYpULtG7ph8Q2KMt87ReGQGNkDMQlqjIDl04DuVhbv9U/c5SWXynePAgRul
c9M+6/SprKa7DfCqr+Mwta1N5JMP+x7kI9KDnryNurAMsgOkouSy6/oMDvOV/Zb6
zjR46RLcVOKSYw7klQel1vUGP0vr7Z1S8U+oJhaLE+9MwRSrbkkFgupiXBU1uGWI
5JkJCGyjw8jVIxg/YE3NkT1SptIDa2c1snhbd+qChFrD2jabgY4CHbe+lqtNnZaM
rxOX0U4xuSAr6BfoquLWA2LBGLZbbI0Ug8HEw5gSLGY0jDwM7GZQun08p1YmMDnR
AuY5tQA58dDPJkl0Nr8/tnyyeARvWsc43lAlRgNLcUC/UvBcqxlKQBNbM+cF4R18
N3NMaPlWlgI3gV2Wj3HuVjJ80XeBMu4PFVFxCzo5t5P35uduJHOw/ragO2yhk6Gd
bvKfRigA022xvn06H6OxEWK92uZVy6dlIDuVzKRbOX32ZquimTqtjjBXZJNasHy1
9nas6jhs7Udx+CieHKvF4rvM8teKZ6zqFTvS4j7t419/E71kIJJSBTu3wEUrvaeI
7T5VvwQgI/WFaOb11OrDGiA2Qv0O3qomXlUqetEljIHGQZNCjsrMa7WuAXTZhicA
22w4Q3PnS+Gl0lccswpu/p2V5a5VpGmnqkFgW9yU9Zfme3oxyParaFJMxsDOAP/1
ZjeRKUJfDO5csFtkOGMS65TihkwV0s2qfVSIXsbTh69YEhoi1tPoWytp1QMTio2N
49VQ7sTyDfqS/QeRwhgPsw6JWzLPyhIrrWjBT/c0oMCZUIR9sfvK2iQKWBs2sqIn
MRU+8ERiK+48Fd1O2pFzS7td8s7YGAhJdWC/akzpsN1VQJl8Fcquv5RT/gyo5upC
f2M31XiMQmsV15xdQ95qOpbqZ821xPsJAQsrR/zbfZmeqb2rAmF49Ai5GywQL98T
EJ+XTaMkcfiBA+kDQY5U1ks0Lux7OH/hXJV1cTWsC1LOr5ZEMMAy8r7qJjSBzwOD
DzTZH51/9qLNqtAefCxhize3U2K1sT99LE4FKlqet84krYV6L6z9QsV+ZxiqBIos
JapPzwOo8ErqTuduz2EZHWjgpUQxXILjgUSxPE1SH52cFwGeoO8pmRVuFfpjgQob
y4FuYspDAA9LOnW9EU6jAVtlern6TvWpuFLWKCyV3+mzXmgbn5eYLHP11C9XDJy1
qGY5NYhHsdOEuPq1PNG6wwVWwYxvpiuICBR2hqr5FyP0loYwm/jtZHGTUekUXlLv
YVfESEEJQb9I2cKkmutqpHvkzAP4EOq9IS5ZVF4EDlni6bg43xy/5ZYYFnY8qfo9
30HHvOXvdP/w/yeTH1XRhSN6WwFZLmEFQpY152un1L9YAcrGv+s8ExGvD5ddmyK7
fdV+ldLw8h1t4EwhURCtep39kD+jtnQjK2qERs9rW6RgOo7OQ17R1EEGhYImU91V
Z6yQLHIuLmfqT48KvDqmXrQg7nmzRcJB7270FjIhZ9Uvy/taaA2QqwILeOoFli3a
3DGgChfddh1rFlCpBtCoIV7k8YYzEUwY4oxkv1KITC5f8NHdcSqLJq8i1CgMisVH
H0nx+cvRmEcq3gLOCAjirVla3PwaxkLMrJKKwHJoX2DkVPtCEjJwaCoEvRHOhDKD
R/sTsD4+0pI+AgnWk+axBpE4ImQt5KCKbiUmPwDgkCjVWBO7ngmVdzX7EvtPGPmF
UqdEW3LTULuX2u1RsjxiLHJHhEiT33Z3JiFkoHOXmj/Ik0IAl2+dGkTh0SJJLWfz
+B4WiH0JA1ziS1+hzDWigGxQlxYdtDTjWA33Bl9c3zbQLnD/P9SYwtFXFzMYgIwv
DGZdZQJ0BSxfi/AfUy0b8K8gccTVqqFUUd9rP5Zs/gWSnjbKtvfI2AGEBFThlaVB
HCVZGAjgGsEstXFJEMktBykSaj2KnT6/BGjlNZBWPmIu7KYseQUOzUtfoNLTl2F6
f8UcvhtZ6mugbMXS99LlciI9ZoMmZ5PxRPVrOPY+yHW8WxgoQF2Mzyyhe9PKeDBv
zMn+T9SpTnZgLIlgnDvviJ44+uMyb3YwFZhVvFgb31Mty+f7zsDy3RqRd/oK8VJl
QISgZeDdZCTqDbuQRUMu53oubYZ5ZEphZgEL0ZGUkZjbwAvmdEbki0NqMt+8hUPm
iQGiokdSYbNh25Q3n/yklUpb6JRT2aX/QKSOdimQoD58lDZu8GbPPkqPpPfSYFJf
WmutE3PODhAjUJ34hfXFSj6IbBgq5iZCCdzQbSxmCsRAreg8MKpQ20DxqkVLwpKX
0oo5S4w8UBvFYGZmvmrlX8obQwFt25NCRMVDZaf+ifbREBuJOmhAB/v3TPlmr7vB
/gHrrAviRiUqkFSySNQ+t9/Omct8FOB3PunoPw++YVvj7G3qFoNhLGGqPtxkhlI4
yry7gBbk6k1R1L2axk913S9+ZSTqg8MvDvYh5LUxn+BkM1Cc3Jopz8v0Ku8amJ2n
6ABEMFiyFX5IP29TUVEYCcXNJK2yojfhlefgtcSAOITZ0IjKaSagjjQwGlVWSuch
qrghOmEpptqeh+uLNtpIGVgBO05GoXqYFjzhZTbkay9RvKqLHkjRz2LXyk+onCQL
qnTsqjc69n4itUP5p4l5GboKHE0XTx35j1/xhiSCQIZGH/zgePMZDyD5VIZV6pnd
De13PYPWmb8RJ5AJCI0QQPkc5xml+9w7Qdevu/SJLldewteTyftTWlcbGsGuUMd9
W/4KQnYp1qmvyQtNgW08fy72x43lCkqng6od5cfJZt+ww761mcF3q258DifKgo+j
h1BWSgNrsAPIjVgds+MuHOyCqBadTGJsMW0sbLCj4XtGQfunRLCIMv2IJc3ZcsA/
1GdrIaDK9CUplp3d+1N69ZzVImPL1oMOeGcoN/Q7yquFbRmH55KIr10SlmapDz78
CHIQSqaBwgVuiSkuT4IsENVFBUR7dZWcgUqRSuB4MurGUiMCDq5YoHyaN/1Z/EZZ
f3QrTIh+ULzXiWNCd10K7uZBn9znzrC+mvXQ38HQ5eRaE1iWGrAWh4FM6/jptMdR
P+6x322oV8hzQfDjciVSF/2Zo/sTdisVhhUTn6qo7ZIJSBPjgkHutjkl+g7nIY3C
aKiLs3KXeoS8UzunKs1RGN8plbmgE9JeohooTm1XpGHN+cA45C6M3PT8suRt547l
XhKJjgnmEARVhOpg2E2Bczpjgg9n3hxpkDF29LrompMrAwB1ZMuZt2UW8ppFNyjY
if5nbZkBixs4l7+6YY4rexJ2Nv9pWmvPKAK16/4sSmtTsNLMsLCgXZwx7zHyHx/l
smpwxgx+cfXwRmcwnH2jqkNXZ47tuG5MP6yb3F6pvp6KKeDFK4mlfFp5EO0iodCN
T5D+ECR7gAg4PoZFI5vpfAKjTFWOmtnXi3176W370oRjsK+c9TwcyPZcPlLNnMDo
HO14hDROc5oM+A56bYKcRO25zsblRTPhG48tN0vsisHQYyIsvfMJa29hH56FIqYv
wgf2APlPFHaNo1AGrYP25hi0kYrLr1iLTqofZoY6A/Jy6okgVXKL7OV9eSRT3YTb
/i5JPkO+uovl0WRzCHUTQ6C6zsgxaQ0eBKPuY9MGGejweAQeG3ATjL1JO3240dQc
P1m0f+nEz/nQu6XRtp+NtFE/Yrspc6JiSfVEAB5iiPqHwahHWM0g6TrTsHCSnqJ9
HygU3BnL6gFWcWd9k9LBV2RZW9wqpgwAa8WhMJSCI9nUCwC8Mmxs58ASKaC0OouP
p+h2FTt7ZxQL4yUP534GkaMEVcFUtY81vnbxD/Ps7qF1tgawQ282WK5/eUQMggtK
7TxjfPHNPYFmnIehqYc9a4GuvjazI1AE3QAVlHLLmFuj0LYcpXeKau5Zpq8MDYfv
Ih4dQFjiUo7KUWXJe9aHf8pNiQavH4B+B5YadC9lJGCac+qfGL/UdWkOR1/dXVZF
8eAmQunsB+U3O2kByDRyY8A7pBstUXT9tsga7UZiotm04xprOVEG8l0kGUTm+gsH
2RtIdUs+fxv9ONb+S7JgCYKKwv3Y98akaT/K2pZZlAnnuAYWmbdjAYboDgQSnIsR
CO56oEysslAm2Dy8nyPvD1jYy7JMe/XGq3OJbDjmNVlJ81igzmc+9ij2o7qleM0K
1SLNtNBzzivQ9xgRsIPFzfMQnG+YC4R8HUglAO9o8LgPu5EwfwtIdhtaccXPwyQz
3QX2d2Arhuo5gPo/KjQWPwImr1X+/sjkz9fQd2+MZ1xCM4+pLj9lo0zRfB5Vz5s/
+jgweBQvAUhvEGKWfO4sjsZAcjeZ/E+2cJhUNPegdysq9u77o8PPu+1U3TnjlQgn
bdZCp/2Sv51tjGnURJ6HtzAJ6DJCTvExzqij1X+Q5jR+TGCGLfH6QgHszcX0QRgV
2HNPGUrXlhzrfdnE2bevdHFWNTPCAVHpY77pXsbeX8caCsCf015LATOipFRc5V7P
ZFdGDBbgm10ZB34Nfek16Ns1CV/dz6ubU8u0JG9whH9JbhFzW6uSPVKcEr+Dln6e
6sNwYf18dSuxcpcJEp+jz2vX8kWmjdNTmn53gtLz8Q3JKKS9Jcb1BQuL6lmvwUjc
eG6vPLjPmsGHtJnZzg8eGHg29xxJ2LGEouNLP9lhR2EoN6fjnzYXE3m1ku+PbTJa
P/YusWV3TIcGBPosQUasKkIMWC3C0xVF+oDJYESdaHhSduiLkenh9qewPjD5CnID
ZY/gUUaOg2CWIFUHw7LDOJlQrUhR8BZmsS2OvB7zc6EajNmWhsgtc3+VV4/hjo9+
P9ivLT1OaZHGNl5Z6u7x9sJ8ANYoAyYzEhODGYUc1cBv6zU/MaO2kMQk9UWaUL95
MuaM5OGcyzX/Pkydy3GbgtPEWrVpXJ1drt5uGuRSAqgGZs/dyQumsD1FzPsH2Wn8
DAlbV94CLOk2eYMhlxH0ltQ+Lyy3mNjT7loLy8toVnsBUhRLjVLeKWLQ9a6CFo7m
Ea8xtl8ofjGWu7e49u7KCSxAs72y7ZGFGgtcaVDr2tvcrGGWZJE9YLSCDG0AEI+N
/hUST37DUHnVlwap2EXKuog9/7Qhwy1DgOz1F89NlqqyDGvUBUGtu+F1vzXSC68E
jTbFkGtvl+DQavR88KTYcQaHqgcS/Nj/J3anaFfOjNWkYUlS13em2mThU3zgvhNW
pkCwC93j6Xt6YAWWmGvaX+azZxNyH0ss9aqvMAZ5ZEMLUOwf+SuO4g+y/CRU7rS1
zgPBvJ6s1F6MXFf3xvQhKB53V3jmM/uMvEAZXqKndFZOfFUY/ZvlTUAhbez82Hoe
wAZqMJKxg0abQAt6GPIep9zwptqctu3huDBxcwB3U+WgFLUypF/E0TC55sOSQJo/
z2MecPDFG6g5U0TvfWxQpRWajQ2rhWc6lLblCF6oJupRP9LuvHgbFUVSbFBnnnug
aqcpT9UIwLHWImkoGMyCIntaFFAI2qUPqwpGcZ1WoUdYfW+SDN+zIW5euGMvlE2a
H74xTEFqKf3F2tB1K6JJhOb1fVr5s6u/WdTmi+EjDlhOcEAtym/NoFGJO48NPpwt
UbaHS6QkOdhY9/1HEeHgYgquPuh//JXKrSzUGqtEnWUdPqmt0N+qnwdBHcTcf8CS
FHsSR+sfqi1jSA7BJHos2NXmHnvPgIqKoc5zyhwAo5lidesdPZ6RH06nm6HprDKe
8qLWsd1wZJDQ2DdbM9ZEZgxlzSTR9fe35hPj1JvsN6S3U+2bGZZ3Fb7EJPldOYJa
crno4fKV26EheaZi1XSCImOrEoCXtVSJmVUkuz19U6WHXptRbrTkkZ6v+lAQ7gW/
p4aZd6OIcWWWPhiqztE8Tkbi13J1a1AFBDYs8NMVSA5lkSUZnUlzttTYhOvpG12O
AdmNmgQoOD8P528S99k77nip0UIIn20EL3G/WXJcWWlXlHvnHr54B5URtHNNtxU9
E26LsR823xX13HRMWYPBJ6/P9kXnn7nYt2nmJzjmtjApwpw46tcF20heoRhHropl
Dpl7+irRPyCzSn1OEGCvPVLaBFlxf67DlQQ1Pl3oB8VyzlqpSRKNuK84XcfTVm3+
gJmHtA3zUVAizCGyrFqzOTty+gA3UVt86L4H3A37iOWYUsNp9B9g+ZluaWfTEsS2
Cg/DIpMV9qQVuPvq6QFgxFnPur6fr9sfByBDZZAmyaBMnZ3Z8t53khOmoI+DIYKM
L5t+Q4yXMNhhsPVOYfzlXOSwG7wwuHoZMhFp8BlP6C8Ave1j/J5e4k7Zeph8DF3p
GMA37uCx9Xc+fhRfX2sTXNL8P5JHCnGjG2WgFZqefKF6DLbwaUOsf8aPwQr29RIJ
ZWOwJirKeC8us+k6MKuMtl7XnVZa+tWXLKGb3WwzR9XFLYnwz7H/8/TPYhlrPDt3
0DwzLqDjGhrLaI0ICUyYsl635STIXI0sjodbccvUKUePXa7e8Jl28+L5+xWaMtE4
2O7Z5ePV1UU//aqNQ43IaTOsSjLRFl2zdeB8xw2RhzoknXD+261gpjotVAceBhj9
zvKAXdCn2b75QFtQ17G5NftQcOja6gegXrqqG48VRbFCmZTVaLVmwv2Whs16RfLb
e0r9pe6NY6t+oEs3m7L8jzxpfD+vv5eZBmY+2+KTxtTFghIZIt9QsAF0GGlQAwjs
rNoLS9nIHerUeg6WSRJIBNBuPeNCbfWT43lH1aeRNTZYFHjOC5ce0rbEB85z66GG
3a4cIRsAk+3sLBA6TIDKdXePMEGT1gYs7uBiMSJXLXxx8CxRRgwUPzAt4h0ZJGqU
Ggf2SXczQG64lzvLr0x0D/fmSU5G4sEB/UCz1YMIuorYO1hlAB55isfbF3iUUBK7
tfLtqVZ6E8vEAwb6sYlyz2ZtIsbW6eyfprWbV7ShQO1lteG50B1gjsn194lsZxC3
bf6ZyjSzYc2dyMNfjY7yFLXy9wOAjDL3O8IUJR5fBXwFBlMr2Hh4jzJCPirppTyg
cstjeVffSzqjTwndTFLB3A1ZudMO7mUmmP7kmac61o7wOD+bHfijhKbbku1ZI8mW
ZXfYxYcGOqTDwk6Tm8SJTvj6Fz3PoOaaFbqI1+Kfb0ERGY9gPlgAkGiZGbby7n+m
5kGBUB3QkJwXiuDzWnJQ9KtcZI/9RgEBenYzweYjHLQziZ4k3Ofp4xR56aORZFGN
leoXBkOFo+hntWoixSm1hdD3+fwFlFLjR3YD7eUrN3p4M6UQ6oBIMMAC38pDr8ZY
nov0necpxqYgAu87XibB5hQHtl1umONOqNLnxm1o2F5fUf8t2Sjuq44fOaH5blfC
jZ9KwNpZsojqZZNZTNZC0O17/2ww2G5pwtcoW4ckmZgqkMP886T4CnarlgdBx29U
bC18fRzlEWlqp6U81ym5nqouZLpxB7Zjc7oWlM1A/WGm85ERZOYJRAe3hf/DNo4T
/aCq57mb60Fufl+JBy+2EAEN8p6m64hrvw+5uZJ+K3M/3kLp/f71L+Laq8UBqHOC
HBibRnYFAsFZPsplwWsbLaGIMVb+HRrlwUoVmezF7rhFByMO9S7SSy7pESiXQEBY
5RI/FnFMIajR0s1R6rQErLw84AXTBy56P4JeHohK5o/fw6o/tiK0Rv4cacgQIdKZ
luuYfvr7J0fsDH4RHL4IBfjeAhWn8j86VUifBrNI57N8zV4StMadbnOB+T9EmF9r
8hqV3f8/bCHl8ADF6P2nkwcmHKmCZRZVsjB7Y3NKcszzayldtxxM0GcJ+Zpci/Pe
hNoD4aZeGCIcY9UJkPq9q0FS4w8jUWgKvCWENAPzOU8B0fC1LPl5YtWkWyZ7pSsZ
RKda+rUPdeYUg1X8ZjUDPIPs5lym25hR/h/xlN1ZLlbYjLTcFhc8nI8OtqkBY8Gt
AuMw7tjR7nuji7RKKGPODUFgFQVezD+i5w2dFu6dH4eMBNnDMie4pvJgR3g5iNg1
mI2Hietiu/qnPk6mnlBqiUdf9IbV9vclyrBEGYbxkkom0riikhEGUwDMkZcVQdgS
+gJ52j88NdJfESI6HxlE2eZ+5O03WTC0sCQMHjdYuCHStSahXaaIugZNoBCl0xOo
NAjgy46900Sh7n0T4BUCCRCqJA9AmGM2imIsnZGQs7oeoo134F63U1CiHAsSnSQh
//osn1oJoVlGiQSDKZ/gtEHPNStEW+H32IHaklMlr3TD6jfatRyH/kI47fx8B/7S
nESkQv4F/aWGpblflxhiZYTSt0vOwU47PCuEjdH4GXLAq0fBKYuYKLV6XgsM+w89
BzrVvM6x0iB4diK5N9kykKS98zYd0UoiYJlXRDrWvlhTMxiLP5aPEdv8qlMNdzRx
RrCvKPDoFDkMHAmQmhdLqpEPZ2JdCYyhS5b0cvbEd260sZVd8hBXxoAdH9hwV3q3
sKYcYTYIoPnuOY6wJjo6vc1JCTFSwDo61Qz2CDvwAwoP9Zx0+VETXUxFFP/1lcPW
svmPcSkHCOs8i3vo4F6Me+E6UN9s7Jffb1CQu8IWf75UnJGR2NR+9TwZOSfu4Tl/
Ayy7clFGfdH0wgrkfr3naCXCzvkaADde5FIeyrXH0YNmxbQzFA8DwbLCkJ/3oCJ6
yfxV8SIU0hJ3P7rG4C1BlK030ZfZYuOzYOfx07H/9hvUlnlOj2fkYhJWLGX3lcO9
+8lr3k0g5FigWCXLD8GJzK6xZBjSTT3Ttrv/XgffAIKjibkLJE7h4Si+LZurr302
nIivBrkFfA1roj31ipZczr8nK0q/9ob5330Ne2IBu/Y3nU60UzwGFXdHMflF1/8Y
qnwBwet4LkdPTgg8W+/O5kbAL4mOdoyg2pjW4IKNm+wn7YHP1T82qxO04sH1IeDy
VznebsYavSkBuE/JDhSyIBs0E75wSE4pRiFTkgjg9AUMRc37H5ybmmt6AlQW1pYa
IkRaPnVlg4aYYDH0CU+5Ck7CXDWECbRegMaSTi8rkM2K9YhqrzigNymLtroBXPDl
9WQ8IBuHWbJC+xpe9TAbitX767nVHuVlSQ2/wThr6dZ0nv0a1WcQiR2k+OuSklBq
nks0IpqSXN+HFQBMusZcdOX6JEuvKLnsqA6AqZ1cYAbJoMEkcW/y3jhodwewMzAl
/8wnUJgXEzG8n8Xc65TwBf3U+HQEAbWlx5gV2mX+2eADXzuHidRyd1V3eURRX3o6
C+2mcXPEvoZ/WQGR7Qh8WgF2jg7OieV+Va8KYLuXx/QCUDMtz4QdGf1YZiKbFVIF
gbMzAlKuQoCB97nRN1TpXzTZS3rrnYQebEqPh/j6LrY7tiESQAlts/ZUDmGgHlZV
a02ISox5FlNxD588J/qilH8p143U1VARb1ia81w/PBL3AV4HVq6H4ysP04CV125g
v/hv/a57QGZnJtVE15ckwaXUyc1g8RG3SuY2COmOJ1mowfvmrUIw6cQn7irXX8Pg
x8nMXFaqN3zgX7eygikjhZP6tC35wmSB4pjA0RjsLLsOFIhrk42rnjPvI6KpQY8s
StJ1fuvYhW+nYImUId02x6buZqYdKWZKwPK4lFizAjUfW4wEkfA9m19y4xtTkR8v
ebDDV9EEZCwdOM314OIWqerk7B4/fEv9+EgL4fGAjokGb5EO20NpVJorYSVzcceh
RUn1B9xL1QyDx+Mz60ZXFp9akeDWLUjwv7hSkO6siZpe+eirlxYuSgFd/vbDZyXU
huRyLHo8lH+S37YAFtg2oZXAjAJw6BGeBAcu+AlK039EdleAtRPhuxF+KTiLbt/9
QxveB2Mz9O71u3dHd2JD+d5IfDR5mV1WwvN10bqg9nfXGFEMBwOdHjkJR3OF3VRJ
ISkLgT/0WkBJSg6dbk+vYnYqbiB+kR+9GA7W//lr7vQGKEaVuACYraA8LAFAj2gd
973UiHM4e3kAjJTaHGQiJalUPcGOfmEb+vVkx7q5RJxpE0GP2jBh/bPHWkyRWCNU
CcdJADF6I4jBX5h/mkDhddgR/FxsXex/kHShHhlfZTH1ahrIFr+yxMW1va1T1LXe
urPQLPRGIV6otGS4Ha1z+Re+Xc+jlAnyMLyClFL4oRJROdTRF9uk1DiOLoF2oZGd
UsVFlrNXeh2Xy/7flyvA438HuXIjVmYcFL2pN8K1vsl8NROW4zgb5sfDgUzjrpjm
7O8NJuZV1kogSAy3OBzwmDUtjSLEDXHt379jcesx/nvsD2f3CLJYxiE/+e3saiAc
jl9Ayiq90OSDLHML0kBtx7HhfFF/aHtGnKPZYy2DYJ6KlNkZj9Pcm7z6EC9yh3xa
yvsN1VgfO2nTiVGsn8HQkyi9xoRn8FUjSWaLvsEQO/J0BQBakVnEgBiTiPMy2KP2
xIi9FzQPTL7fBml7osbeGoY6jFMZwYY12B9BproI+ewwcr1K0iZx4o+/RmcmAskz
Sf/8KPHiU2sjq9OG+VjFh9GPS5V9gebf2HyFz61wOTT9Um633ByJNnXRpulr2EPo
c9vxST3gWcAypFrGdTIg8wTPdLWdKyLq8E4Bp/xuzTNh6uMK6/8nJyLkUuT6QGh6
WWFZfKlYp13YQU1Kn0kvehx7ggydOGtcrv3JEBvLUcYHFFu8yLrxLy/sibg6mqjm
gKJjZS2SgCnK/edW4TGVWBJLpmoDocpH0WLxT78wIB0kGytNc4RQRwdeGjq36uE9
BTkc5pZ4IRKqnBVeXdZH3goc7W71fsBlm/45eGxW+TGYA/mVVgajn1V4oaXfEpQ/
jA/dmJcIqhK83dtCBQWbLtmTojHdmHLRWFVb1J3XAbE42NDDp6P+svCMkB3tVcvh
GEs0uMWSO65NhKWwRK2Z4Ohr8l/rg3k3YlXxK0rAr+1zQe9nWM3CstzfgJusOZSX
499iVmZuZ23vmyah80SCzozWl2wPpd0tOlCiKDZsCo/eiGzqahBFklUD1RqMYSaq
eIDh4RO950641JSuT4LQjJHOJ6y48Dn4KoIb0/sVhv2h7H5zJiIjU99BjB8F8Qb0
WYDQld/oALiY7l1ZxRV/7HNoJQi1c5ddSS9j60DBoznLU10Aaaky97rct5BgaNJy
+GUevGr1QzfIUXYY4L0xtDT51fQDeEpLuO2Px074DB6h8m4dLQSB+VMDtfpFEjzO
Da4KFJm4zn5yR0iExWt8EuoIygC6QbVCP9FuLmiJdKzBWpa3ydCFsImZjL3P7c5f
1n50jv9doALtMidnv+Rq6rooeaR6uh3Xn5zlk0pNj3V4+mnaK2iVzejoDLavRvOx
Xswr+rh5wjvd6/5c9ryATlfSwanydniggGcYt3k5RxlExybRhE04GEiT9oA/7v0D
oi4HwKaQdGUZDBVBfBSNbfJd9EmIWxwiUTMMBTgvWeS3vHEA653TPC9KcP8YleD0
MfAq2ZGBZ0RkVaiyTZO4ZF5Rt8SFGGD7XVfIUzr5bKkkmMDEn57Gb9KV2DZF/PAg
+By6mwe2pqGsUy2bra4g6mk9a5juTKNYMdrqkXPTleQIP8TecO91d+vrr0FuBDjK
EGDoPXi4pljxhLNC9A2HLCGEai0wgf7K+I+4kfd0DSP62/QZiK9urz7v0DmCJTVW
vk7V4RZm7xymXmPME7i12TO+Tp9dCd5QErKQ0NbS6YSN2Z+JhUexDTJaFP7frGJG
bfKIN2aYwkSyYFifkdlApvIs/WoDBSjZ/4UPgzUk+xfNK2xxJQ9aqxELEvvsUzFM
UmhoftceK7kuPBOB6o8ug02smhPzN7s0adZGdQU7JAEKXP4w14KCTYWIohkXCuLP
Hj5X7vmdMLRUPpaMT6sRAMElCFqgm43NdigkJh9LLtwnONSW9NmFCPynFQ4nc0W0
u0oJZxhWvt/qTkajbNuQSBgb9zOsMcnG0vy6oJZe/L26MBZJnEYguMbXXhfm0Qv1
LkuM74z47/is/+HnWmLxLrdKpLhYisbsKICJ4LV28NjSzZM/Y5DN/R59SMXJVREF
Hc4lsxI0UNlz3dxom4wjCq4mUj+hvXG7GQ/Eyq7hdfSsA9I4Xu6c6Jmu7qNvPh7a
z5bI+oD1Tfks8bJBBXf0m4oIBZ7KsqTM9jvF7r8g7ZL/02pKQdTkIUsQkozX95os
Mkzs7lQhBQ+AnzSeUHpq/2gRkhDSZyhRSOPBkfJe/EiiwcnDc/cY2QGYWQZqYUbU
qN6lD3YxS1hXZqgqEKXXEIdR/imx0Oq8XhPnhx9jpQ3njGpdAxOEbEXOBPQ9w325
rtLxhMo/KGJv4sPm4tMGMyyBULk3DDyKbeZDv4Ey8qM914/JPoQ/TLNVr7sfRCWM
A7WPTNd1dmvmERHlPmPJ8bRMIHusncnuMA5qhHr3akWF4U6qoIAhUFg9XuAFJd4K
AU5uaALASvKMnvtf9vuxRhh1tm1su6UrIjkYPp8m1Z7NRGCmaUrCHD3HrExrh1+k
9mWHquOjShje3XXlXDJi4uwPpditD4DG43KjmfeN29dCtx5XOKUIuCCu5ADgB8m6
nZzJagK7XLTfHOF3ioE6lhe24DAPwRXib3ffcdje8LU+FFuWf5w3hxkQoYINLPE7
2x7egs5gtftlL3t0SXcGfS0h7R/9ODanQIWFKLGo9HlTjRMtJH17ZZExTuEQk4c8
SPCUMufuqQXkJq/lzUAQWBPxgS/zWXiHOWpxzxMRArzeSxsqqH9xyny2eB6UGs+B
J6h1qMBzF7wDLjZoXiMkh7C++bj+OLWyrVlaEbDOqQeSY4TL1SQCjRcJtPGQu78y
OnMYy7JwYZU30fSz+IXUODasyMsu6BWzUjB0cIcOUT/dpMhm2n9NTmG5mKQq7xXG
a8WX4HG1GcFejQS5Mv8Rcx3uTPowwVEP3tUa7lHQu0EXCIwOpx1kuUllynJENDQq
tNc2F5SUJRgcVOA8zyFqRTS0zYlsieSt7PF4LJNOJ7XR0Yo4CReNxjPjjBFZDmwV
hFzuSNeM08USKsmujCYtteotRdBcufWSLfMQK0qoh8wMclKcVcWXnFXi+jXcra7J
+dwKdU4Aie9/tOucXgyD8IPq7LSaCINjKtzbXqj7dk19U/JnrrFOqP0a9q5l8CbW
kgPka9BU/g6pWrJHnNk9FdlcKQ+ZmKxrf0CcQbO7cV6Gl20xVfD1f7MThtjzzpJw
M4z3i7SgLMbp/o3nGwxnl74MWWVdlP7d7JMqhfkFrKwVMnRIGFRRCkK90o9OqCo1
5FoTN5X2x+1WRcjRH1ia7iH+B3q7zrkU+j1xnsBqyGnBJbDbxkQM2keugj0n49cf
K76oObuJXdqEh1CBV3HKF4ueOvtITjeVZ1n4b0sfIao8iEWz4QPeHkjr/iyakUU5
w+Y5oBnyzSrj7WohzsikUNpBFeg6qVbXCummWh6LZKxkTR4GtUtDrHIT9GzmS0O0
KkZpODcaZ1EX5H+vqmzaqm/4BrnUitWl0u8CAUYr+NIsEB/RBj8E1WfWLi713sD/
+04CLmJL58BHsP7mJELvYYcs7CytadPIV0ITj56HJJ37JEv6N58l8Lc7vDu+jVTJ
k4sVSD8QREMa/b4QpVVORSfAuqWtVI8Y8JnlWK9c1VJgl0fLHtQDYhjHyOPvvBW3
6N+iuizyuY5nkr2qmnuSDkWvxvS3MDopQ189OmZEtn3S7i+bhOvgbGxVJWwxCLeD
xdtaAjY6rlTHzqltxlYwK7HcOxwwK7cYdqiRJlwap6QYn6n15Xidj3CM8Pb6VXq5
nU+Ej3BDnQMOt1gHwapn/exKjkVIzlZzzhrqu/zpYJ6e8pyegrSU19YiEs3QSJCK
/KLvN8XOtoh+IKPC14OxLGmsNMQ5rZi474D5Wy2wOA0x9om6AG/V2AcA4OCv+Tn0
pjfruF+drMABk8rV/6PMRRjy8uBnfq1vgvtv5xBANgMe2jdS3O0zYHBpVJgTv8kP
OFMnTIpKCQD3pWlv/5of5AD14OZdptyQtDyQxx+YuL8il/JdJVwRAheJntob0KB7
zlGEhGC28wMRhTY0nWnC/RO/2cn9gB/V3ANdy9naYnnv2Taj1Bmnk5npjaBE6N6G
pDQwKD9kEs7Mq4y6N5iQiwqmheaF9jGkUi4sstC2eVO3Nq5efFrHdHWx9RrJeuN7
5Qjef8i1V1JWnLXnhoVa0h2f1YNzLR8b5F+hl8ur7o2hbVTKeI+SBKVcydAf06oF
7kJIXop9iq+zlkRUEyALjmg7CnpQD72joStmWsOGmP5NVpBcOAlZbZKPT4eSbyb7
U304k54ypAm1Ya62Nbo1cFAHvg030cNNdtdiMNsMtXnpsK6PWLiiYnT1irLyf111
yjQSqQjpWDIw1kL9UDccBS7JjRPzSaQVq81cGsQVAB8tOK7MzkJEPn9t0AVv2XyE
huRlwkD8T1EAMC4ok5JPhUOdTRlaMWrZAh5uWkUWk/x7Jn/uekk+YUPbJ/+S9NMe
UZFbiR0KQKn9Gy8qOzUFb0wk/f93B/0r/2rx/g9p69xraZ49OvUgraSbBvY0ORs4
NndMvLvY6jEGCs3eC4cTIfspu7P7nazICynkM6g3wdFt6lYcqLTcayGYOG7422LR
JVIK+dq91iTC2pMGb11qrUEg3VkdVApIg9nTI9/+qzqbTiOFdUCcJWnZplIXdXnj
jK4SJwBhGGK4xh45ZJTPxg9M4YxybGcxbo3kkQJ4wPk2R8unURlLJVN/0PCdFC4n
y715yay2MmFHfrwi4MZWUUsHZTab5dEzJSoXIIs9fnaOPOlPpvgico2onvxvvwxi
Hhwumhg7nqDmON/u8bTqzZHHCPnd/lzbBjqNIUwh1SMw4RSkQU0VePkejDkW8ui0
Pr81Jr/rXpnzUrRqJdK5zNSFXcmm0Ve3bPgKE1kNXZ8QN9kOFhv+fClNuX19alG1
UY47GayUJWNOK7eISHr3ccfS0eWpehspVN434kGc9ahbopZiKgrcK1qlxrBDvxQD
uAO9UcN9ofJ7G4f+H+9opFDlkZyi7yEGqqYv9fkgO7eL/R/xzg0o5iPAUF2fv08x
cy2WfOo6IKgpeQLhrLwuxNLb1HemIwfkD5rt7PokS63O61wy0NrunmD/Bwabvnep
0ozHAenFV6Mq18g/Cr13U6j1caTutsvDCGcIjXTPEfvqr01Fl9YEZfLmhyJoDrMy
JRwZbYD6NV6xYbmNEJ0IXNnLj4+QYty9rWVAZR7xVX4IO6RXaXF7CPmL51Hex9SD
vrTW9EkcxBTp9lnq3ZSjJXfechVptw+Iwd5WeBP80tgW3CmP44yliReKj7s+k1g3
pneKKg52+UKvO47dAfEaPYN7BN8huBu25q0Ijd7zPhKoIcyzf5LWMWc4z0k0rZAg
NJcz/WQhn1fGJbvkLXxupTnBPF1W2tTmxuCDxblPHeh6+vTn2mHkTg/fwHRh4SSV
gJnYoZM8MDRHwP2k5bzGsduUIsu3/+NXyWuuHSmmg2I/Ce79zl6+iJTVqHoyzRfh
LYkj4Up2FBampuTgwX9ptfm1Z1MRW/oVbW6UBubl1E3RaE4TlHK0w4nu/L8jnAlW
gzcqe677FaKHtfslyWQDJQzFHwYu78vi3FwAUZ6GCslbY8wNu7yZg8v3XaPADv2v
H2fFaKR0dOj0I8Q5xY7VRmZqPtDNSUwQNREG/ynz2Rq1vDrFurKqZ7CymtI/8jDi
TtNo5uAPaPKloZiZJMwaCeDZiFRIFBHDq0qkvTaax8MuVet3FlDeDZPMgKRjCaeB
JCo/o3VGKLOarUFee35hUdI/Kc0jNXR57sWeR4cTU0ipt+uKE2p5V3xhQ+PqfqDe
iK0Hfz8SNc0K3R+wQ06OHcuPctRVjz8g/2FTjnSOuV9d27w/a1xbChQ279FVNG++
ZXaAHBZUgIvo739WjJSxihIcZVO3fS6p54hb2d4C1f6zI9+veSJAC+7lk2HGGJjK
tjplqDiy0XoBxLw/nEx40L2+hEZWqE08JJiNU/PW9/tM8GvjAgpD17beLi9CpcKF
qdnhakRz5sBwQyVBfXAUwPrGnKL0xidMD2biEWgTO00lbvgPDdPE9VgsJXYcucOn
wSiRzj73RZCsYPS856IUFgJN1d4ZSnbfhRZBuPUFWomoL1CRACJMVSuHZ28gVn2g
D1QY6TzdAUaHrktFHF37EbuNbuQLIVk1ZwqblUgBHlTprzPZoYz4Pky5BxBZ2a/5
VePbzxQ7WK9cMC/1h453yAXTindLUkiVJtgCy7p+IhHLtMXu3T2EDp47CBMicKXd
EJ2ey3NkhTmHwXHa4oXJySGSCq76c8rXveoGwgPg1jtHs7OaSGbOJVMd4bBL5Y+J
DUNgry6N3pieJXroLPA5GqJ5cjhBxjRE7HxJr/rR06BYAaanVnTnM/oIi2qJpKiC
w5fslAHQ8uN79tccDuPr3bKwIVP0TFMQBt/ECAwLyb0Z4oR9M1sFwX5uwU7hvcgP
+Rr2/qR2SjzVrS4EyQYVS5KupGv/fJ7hGrsCelgUTX63w83Diwf6rsuJa15Fgg9o
Dt0C+33LNoqDUGgps2ywIFl2hQWcPTzI8wEIu9hGwosQGu3rmHtXDOduYLV/iAcH
WPzEXdnRr31hwbnuzXwUDPnvQb2WG9RpX93z40M4FDzpnrxWt9XtPTlZzBoE2vA+
oTKEjAhFCga3twcSUpLZOzuFUWKv7SxgA3ERRV4kElBrn12q0DtEHoBOydTqxmkJ
r4Kyr3BvtN5UbOZIAmasmRKAxQa14aQxdWYpKfSKXj6nDF2MvIxwghqB3JUS/Lw5
7I9pdpyfGazC8424uM8jgJtX3tRID2AJZocf8nMGkdkRpe5qSJwYH+sKLa35oXoY
/U8I4LgFRKGWxKwEbxrMCkvqdSxR51PwdkNJt8BQ7kn6X4oE3rGUgG/k2qhQN6r1
KN5wDvmEKk4kwt4pQRMMgwamzjI8TV1KaxxBzd/o4BSPrMI14fBV9+/z1U7kJZLJ
D7jzreBrVu9slc0daGY/HyP/3RwxUz2lzl30jKoU3KuNNusrUfUfAAspKNqghLc/
0ngfLKYZKA0GIpKZOLiRBpHiY8Zc+er2h0RK9nupqEBES9vFVqeJfVABHcLy58Hq
Z/TIamKnYNBfDKbnVIiZ/7uLvpO4nr4WDgLOJgjTO3m3MDBTPZ3SvLr8ObR5Xv5Y
FjOnbUljNw4w3CqrdWMDWUIEfjhJXxOoeOO+qg5aiJ20i8/u0tRwQT54hjPP3Xzg
YuiKi7cgUZa4k/y+15wHCAwKAbIFrm4rJmrbEaddDItcxNntRh3Z1BSQOI1ndO7U
OuiqjaoKGCClANEQpFcu94kNm2TD3lRbS9m/6UL4nHBeIwLQlQ5ec0HIsz4HDWpP
jAgkzzY0a05UaelxCmKihn6rID1RLjfZt+Uef9Tu2okBUK9B+HFGjz2p2ehyOUDb
i8ZH60nNlL7WRS4M5Kohl8m86NDnyOKu0WOwvSi9afPp14tgAekodhEmECLA4vuC
1yvpblLhLRBLRK3h01zcRnCcc+2KZs1Rkcoj3TzNlchK6Ru7ub196D1eLS+VpMnM
mnRwR+/BC50Bp+Cycxboo+cvZ45q1F3zxtS+vPcPbhxMrVxBgHN5ft93bXsuT0yI
L8v1k7iUEcsqSfVW1IYWrabec71Na6l1Wac1UvsD5d0bdIBje2/ZFbecvSybDjDW
9SOhI8D0OGv9sVTpzFXFElh1ZYtfXs4k6Z6s/k6xY94lgUPXAvgqIXKFGpaq6ru7
Xjc53IVxohcLVXzW0SlY9BF/5ACZnOW9e/tYbdXlWy9zfLAiLGLgFeMIKRjs/5DI
yIAineVZEBaeA9xOsUy7+Ne8kGqYKCtUrUm4fI9lazexC5SNxD0DEiF2eS7CQPM4
nmxeXzFKe3tjq1JX9n3yjATwikosKTJWm6aiqbQNrpCAR3maMS447cumrbTqcFF9
4X2ZzeQ6pmcJ2blvxyNgor4wuuYVt3gSmYSkgATVXM/+ieOB0iHdA7/yCSMqp0+3
ILwFbWkyKU3X7vsrQ4VVIsHgluuNsXVU1BzYzFdvXojUEO9dLIJXJj4lC/L1v7KW
FosGlyXJb3MzcwOb/OTsmGorNNS3yWiKifx/fAqqHjQggI7aDQVqbL46m7fYyDIC
Q6jfZmp+/kwwYptV6T7baFR/MvTgnUb7IK0pwz9mVG9rJvzjDkywrp7TgrpdUGGM
0vLDs6qWPylYHqGLFCAkkoI4122Qc1Q9JgxH7tn2FASD17rVCYZCqGMlCRCyswLn
ckToj+krgTQvp6DIiKpl97vZ6QjZIc1gZUtN0B/0Sd2hjVLj6VQBMkJJNEkF9B3Y
kZsAnl3vBwtjAkzIP49+sAxQH9jiHq1CTvuKZO6ppQdIGLZuU/bkACpilgZt7mde
qcrufgQgDxmCWUGUuDIGgZrZNRlhAkEtW+9gCD4hnnvnn0pxhxeh6uStwm5ThOeD
Hs1QD7xD+TFD9crENI2Ux/EGcdVjAFkA9EwFlJTN8nXAoxDRXlgw3smUIZ9A5NED
1b4cD7CT/7kPfsDo9foXof063DBCOyf42TNLcm4e9TxbL+8ubwaFttPpKiiYSkUV
HrVT9+Qk6qSrMMML1mh9aRzuHq+xo0BL7oRGok2A56nTDEU12He7PUEWvXul70mN
4jqv2ImrWR/vq3+FBwYFu6CYqh1qnjOIFrLeOhtkQFSmZUqLllynYoLXohxE/gQt
ZlY3+yNWJJ+cGL8bS0fGNSE124ff5DA9W98EUhUT86dZIverb9Lw7H4Ov8xcjUVr
N8TKGRFevI1is/Qao9jAgz9g4M/63Jm6tGNseJa0VNq4n7yhf+IYc0b/4ybIkEWl
Tg+Igc0SaHqaAuSx5Od726IuYqxPhOfTNLxCV5jpL9ywRR6qej94HR7dXot34WM0
SYXNKyIbuRxfwouctRjXwk8UJ7x5cu6mfszwHAhOpzqp+cG9DWT14ch3nNONRlqs
LfCYB5Ov4xTXVcEhvb7QZrrByQWiPuSrJx1JBf9AyG5C5w1HUU8Ap/IwR8xS/4pG
Q8NBIe09OqC5lxc/ZrLwoxzQyOwdOujlwrGuzdkjGjYW8K5+LT9mawuh6nSR58E6
Xirk2NguqDmeUtMkPtahgN6WHctdBV134qbdiwWvJoalrM9uu7zg4qfVwz2qo+Ud
+541x9KPn9tUWNk2V8j0pHt021Zdc9Nqv4sQhRGaYE2ifJH8jI9eWyVLiy9myLR3
9xXWgzmtZCLnRlZcMMB0BmdzA/cNvGs3+okag68EtFDbt3UntiuOUp3JfwsUd2PD
HNqbF8i97I3hRygj1MkGC7JmtPj/CP4Rs8rh8QIFXBekBtibOHaKw7oisbro9sTr
a3etQmsqyWEp475exJsAZKN2ttwGry2YwYaLD6z9qXDVt5np5NhZ1Gwub9HQ4Spn
6T/wmvEdhJuYhpfUCq3Oz371ROjoo4sPeFKbImJPY9vodaQGbmtz1auMmCcSXrom
ud8Xe3cL/dYbSGphQG4OZ2U8NmCfQzukPh6W1lHt2T5owQbkOS8VltkKdp/9FmGb
5+OBNS4LEC+w/1YE5sMe3hw0x2rXkTBqCM1H04m/RlbcAzfxbp9nnCc/qCv+FrKT
vP4Icae8AQn2reusGKOHv9XNSLLoFGQiyh8nXfMlhxtamCrQuJfymLKOwOkmJOrW
RuyOZQs/SOLoir/401XlGx3Rd+tG2hBtH4ML89BmOgNqK/H14M9yPrlzo3cTwQ3d
cNSD7Cqf5xkr7M0dIQW6B6/yP+WLqW7zHVSyLDz3ZlKqBEfJQCgSrAXhnzt865jo
cTsexM1orIrzXH/EcBXDMNH6wbBTvvdSpDcoNeAvwD8B+b7V6v+kV4+NQ/N5xiJt
27MCiTanaLRZk21AE0yTBE/vrO4ZfptEi0G4ViiDflF2xRpzNlyxPrAvHOPPClQq
O0dKTBS5a/Suny2wYuqjaWWJ8uPpCAfnUSFGIb9nqyHe+vrspQ3j0cfiYAjMPzDW
lU8cqtKGE4eOTxxnJNzC6QkCTcAMe3MrL46t0xfkPUaYfQkyisQ2SGOS+l7TR0y6
VphEwXpx8YXNU2qbsZiENakHBHPrE4rcx4T6P2jVrQYvlX/ua0q3+pC8b1dH8/zd
U4JyZC1K0UHbToJwGvwh3d2v7nlePgNfz0KWuaXTZR02rdJiO0hbL688C41zQmaY
6yDIN+krt+WPuDl/KQSrTN2t2vyP4a52Sbi9UUVZ0MYoD1jPRd7HXAO6utiIyXpJ
vrb8wb8kJw3PsGxWGlbsYcwxN/4JNRvr+w6uvupD7jl3ocpSnRM9TXx9Yz9nIeaC
oK3KlK29VKOIPAONZZ9EeUAOPr+I9d/gfhUXBtxOyeswaSYf0mqO5oYCzVG6HsUP
gipozWvR8HsZEN9yj0h1Oq58da1q0OP3IUoMhk0z95+sNtbQBVK7Olg4H7tC95Mq
7rt88nCWCG2giIKeH6F0L6WIZoo4NPY9Kgl5J+utoSf2aJfykWjxH2TyJ1PSvif0
tHhD4y0MMIujvLZtXH4cSBF/SV4nIQ+cWnbQXlaK7M9XPP1JzQ62+N10CPPa+rnJ
lphsMxNrvexmEaxqYJhhRDMDEvo7tCym/20z+DQ5xF2d+yZHlw5/zz9vknsX0vG7
QA8g12szDQZkozyQdp8YK8hjEJxON+MRgfMt5r9vMSju42IVlaWXtm7+Li9ApPST
1p7TavWIdgjRjD1UFK07AFxKWPpXE1NrjU34syfEMc/iilpXcfwIB2i1JUuJ3CJ9
v5Mv5lntezTRPpxr37dcol6EI4Ipt/o1W423+XLPMZ0GuqvA1eRnIFWoBIZ4coVc
RyNYdyAZtNncmGeDbfcBiJKIIoFnf5h+PUUHsQVBSJjJeUT5ReNIUKoAUDSrGLLg
XLeb6aLcrQBE8x1cFdxGfxlGFpdI9fLC+OaQDMAdNBqzauiygljb6SbjxZv6l1uH
BqaSHUJ64OGePjH1mDr6BP23GjRauaf6iJn4XaX7T353l4q1xhk1j+kpfLNyLYKs
/Lsm3oQIMa0TLQRdBT+n9SBOvF83BTJX+uX4Lf6pL6pQJV9lqZQFe3D80Zkn3kMg
FLxgWdUNU7FTthbc3uZJVB7HmSQOszuhIIzU8/GTl1LQGfmxL2tBPRlO17HQrXFI
bhRSYjg4NvvEscYQbxhnhx2mucZTQR5HsbJLtJzsDETSaokgLCSA2PyTO0BlAv8L
AVbDLU6RwwYREV8nfNUo/hQadCPgQ0eF7mtAa4ZGu0fPzcfIVZfzoiDbV1eSzlMl
o0uQ2La6OZPsoRQl3xuRaFM7fLyYr4nZik2MV8NE+tW69Q4hAB2Gfztu6EDilig2
7Xy9QznVZeu7gj6rx9sSKwtaMruKOKXe3CuD7coR5BtZe3QxmOGHIqD72pPCKt/h
KS6B66oeF0HOFKrtRtHqxBeUcENnK8ZH1r6Zx3qp1x2kNgnA9b7cLbx0zWFzuOor
JuMsB6x3jbPKciC7BGmteabJGkb4FcAOUB8v7vVj/JrP/+f1MtenwtA7iim937MQ
Hfr5D013TJVV620BdFzXe3XKShEAJ3KrGxxxSv3ivKp+gfL1HGrDmaw6jzTSpXPI
unJg3VlZUdhxsqlM5zB0/A7AoGrzBF19kyrEO1SK5ADV+EspGLNotq+pM3xPXvHy
TFri82D28aqwIoNz11jfhHzqZqNJTmbETCv1iQ+0l1V+KYu3nDeKAQgveLQCDPBR
ZxUQNip1HtAnwtPeqbmbUqqUsOaXobPnWZGgPf+MYrrsDLY0riKZbL2YJmuaxvZo
89Gl4KTGbr/hW0HMu8VWM7a4smAxCe0PclylFdv3svy+nNL2Rw6/3hfGDZsW6Eqr
Sx4U6/MAGhsEsdxr9EIQJdWhUOSjspTVJLVW2wONVq256MCWZ1Nn9L4HOsVxXtqP
1yqzud5Z7j3naj0xo7HL1lj8j65W4pBxXtMPPQtgUN1YJe3uDlhRyqElOSU2AMbV
QasZIOpEwiqP6HiSrmAwH8WpoF0vYSe5VQw60tGsPrLH9LAXyVSmukV7lffar8mJ
/hE7t7Xz0S9iMKOHuvkokLIBBw+Y48wucuotp1v87FPcB4JRSrW1uziv3deTNLkV
nUQDK0oDzgx64Gs+HOQnm3Ku1YQhStMmCnA5kitniyj2Cn9sO/GKfcNUXm3XvZ2f
VJAZP5LPWet+G0OgP0bUOhkiqIIjw7pHULwcVHGkchF1fEvQccMFlzojC/3DWo0s
Oy46GS6U7fLhYN/O0XLX/8EgwrmWy1CInzlC/DE01n3O2H+WLz0trJ/wjPfIsdUm
3X50FTbX+WbWS3xoLD9vGBGXBSnecUHYbB/lX+2U4rx3hnM6mZJuJbmhfUsjV3SW
E5TB2h39KZZ6iDQuvlMrPRf3EdQD+TwsfmcWiWrAAvevBYTAwkV501zZuQ/3E5Bk
yJW2wOt23FhHsewaJRIKezwClCN10yl2ZljYjbJNP5Ghu0Uo7co5E2R22K/mWXfw
ua+6FKedyAnGXgWqP9Lu21pNBwSYLXRYl12CB30douMJ8nLMZFqTwnlue7a+xmZu
f1kD7Vmhi9AbIdC47eYk/9y4/YAvpVCLYrE4CNDZLQJ2Um4V5bWgiXGF7dcOVrNH
lMp1AzR7FLqKp7kUilT/TbhJrf1lQbnd6krEZUBFq/MPGq5w6co+BHYZNu5cII6A
E0R2xYA3px/w8suXccpSkY4RjYXTrqGNTUUJywPrDESV775NvMKxzIuGc5YOwte8
RdtdC4X9f8bz/dUsV0DbXu6dPhUoqrva7cnh9WlR858NF3VxTE0TkbpkoiqB6+h7
IJR1Q3OIYEIucqThOCowp0Tev8+5ZOUxapgT4RC9E9Y66gdbhDDyqgjZNCBv0KfZ
7RmVrVuBbC1V5uMXSvwPmE1Hcwz3lhSTYtJjHIvFjVsZLy9sO+xIXfLixVv+tfJ0
5elX3DKBuVVsPwIOvlKWC4qf2I5z9ACSMlsIJeW+IIqy2kZaJ2Gy+sFBlMkPmLb8
KrC/gSi0PiKvk/6MZiqis76tIUEyKDF5qNZddR1qPMvdFAjyc3Cx5o6asya4+WxT
0/EsspIb2ZYMusSn9SLsWfyvEAQ7SBqw2wpbBSWGxjaY5DpZNmlzsQaG4Ry5tc3r
zzXkDr16lRSxOIHoPBO/OHJUloiirpYA9MwqUpTcxfDrRAbA0vHTxVBz2gOcFPzx
h3jeHNreUcyAMOkWmpJvHCtixQa+h5WVChgC3bdK2pLQKM7RgwnryZyG6NmdGSmy
Y0i5rKFC1+1Iubgy7APDxJyL7K3/vE3UvSmxllRn57lUChTSUkZ8ALDzKxy13df1
anmyq1r3Y9SlcsrNzUt2QMsgruvUexS5tTwvUissu6P79b8Fu63wvAPA28qEojf2
4fLw7w8S7VfuggMTbGzME4XZlQTmgNC4akttEgQLFzhRhgV/AK9Tbga2OU7GhbZh
YF3dnrWr4SlnzT0Kdbmcs2Exg8SDcVr75Nzknro1WQCQwPN1kLd3wSmFIurq0v3b
MZZOMasDPhQfFO1hLB7isrOTAAoPhNQTkn1OryHGTOVs68npACakApFBsfWgmqvt
6jvHJo0/+8o6ucfqVtKywzdTU8gNFAPyCFHMmUM2y5CXi/TkksGcu01B09CoLW7Q
YW9q43+rLAbcVnvRQEJYFTtQ/a2DMl8kG+TLj3GqxdjkpDwwkZxPCCZBJnuPSPBf
T9fsoZmwm5HtGGERsxR6lLb8kcHzgNzlCRUk1Sia8UXEgefapFD0YND95oPR+I8D
VcplEo3UhOierR62UvCBQT38ZrQvtS4mFaWazBqm9lgFIjeYz+A+P34DbY64NbKm
kE56XHF1QRn7SPPnaee3b7l9h2HS1Q5yCbxZh4di6++zHkjrVZCbKnT/IN9ep1DF
atcNWgFxzQWtQfg5eVXuOAW1Z49rKuOPBxle32ciOVL/3dImPiIJyZ7NvMgndv4l
DL7FyFfY3hOegbsl3ksSreiP59qQcWvcf5vm6ksKmX11ch2usWoeAYnWV6BsqQl4
ZxjdhQPG4slzchRHHsc14AHVWlCOfkylhDzvof6tknjHQIe+DI5LrrpVrQ4OuI7w
AHaATkjEXAbcW0Rwv0+2SGd5+7R9XCjrU7Ot/O2ea1kPQRBrwFY2PU/tWZQhLBt3
BCjCwEQbVxDfQFEhjdP1hllMPOiyTvUCxF1XJbxEPAPvQImTwtA6pZ6Lv9YhJIWG
mF3iCBbjxJS5y7aWq9Q26EkFpWlCIckOO7R9gn8cfMH+oALAVaIMtzD7RJ2/hPpW
cV6pz/fwV+djHEO+YOlGx3IRR0SLfbJynyE+uDYBpi+FluzGoJ4hqaEr4A2pz18y
+4/P7fjMiAOS0LJGWXDrp6sBP8RqVs3cBbpbzbBIGF8AOspztOjYIs2Gw7H9x3kJ
JMz48AuWLFD7CARI1PjxiAvXdszvL5lHf3ys/w+k/6Uc8K2KYGKWtB66zfM3aFY8
k/s502M8uZuRrYbxLgkOvmekGwL5DootsYigiJFqSO5sIWGVw7QssY5ohGngweHI
zXOR0HvbsNv/Yt9j141gsDYlXESDPnBOYZzenVzMlFbuu/JxyVJAWkN43Vh+PcIB
dahGYbz8m6QXLy9ZNbbnoWu9uMYSeJNPx1oCGlz2CsR6OZ/1Q0E7TKB4t6fH0Xwp
vbDHGoGFbnM9dBVlAqmy8QJptDzfSpyAAoEDgw3CJ356utCPacASelHzl+8LxInB
xTGA5WMUMrZbTxFgWB0eP6Cd2v//FJYaTMqJkrHrG5N00P0FAXswsBAAB7f/0IBK
m0Uu4BGdkjg2RPcMn+yFzdMBWVCkwMx4sWOwqq3UKEJIZssx4TjHuFxEb6DjRnzd
d/ihHlbP22ucpmLtmhFsOfbKYcwe8kQZDWeyoCRVFZyvjm/XbRX6z6CqYZCQ54OV
szUqSvKRIzJsoATxT3TmPj4Ocbtm2ZUnNhqLo3aSfBKvXVO6iMY72cC3APb/BVCw
7ORh6OEWqKCVv+eiC5CfI9UZME50rAkFYOqchMesd3X1EPDqqLJwCwhHlcDvf9t8
EMuVScN6vAUKAsNcfUAEkWH+U6KmzMcJ+KZE11OIkcnnFouC5QE6Q/pHmhWE6s+n
q4cOCaYCjgqj2A2lFd54z/FteP5h5t4Od4Tj8mPpqCGtzwwe77Erb0P0nWDQKabU
2iJ7tnZtp4R9HTg0P+5s33GNfMfClsbxmpj/ODaLNJ9yigAWom9kuBXFIESejhXF
81WTlqBB3cJwbkrtaUGMUyb+N/VV3ouO5OVsFP7Iyciob2gX7Iw32gHt0xogw5tr
WEgPZIRFyAJ3T10P+JvFxlw+ZLfjuzRwCXQx/Fowp8e+Tgx6Sv9B5o1g3DN1SKIg
Nt4Ova8f/jX5SgujdDSq3icTDfgrUpw3jYbhYUwiX/wRnrYFZzGFbk1k2Mc+aGC0
xTDp79zOixb7twMudsZZA0jWRwf081xRrmS7L/atX11nAQ1gR0k2CCL3q8n1rw2t
YAsxUQ88lFuHJgrzoqjzYwLfWoVJh59EVOVv08Hixhp26r0WSEdkWRxQQr3jCkMj
rfy82CJkc/AJGqVFV7OinaAq0VXv5FMpMub+IzBp1nCT8riV8dqOSBTJ+g8YS6O8
PJiHbhHqlRdZ61rC5zCB+sIzBfdDkxXIn2GJlrn284TEjkpdduaNNdQGl55ctAYZ
qu591wLBEtkk5AKc3Hnx10KfzPejgWYdiCOdRMEDE3byyZIEGDqJ0fYjsD6Srnam
l8kCZfqYsfTzKDrUd6tbVOskgkaxpUmul4XZefJzA8YQvdNgm6CNwbdFeFUzy2QP
hDNcpYK24qqem3x9eN6jJ0jwnJz/Cq9u9DDSEOjLY1hyqV2OogGBtpS/uZRbkyVv
Y4UoghR+lovi+/3e62QtRvylwxh7voy7oEFi+fstLk8ReG/7zXbQ5Wv4uaKIje30
Fxy/K+fRJ2fnDIjDWgKgyIZYwXKTujBf3HwU6x5H+1SqIM/f0SUkUyzeTVaZYHJs
0FvsO/WW1z3jymkQFnQix3udi3Gyy0dgsLkYqzZ8uKrz8cI+mp8AWVB8PNLPinYy
xP7Z16l7M6hTc1ZtO4WK3pMQll85NRdmS9v4ztm+k/JRm+qJ29+8DOZ+DTyusDMT
f1OtPxCFxK7nOY6ANNH3fg0JbC9XJrmcPJ+2q9D1rmZ3BOoD1SrVMdRbyNIPvpVx
1Ebg/t84NV4B94Dvp0Dk9cNVRAYwbuiUFTP/krzRr+iCs0bQgejOI88hqAw7S0Fs
DU0nzA/qVEil2vPdu5eVyxPtpFdjV4iTbNEDOZ37X6fy5lDdiLtTaQsVqMMD4r15
PFKXEehqWO6k5IN4Wfp3FDTn43pXCVy9w8erQ6vcuwEW5Zd9b6Qt16pzFfOi9wKH
ivDTghh3wsABj+C8LtC+zlsZTLW/2hyo547pFKeUAk+C23GHZyDpSrZgMru2VH5H
gl9SdGxaga8L9Z5fT5hFhHyF3a78ZQxsh8smQDL1sXHCfUuYyuwceTcb/feb3dEt
YgnWHPXF/9+xK1OEIWmdYMmpCeIYv/57C2wP8p+liQ9c/1f5P93Sj3YjqLmX5KGO
1uj4RoWUlU3X+PVHnL7PamupfCD/wAe/eEPZV/UmztNz3gKpvw/35Ozl8y+/N4ZB
IknklfUONU/66BlyLm4lwt2tfIwXxJpmIy0hsS2jrZgqkYX9JfLu0d0Y6RRyajb8
36z75GyfeIom12uy6XY6jgnUaTfasO8BSKO6Jgl0hJkLzNO4yzFeZmQITjws5Ox/
lJ15tDy+jOe79Y4c4Osh8WMwx6l7Ds0RjcrTiqK8gz649R+eCarnMVQaXxc2qqNJ
kDX8wFfiViez7crN24QkW+L9KacKm3Q9fIfRAaJKIyVhGHvaCZnFa9RJd6GxRDo5
zE6TKKSdRd/uX2kqjAYAiNRrJOXaI9WSpLbjY4s719y/LKqjv33yWv2ffnEsfwqY
F1P3YCxkPWlkxk2PJITl1BLe4hcCh0RZ9bCGGSEMMKX4jfp6wwE0ujJxt7GzifYj
68hRuq3L5HDUhyryJX3mZsxwqNpCGeSMcnzS7DZ3uQGEBYIMUIopLmaOAmLrm5jq
Zy53p/8yNIWJbisNolJSPrKZQir7dUHGrECLS3+cFRBDMw6d+EgjvdO4RzMQddPL
/rYsdvRHkokinI6R1u9x3OWJTo1O2fViQYrUNSaMuJb5/vmxHzNDu6/wYzr9lGOu
6F1msORROcZBYYgxNUypN6r6omjxyREhUbbEidQybYBszrArvj6Z14WeeA3MOoaC
QFLJtaYaoIJZ5xJqw0d4wYS4QZfAK625ebzkI7pb2Zgw006dqSxW/rb+38eBSTi4
jTB90x7pNrRiHVTcn6HWsWqmu0QsNIy8UdnWI8IhE3I0xS2svpWB4PiQazkcUFpG
bUjbk+A9lhpchdcQFZQkRRzZBBbGyT81y4JY5ltTHFXK28t70oIcBjgqIwbmoSlZ
OGif9Dn87DBsdkA5zTnWIT0QXEM19E7oDuOs7mQyKOgzv1QvYkFyzlpKsOa+CL2S
xttAq3QC/lnWPiDUXys8/Adyrp21dP4OASo4SFZRpts6ecp/8J6BglfmlwkNgO48
IApaG4D14B1RvucFDFwLKTok5tPoZbRpuewRa63fYov7ORq0WrW5bm8NZwAiY1/i
SBE2Hpr/Lk+qdp6Ut0sInSuh4NnpDRPtJHqwwYy22JJCl1hZ3ktV0YhW7IHAmtbZ
ZlH3+SwbEwFjVh3RDILlvfuGFO/x2478Jt0WyaHt1tqW4KE7sFP6F1fO2unspnD1
R6pIZEjxMe5jVz67trFwJcf2ax/fD8fHfyuafAyPexQJgwMd43A+4ak6ur2+SMx4
7YGVkEGrasF7Voj0CtDntTIS7b3Wh/KC3KnaGa3EVNNAe48P9/A1GsO3L7aX3yR/
9CezOItacpaXLxw3d0MGTwWsl18D/acmCnSL8MJK71u4Ywgh5UmaTEYHhSJmaHtA
Hxxmhy9veegW1+8t+elywLHhBAaWk9sEY780dG+wBXTdtwhCl+0Kti6qfTp2nWAv
WG11w1xUCF4pm9Uie9VIcdMy2SO4Zp7AZHciARqmIPtV3bZmROyA/x085kI1UEme
Mqr7BUoGlUrJ1co4NkEuKh+Z7BDjM47fO/KRxr4jnSYYH1ICJn+DMjCpNz/uVt41
ybsMX+cWKz+fmkWOd/3Ka9jRcA5ikjLQ6L1qZ6al7Jvam16wa/njBYLY+1ib5E/C
THliUPCRlqe71AA86966p3EtWcUN0uUw7/KWri9BLJyOMtnbdfyV9rl+j0Dj+nGY
S6+GXExqRlUPAbRnDVRe+6wGhYN4OrshjZpqeJ/o2cD1aYzof1G9/O/5Aor9QdR6
3iaqZ5sZ7JJPW8NmbBbQKB2yVh4XCC/yybwRQaSFsO90D9h8dCPlE3x7XKXOMNYi
iDp8WAgOO2LdKao+WKiO+ySEhsRB1KHGztKa9AO/QHdMBhNPUp345Re0vc/OeHQL
Onn6rOT47yy+nkDWNxRKXCM9t5/C1bRTerLk2L3dVIVs+FR3yxV2XkAADeFYz1a9
Hnk4lnWTcd76y19pdN91Z1YuBexiwgrf72RqDopuwOiT2B6sY7VhP8YCboPVcNld
RJA4ARK3iZfI3P54BKDk0BaGZsSpN9UxibJEKf/UMoHfe7GQk9VmQ71BNMe+PGFX
hTD1URdvH1YEUcTlYKjdVXorDB5XufuhmCpuCydh/1u4tq81a/mlW9QnUN34T7uY
6bd6YOalDnwEiD64b1L+olK/gy6ta++k2RetfEq9wpB5SfgYSw/gcii7iOzc8A7K
4JVCEtvgAsT3QSDc5pOXFDAKrVwmf0v+NRhndQfmU3+3ZyJMSoDP5CJY1w09Bilx
eyqx/uRDj+fYxZViQLzLL2XhQDRkGmSa6KoDUv85KGKrOLjY0VrsNrOgJlRRdz4g
eru4+jmBe0bY94H8CnoU3H/eqmGaxUl41JtP6N8fcIvKBOErnZDXlweEKZT/qszt
pULNHkDEDPjbcScCkoRBrhpvaI60AlwubeUv1YrooFJf/J/XjsutgN5IYuKdPpn6
oWv/XBuTIEYI1d4cSnoVix56sid5yeafaSR3ieSR3vsLb8Z5QV+PuoXuTHjqvrks
MUAELf54YNEVJK94wldy81FTpEB59zCnyFF/Mi/FbUxbGFFkGHxQz6s/UEjLPMDr
g7yyffg7mv1QJm2L+j25Kr/bW5sNJ1ndEuTh2nitvSx9u2XPYdgxLfh3SRb6vzht
wCbanC7K8WgnGe5JgbnI3/jgT8n/KWk7QK7SB5WrGrPLAUA+VEIC31XmKgm4AweX
2zeFuGIP/ROPKAH/kF2jYp4j8/CsUQgQyBsRf23KA7w+SiBPTrgvRdh0X3Ah+hly
m5aK+sFToPicrd/1JCMvAt1JbpeL6cSEFvwVgajNU5VXKptoWNt8CP2706z8Vg1N
fdWlYLsuHP2Dw3viAC8Z/I/xWJGva0Ul19ALs6Vns4Y=
`pragma protect end_protected
