// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lyDdoEIijKdGJQ5Mjr3iH0T6dN1nubbhPTU1+Vw3R347lIJme9uy/RrdUKtpHUba
RI8Kt8sQxdpA/R0S05IDQBygedGihmaFSoADL85mhVXPQZ1fFLUKYTHnFCHE9Ifh
qPlBdqOIp5NFdnc8Px//yYu+8gWdCfGk/UFnEGLybDc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
P5x1Iq4Fq3QZKf/VKwReY28/6N1Drcqa5fWNl1mxO+VXYqrA0jLLXRVQ2uyEd+9M
QrvLwS4yGKjfia0hmeP5DbSW6h12AiXOfrMY3i0QobJFevBf8bG/KPcYtimE8gCy
/eePhukeqq5z12G6cKBPqDEChmShTIKDNprIGbzJHLmx9FTC8rEm3pzoH3yIRurs
ViqYFLzPJiuOHzJrJs7uK5D2Fx6vLk8UPXECtXwUHt46q7r0hRq8gRAeMk+S1k5D
EvXMdYDAAou3oTOk6C8HfDwdK8pR3PBjJl2y6D/I1SL+mcaCEPsXE9smAF62UHA6
dtGcITflhchxvRIIjXhypCVChoB2IrBQ0BiNbBzc5Jr/1WUVUdpZNJnnXIdXKi02
hUXqqDpciaPaL4gFnUBcUxyD4ufdmpYPtqIP4sRuHHbXcCqRlJHXiWdXMAto8Tfz
SMWei1JNoAkVE7tGKPM6voUGQG/4VhiFtRNTireveKJ3nmxrKEbRQVKzeBXc7wIC
Ozh8Jq5GJq4wppaxkkj9eMsRIfVBUMEHztKn3qKq88UCS5SC1BXQSy6V5erV1z1N
raVaMDsflTuwntfzhozY2/KR9GKOFAf9x5zGwoDA0q8q6/f3yCzQBZM8JIXRNY+b
a4ZBXrYr81Q/KtQDfBvJKx6R/njZaZKB88M6n3J7ZwualpA4FQwQdaG8zkdYM4SA
bTjEyernC6rwj90nwcujuJLUgSx0PbUzP/jOSYURUW9Mhiujr//D+GFgOI2iPvl6
WQ9+c3ff8bq0rt04g+hnnus0aszJKoeYWzimBmWUImBVJLdFp0NRsyF5Xe8TcVAb
ee2z24viwnNP0JfEtCbWBLQaNEbrchTEF4Rb0Q3adejk/tkPT2hkxsULIFh8AVeF
yKpypS2ZC2gYSNa7r7MDwfI5ngOAGvJ7pDkpZNBMCFlCI393guXUZ3MN9xc5qR/d
8CYpCqffzXmL0b7Ojr/iIW4DMSypyLAnTuCn9uj/iYnJ5lXRR6R1X67yIQaKcGL9
5j20uZrTXKwcmPl8eNu2R9CoFExw8/KJ2f0yHve3h3ZiLH7kygXdEmEb1HlKBQth
0ufWfctkPHgjA0vSmHHuopUjOXxm9pVFyx4pdxy2AeG1Qnu8PGBS+Bl3qPR+4dSi
EA26ukbx+dLBV+gdd3OHnhQ8cEkHGLhNys9VYZDK9rqq0d+q/btfq7fHnT82xzxX
VBzjwMWvGFrZSlSQRslJSHjmvVkPAwSZXsIK+ibqk3njv5dNthdAr1TCnTlJwjWb
IQ89tKbtoxQjTi3rKyhZ+fXiCWvd+D6wHhBSJkejudZl62qfK1OpaPWsgGHgaYp+
LQLdQP1Kh8IinYpp64eaLu6Mx/jpAI4FYcHQqev3Pjm2lCpYu/MA/Njl2Io/aGuR
ssDlqy4pyl1/CqWYp/8qv6gmQAaaXuFFzjsWc9NZk+z7L7j/hqpSExEXMPMqTSaI
4ZsSXxO7aR+ucOczsH1bM3siQEkktRVyRLaiwR9Xfh20Y/2IP7QJKdYWvC/VH5mY
L7F08ScDJZAzwyfiXrf7SksLltrujW3z+TWrzQL/WHXZsly6KaH915n4Nv4VWgWm
JQC0uJvTfh0QIKLkLk97HVYdyPHTENQbuhC/XbFHDP1Hf+q4Mkxua5wIcfgePeL5
onnymeATKIW5XxLtmxUDA/y8xYEH0SZDpwZiLICE0PbODblSpWsbYWhR4sIPRbTj
D0aHY3BoMVURGOPXmuUFcQo2vFPWGNdKOc78DeJA/C3S/erbsfCM7GHVDQjSBQWE
+98esPF2z9+MLRzZk+kXz8dhTcUJWtABJO363lQlToRoFTsw6LPwa86im/zHTHkI
+mxlr5dmDOE0Cs2/Oy01ji0W6AVQFV9vMjrUJspya6kQ2Xmi1gzCGwBw0iE/9Xx0
2iagCNQv1+zlBH1AKc8awsatx9ZCBRozqZYEzfa7aC7LIWLkjUMIDFIEUZh0TUG2
vMtSsxtl7Zn9wluLDugxnQyn3AEjrFQ+xwIu+1CCeBTqSQpVnZSfxdNqD5gm75Tk
JsLOpvovYm/T0m/AEIp1ACxS2HcyN9pCTB7IUWCVwbK5htKvBScyGp0vkiJFd3ul
ZJ0ylypF6dXY44/gcHXrxnyyyd3GXvhwL8rstGG66WK/a0p5c8Y0WKDUHAOHmgAc
MDK4f0dBRXJ7NKVFJKTDDr4DpZ15gArjee5Dl4RaYpMMFhU1MEfO7a6tDPXamxFx
ruC3G4KxfIwVKXbUJP40RA0gR/ZmMODsudYPTe94E92gpQw0sScQuKMxa/OtCX9A
4V/zYwmaApmAr7SUaeIQb/geEniBicVRQ00qy6ttAsz3pA/AzQmVTTZUcozPDLL7
GJdAAaVfBB7ptflTu0IxAXLCvTDi7neyFfXKJ+Wz7Ut6Da2ZlBRC/iZmKlmakr/P
VbzT3ANvYweSCsDAgrO/r/yRFP0qRZCJgXvAaEh+FDpJUY0rOnaIo7Zn3MielYCa
FrqvcU4Eb3NhBXML8kAPlWGiCIWphC2RQWB2bLW0hJ8rCdbAjFccdQcFayB2Zdnp
p2KSDBaDoh/AeprsaHY+JugOdbfSrPLRB7KyYHkHgs2ArLAMjMB2bRXcWrblXY2z
Qgohw1Yfu/ZwaklpDLN2F/ZJvjuHUhUukm2dvWpZ9A8qqx80PlbgwGq5h8YqoOdd
oS7sCEuYwonqG6M3+QpkIzD0/Fubmx7IJkbNEOd0p+OCoj2svzLRLAwqJKFaFoB+
4JzhzW12HPgDQfL0BHOLWbqIkrRAOlWEa6CD75rSQIiO2l6tndr4IFLRkP/lqT93
4RGK0oHXQBQyOo3gtpHXA45bgME9qqlQDM1iMvQlyeLxFOq85r3X/qiKE3EFW6xw
w0tDBKvxnQ4Y9DfOE4bnKimCdrbtScCfdUSviINnXKISLDlbnBSZ9r8dxpgOCUet
udjME2J4cWqjr6F1u654Dx0A3zgVXP9G1Cu1hHon5C2qlZ9y1odKAzwNqcmTSFaZ
Uos8R4CdRBIqZq043hYApF3D4cbhOkpIRjotW5y9LBubLx7mfQyFU0ZB+lUofUIr
l/SOCIZAhiiWMspIacLI1StWBqeROX/nWxoW8+shScKUdCQwdTkvYxWSKXDSJ473
Aw9zzP756WtcFXkSJ0z87G4n3p/DQ5uEAwFQ5TIN0prHRP/dHvjsWNRvQ06+IccU
8A1SeRBaAisBsyKh4rMJe84kzgqeRgHu15rvaulpgdRbzIK0nyuZuoDFXoBY1Ols
wgqwig+a3oNSLnLUABRLZqIG6Il4wXgHpS6LeaP8i9FXpAKPCARg/+ToT3MzqM8a
7gjphiN/8/2GiCVx1c0nOc4nAP7e9IK7ubKhPSvuKDA102kVmGf4HCQjxIJG45gC
jK93shgPL6wBAVp4/fYhK7H8w8pxBvHKl+2T+0xRlrxUHEE80kfF8Rh8XVTUqhBy
fHUDj+z9SaiEm1oVceapGi0WoGSWwzNyHjbwCxFmIhXauxy90zbK18CWNXfSVkCi
D0AQfUP+9jNVjPkZexbDMzc0DbqQWtiyoIsM5ij1/Sd9+AiWjWy82p/PXG12iumA
s+64JB0zCmvLigND3foMQ/bVZZYXFD19F2KwfNF5WPToMAw8xYsUCV3GTcD3/FzE
WuXtzbOCj4BvvbXtWr9ayyvLcs/zxs62jOwdZ4qXOv8pVx2m4kmc0QYk33f53rpP
QHI1MQVySU1d7ZXNyn0s1b+OqraHyGhUKVrQmuUZrUe1YGI4BK2GKiVvfGFDuAeD
TD9MfIuhTzDRq/MIrDEwvMD2TmOWyTOvA6Ng1GLy/Jr5idJnRaRDOG8EbLJo1HiP
Ylr6HfMmonrUnYIh+RV/3cxUBtUtndlTNHkfQXmdFtSe+6qEgw5YM7+/tCwWsvNi
p/ihIWjBVX3olfgYQLkXtpO7Hosu2NG8W/22ShtYzKYaiCN9RWRbgujvEezJuuB+
hauq3KrCa7q1fKJsNXjTIg==
`pragma protect end_protected
