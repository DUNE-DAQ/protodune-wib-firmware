// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eEi0ocPXrmdCoFMc3myPOpJ5xNN8wx5glRas5jh0wnxjzmy1GDfGeIaW969DXHQQ
f8IJyMW5l63HnYJoksjlVJcgYdoV2rLUgdpLssktFETTtksZYp4415jM4f5yFxN2
Jxol5xeb+kub5KUSRJGZ3g0mCz0+fOWUE36R5DpPLBw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27696)
Bb821ErOcZBE7Bc1I9pAh67i5QNSC9RkiaXn+HGSOoXkzyjy8MzWiQp2yb+uyC6i
1/p+Wcq+rMXQTX3yBFlKSO20GEQ9+EU8db3dowPtvDnc57x15XN2cSeNuvywTYpm
zcL8s01/eM6Ibap+eCBSbgItAQONMr91CoskIGUUL5GxtnBzMTcnWzF1jywy60/k
1TVLTta96Ku3m9ODyu/6R8W1sg64cUihiYCAZoWayACNtqkjeSQZAjlmiVTQ3rIT
6XqCQHJVUAlVEFYCj4KlAyeTr6+C5+SYw3XtwbjUiX4wQwNAxsSO0A1i7M1QSNBG
LYZ2qlZDtIr2MP2UliFBmoWgBgnLPeIru9vbgnHxZxl1jlZfnWHeIkoovR9vcR+y
B3hjwkBwIp63kT7uY2o6U+Mn3zpQU3uoM3Ko5r91ZlO2T5VIIE/9x2a/yd78s45R
S8Ae7GKoldZwcITtj8HY+wpmHIJ9mnOXE0AHvjn62s2HszU+zCgd+Mii78DZD8hZ
s4r1o2vwrKYNHMGKbrX71gCkC+aJMoWVv0mGT+H8Wwk80tySyhEnnvtBztqIK6LQ
ibP6FNy52ENcKtdabNbIlbePdCgQkh1zwEtgQ1/466jTbeT2TkMpPVrb9xB7Mg7b
BtCoPbUHK7LKFVTjV1DMQWo5SFJnXNOzvejIO5KeEQng4SB4Zf+NaWTf/bb+LmFf
2oNREOkkxyLe4vIgCx2HYTTY2ZRmLS1wuIBhnwns7hp5uTQJZBiSUbNMPNwi9fFQ
Q/sq0iGKUh/EnX6XHQucc1r70sH/wKIEV+P/Oe+ePB8tGafbqlNOMqYnpjbolEhK
reVSlS3B9ceHuSviJPGz53dupL8W4TfcNxy/WqT3BG/qNtbUZgdELN/rgHgVM3k/
UlIws9+5onXxvPacsj2jDLOlFmEugbPcyF5DemrfF4V50YLP8aRIC028EEZFBcQa
wrR5rl5JafhhLjgiWEly4jVYnqX85uq6EK+8JGCek/iuKwSKVYOcIZRHTqtGWTNI
MbMBWCY43/K2xWuw1Vroho9bp+X0Ys4LxavIwDRViOPkyySS0EqrN0jPk9mwVDVX
T7Dz4aqT0oX4QOYUGm3WpuzVmg9z8JBtpFBDT0VkFVDtzpjU+eZIehW7rWW9yZk1
75IP9QkYPqSPT/UAee0CNmPmrXNG+1rrepeLth3BHhgOUSJQcNjQrIsWtSSjVeDG
h3qgZIoTH/NeLEleqR7AvU8wlrukRAZDajlrYarimthyJ0V9v5Jvp3JTKnjMumt4
OgHCuU4Bc26pe7ZF0XjnSher2XN/t5bgIY+c0BAay6+ie5dF4GJ2TgtnAukNg+v8
3MSXJGakXS48ovRxGl4eCPwIfPy3fR170ZZi/ERKaP3Fpejr3XF+HtSrRxhq07Gt
/hV8FKHPAKz+asGevNofya7Q3I3402+weNglW9pMX8hbr9/YrroM152D5xTycIAh
0UE38tJ1ChfW0iWl5iJv+YA92aIpe02JemSQKnn17NXYzmk2DI9nE/ca3cpw4gOc
gCXn3qE59+WIxH1OSz473Fx2/x0UtryegsbuTlubzHaRWQT0QwzYk5OkaFE+frZ7
Pp98qhPfRtsTQ1X50cnAZ3mFybG8g91/1sM+HgSmtWbqh28075+F2l5d6eILaoiO
5Emh3NLTMdj/LKR6czIvuqfZc7ZwL2d90dMRg5BkGzTr3EIYLkMA8t5Qbw1NwK5I
dLAQBgltxRHUX/91xVSF1rSJRvMZgDrfybI46OkuUDFS8PDdwKmvnuvYYlpnl832
hJhj4ptqmPaC5pUIjUtaOOLJGDTMaEg1T1TRXcxmi8btJ3Tq2gZoo04gyUZrWcsR
urXcC0I5aL2yeQMrLfV2uzC9YDyR8ZBCKZQAN38nDQGdkpvclxDobds9g9R+p31R
Cvkd8L7JwS8+srkls1kZfIXFY2VXJWGRU3ZsSi6nTtg7H/i7238wzH4UgBGOho77
uRQwsA8rC2ojugsYYRk8umWoFp8LlnKKfROC4k0rp7OxpBOkwUbHo+TVef1ZgILL
cbcZQcUafDEnXPrCAkaBS/9xln0ETL73MEWcH2eB1NXro/X2ERP/nyLI4QYHWqUu
Y4S/gzMy3NF+RG76dToWyDPUVPiBFpoxwCdhBkhQ+3i4vZqK0Y0seY1ja3wneRgw
R5VAIViWXVeVmUHsOnUp1gtnaWPaLgYFJjzQTWt3O7t7wdBgn3p8v9rccBP2VGvz
dO1eplmr6Xo9Z1trHAdX0talC/2aLqh2RUG2nyK+lEP1OzSJsC+hq1NMrFCEMfyl
3qIEdV6zgjc/HJ25eQFD3Ql/nqj4mJZaKWRhmHdAvBF8wUFLYMvTKS67RGs6RvFZ
4ITRJ/1iT1FB/ZJQ+wvnYy2sqH0bYESm3kM/Yc+aP93c4iJ3a/fjvqXx5zofxmxy
beCo67i4/oRK+QfsJUv6oD0fLys9zjXpg4pASkZchemqwLebLDbIIQ5qUPjCw/YW
wJB6NdqQltoPzBkNRb7lrySq4VPsULiDNDHLco3losjg7nWJa0h596w8sulGdvN9
kcrQ9Zren+KSqHWsSm+afuwAwXN6uPc9qMDNDg9mTYW/46vl8dlhENCykCGg5Bk/
N0QU2TB6WatBe4cmF3JpOMpuIqwMeZfnlDQYzkhaQMCH0xMdSGRLRMb+du3qzV04
iMTj23D2RUxORkSp1CCHhBeg1NGy7yP6fpjKYRSSDjXV6Tk5HDrz0ZjrvoTnScvK
Ti/gKl/OX7SoeZIlbFKaIYxyCRWLmH8W9dP6aGhPh6K8+5gsMPW1ykDzXkGgqDeW
T2EC4LI1UeYXz/+oOlaMmGH7R0OJP8UU2w8MFz/fRTSlsd2E9FLM5EC1J5L4clqI
36HdHtn0Nh/53UVVH5pblT86RWrhxI+gHZ1KxzfH5iZhXVz2jGWyFx8G220/Zsjq
9dyu69Dy3xGty12us5Fvi/15cU9ugqqdEN7mgTpg4+tot9hLqyX5J6c2hhYBVGaF
TWYq6GT86enIBNrZnVheQ1nL2gJWv7TD8VTw9RN1aGCqomk9y5btNB5ewlnYfguo
upmbwFq52B7Dw6+R3opR9KsSN3PrMv/alJeqrk7+TzFBcaPAmYeA+OKDHpTLfqwo
luAR9NJJ4tsO+D7fcHjgfPNF1a7bbpw6KWxH37Sc3wnqv/E4CKSFIIz37Rbm80IQ
KwVkKBPtwpT3h5VOWxhDCyLnAuvi5b3kvrWUYj2F6/K/8wMdoJwOOyXt3V9Oy3GR
vsSGDaAke9dhj4luOIFCOxdolXgqZVkl1hpCwJKW+dOiKWjigGsyhU3T0ry0+CVP
BGXtDWZ38G1sYCr1rEUeyj3mIQfjfmfe430BLfMAcTQuKRS4iiqsqqhcGm1OjrP4
CK3+oKoikKo2esqsw6e14SvgeTPUa79qG6C+kqoTbytZ36RwrFIXWRVOj0GvGeM4
mMtaXJQP8dp4mMnXehhcJ4vf/wudbSObQbtKg3GmaamyGcXVOwHgUMVHKPn1STVK
d7I8RoetNdf0tEVn5C/WJAgBOZtQliAX5ZPWm2yHq3erb6gD/t+DXrDfLbD32vWM
kvUaIUbsc9Ej6ZXzsLTTQCK6XQSvOgLKbqGpQ6vTdy4HXBHsh8pqs8/mz65QBzZJ
vZz0nPl6ClFso50n6gfi9XIKHuSu3+gaAh9bu/i1ZH9G/hz+ThsUfyF3XqVa2Pzw
0eSL2lisbmmKyIwuVjSjmwoXaxxQrvuIRgH079rM2frXz/2P1NAJAnTyjsSt8eh8
JNPiXasg6BI8ceZI8hzdr7A9fOWDsnWJ5bI54YskjstiP0mTpYSp5E3kTdog84mR
7QKXyHdzcHeF0bCfd3rzoxK1r6iPX7JPtCqbrfPUPN0LBJfQHQWvBqgdc2KiTG95
pIL5kuzxm16ITOiGSa4FjNmg7TaGDayMgszcjoCpXyOafoWLb7bzMJcf+GVW5xOu
L0GN9FTsq54qArdPCpus2YzNq7Eg5Cc7SNoXtscNV+u+01be/IRHv5bTV8t5GsGf
uGmnnO8bZP7Y80NNmJBcoe6L60D24FJ2tPLu7RE7TjklNYBPtrb9VM7BB4/4NoBe
zEKHEkqjkofxOnSiQReDpFC851tTdRS/KcVDia1H39082a4IEqyOZMjEom7eucJ7
iQRuaNoPZJYPBTaxgoq7i9PzWSUUa+QSZV5MElgLiKXz5a0KdTrJb4KSuNjOdhw1
ckl60fq3p/5O6UL8GXkS3Jb2OxvGvNdjI/ZSuBtPMklJ+R0EBUloHCYTjzooJ6V5
+Mhz2yb8tUDt8cQvkwfkeaK1wMGyJNVd6yvIipE6AvNIO2P8fkqdrcA8OFZYpoGq
a3pNZsFOROpF83Vee9flpr1eJGC/nDPbxAyTHLIKV65ZFQrKXChkH9aHm+dWIGol
HNYbIRQRU57DD9HBvzDABpZmmShZwalAEXWcWRPJkkg5VyqcRnb8tSFsWp1kgA8q
RGiwZeOikJga/NoheSJMDNYdpk4WcnWAd7PFP7eY2AdC2ml1m9EuN9mphDLC5FC1
IwfkFff8tM9fjkihNL6D2Nt2P0OuP+DAzjqG0rQ3WTNGuHmlGHbsWmOkR04L9vFJ
UEgMuj7+kgORMPxFWJIUeNQ+G5HGL2UZEIdnjOdSihLCj6AonjOPsvBo1NL3ODrc
Bqtgy/KzZmJfYdReQ9lmfCISzOIu3YIY4zA2qB1vAWf3iAT+Yg7FKic5iZqp4ZQF
LTHMBZbt2Z7VwN6lEUMVLrCeHYruFx+gGC/B2RoSK/Z/Jw1IcERVUUs6UjQTt/X+
L6acXcm019Q6YiKxAZqwZar69BAf67xXLxKjKxl5pxfjSd66SJHb9eaQV6Ox8aMB
UOrxmtJwyr+f00dOnDvP/QcFN7VkL9CL0VPJ2T5cQSEoE6Y/NO9i3/cBtF6fE3U5
YsHIhmNM+K4dTJDlNo2xSPP1WCeZZocU2gS66cmAlW6Q9xIE0486aiP3F93SfhAp
3LZ+Enue1p9FRpmV9EJzZZFRRsjf4Sg94vnWQq9yFQfhK4cWfHoepEpMAXghQu8r
kDeY4ujAp3z4hsT+tti5EZtX9z/OnMvE9lWv9HPIHr9a6ZfiZ5vaP8ZPSQbm3kgJ
hTrgpKYvTgCjv/Y5TST1jlphP5tjPvkFCkVaodNPsNML8oOFwpR/yzS1UUaqf0mN
wK+FOBUTTX8Vd9YowFDZD/DMcddq514N74oe09BKYKY8/WmkUREcRP2e88PkdLUq
nuFBpmBkHQNdjBUnixYBpJR75X1P6DJqzB7mfzq4C+sTOtYJLaEUe8bfBYMJnSU4
6DFZEgQ5vIegLgXb/nC4PchgRL2DOKehV05J7lKnMnh4XZ4RRToSAUInd7zgjCKI
4JjgsprKYtLUESihgePLJVdaCl2uf2TWeTUpT4/Br1XuTEZfVY6pcIQV/2zriH2n
+6LwHx43+mLniKgVHp1ISPoBHB1PfWy4JA3tT4/n9SFVe3W0DBX4+m+bAxVMx5Gn
lLD+OhTwm6tRF7Emk5jd4GyNuliHUv7qbl/LzXkbHnxq1Ju8d+iNZ6+CSSVoCTyb
dixDlwyfUjM3Vc3oK9spYA0k9iHbTmCAeqqI3gbUvHzwcpEsDpF9H68y5g8wRhkD
WEVFymDOB6kNtBMjE8JE5mEmZ1RQeJ86fUeLUEHlReTJrHmGPL1WwrwgBndjey2R
grZ0+744IhVo285kCpTRetGgxDePhP+QECUFKdhbd43IVyx6sMMhZLH1t7OLP9/y
yQBjT+lrfgm5iF8SNxqCF28nbyn/jIXYNZiwC3YR6tkg8hxJYSKIAR4fCxz+PJJE
1rvQE93vrxZP6ag6Rj1QsIm8Rkw8VDmXwI/otNt3NEiKqweVFEl6CFydFbsAm0XF
Y+596x7NrDRslI4PbKas+ZZN3MsM4wnRFr1pkaCEawlOCHCiJdluab87APkzENiJ
AyGqSloFuhFMgnbuzYvRIl+AEmI06On0hO6Gz2dTBLAFTeGVvBdGSIz/rPhI55F1
NQGfBZqhjOLn2TD3+BB5FC5xNc7wX/Khv7pwpNAZCsNaUw31pBJe9juXk77SvgAv
zR8UDxRH6efKZR/c3BtLBk6KiLPCuygpgmMOoMynrGmfPJj/40BHt41xH8dMi2SR
qTk/GBkHUQ8ms+YgCx22OYjm1dT/7tT4AmurbyIrwMtJq/jafnr3wRzDOI6fyBmm
DhjV878WB+iZQQgBzSZ9gdrOsdMJA8fF586b1gHYIU6NfbI1KJuroIR4bfbmmmNH
YBsozrMkDFE3FrCT49eVWXgZ9ABVDcGMDtlZWE7D0cMNjK2xx2jd16bYbWgYdLkZ
PHi3rTwcZg/Pm9rq7beVxiFXMB3VukCo9eMHsAfV1aNKjwvulxUgN6xczM/xQP75
wIM0MYxgKLnoPmepi978/mHPqn2n3skqQiiRkJQ9Uf734Y8v27WSio9NsWkB8fVP
8lcdJZUh3C3bOepWzfbTRl/eQjHa8DQPmalPLLcWl0J2NmRlXQLOZj3laPl2pKrT
quo6j/oTm24Uq7fZpUfBNgxeG7NkXaxMLo/0mbG0YW2CZnbDMdk60oEpkjsKMVpe
wcFk7NCvC6S4YPtz6fzHkyl8tR/dd0Sz+K/h2pRnn5M2HcBWxocXYltC0REa1vKF
3nMj0SPEDX38LW4Tk1GjSG37o/Im3oWsbmrBZgkex2XHANEXKHctVfeo60Q9X7rg
q+UZOlf4JjXyFOR21dm1yEBbt+/QNgVmS3VamFfLjT8hH4EkQZJaqlQR/VBGVEtP
KstFs8b2tfjz5BPOv5zaNpYuwgIOv+4aQVBvysU3KlaYGH3CV6wT8Wsj3qwnB1wb
4mIyKpwbUQXlXRKGiKViZlFB744t9F+Wh1kqIi64S8HmWuBH6WEr3UiV6mKDFtPa
5YDv9u421/67Z/k8Bj7S0eZgrvuaKNt3M36EHg86l9Yol8WH1076yw7oCzYUjJ/F
FmE0LAAaj/tz3m6IuErWnQSiJ9HHQvpFUIcQCtETRnUD+0N1YuSH/KGPO4OksLOd
lS1gQ33tYMGu/h3vkDiouUhU79mBn8RzXxfwaxwiQMmdUSFLrvebx6/SkYje8IVz
0jnNBulTTBR5Ym61CDcErI5KUzxDNID7b7jDVI11xCd32JAScLIgQ7ocOCkzr28l
WiPZSyORAEPm+PzxbGNZm+SR9vqmkaU+s8kBt0kMduXANAyFUWvFqSfvaLK72D5F
jgzIRuTOnyRzGrur6nhSaQDm1NKfJqW4QWp1qWsTvn7rJk8j3MLLImfv4HK06kOE
1FtRoTU6lvlBQYK1At2Nc3bE05HxiHfkntOFT5P6MOPJHYNDL0wo6CmvilXc4+yN
cAJtHk9AjCJzPBliNRezShfS6vE66RqYl+nwW7WwMiXVcFQ0C4q9qyjaClsFsu7W
CXK3nrDHeXXP13tjpGU5DFoyO8voWgACbKp/22jpZ86dx7CXeMgJBz0ofN3w7OWf
otB5bDbPKHKiTcZ1cRI4IPidGv2EjMHoDDFrq0bJx1cpVCxwcOq0nPUQhVpclmCA
taa4q5GfwIshV+lnsZ/GghpJwxM+dJ3DNtOcrkg4yi6JqHggcS9T+91mPxHhT696
ocqb+iC/Yynr1/8a6SDCOw68IIoOwqjDDtmMRDdZt30SjpWBdjTEDaRreQZf8lf/
Z5FN9+iZmq1w1or0RFUQTn5n92Bv2/ZtHuS+3Ne8NA+6mROnzDAneKmay9cFXmkG
FvYAexWVvO+uumYpP+h5/okXDFTjLLh3bPGeEQmO+MqdP/i9JRGk/ptiGsw4wO2Y
GpOgoMnGCJo9ROdrRd0TQ3LplSyV2dXmyPLu9xOyrF+DCd7ZBcw/5Ijsw0zCGBdA
ZW0s4gxBU2Li5xSBZEn5cRnerGFvf65ILGdKawRuIj9TurBkit2qt1kmoq3TfbTl
LzA0MT74vKmsZm845R/s4FbT3L3ZMxrW6ggcX/9JxsJYqKm6hx5/D5wEBUWjjvAV
EPobVVuETyCkUkoXrwbTE4+5wiosBQUMUzV4XiGoej1yO+kHTgOuTz1++Zl2JG72
E3pV9zPpoiLuW4KYu70EpuOhvD3PT6GR5WuypzZhWm62cqgHlDfkbxILF1EkBzyX
NKLjXwriT8mUZdiodVkn3cejjG4sYDNw5pcDjIqimCU11w+4u9c83fJ00VjbwveM
DOKfji/c8FsrIjs/Tj1Kly1lWUpkn6Sxmrtl8xSmf7Syo2upAg5f09+76sfbzjk2
2YEzTg1lzywwfqyZx5BkJoKojeTAFtSVlBFsk7sfrwifco2q+MWO5/4ZzGOvkS90
xdxCJCgRnxq5STgMY9ztvkfnNdY00knxkUe8XTb048IuFfl/4ZeEiZsBOWVKYJuN
b0gpxEteRV/ut6LCjc006tQ4ztURR93xz3/+j/SZLeZZOOraE2eehDNSXMg1VDCS
EUwoth9bqK4D++n8jOX+8HhXV20cHXAHjlYEylPiDyW2I0g6lieXFHgyuWIDiD9f
zVVjmWSnZNN6obuOLV1OAlVTRQObiGIJlLmwL5dHgwj5ce++bBcDAcEmffDZzVje
JXmHiDcWJ2s91TfQpm6cnSxCwLuzqf5SSPLPQZwYnbFE9YAf2/IYW4lWaprcItOp
DKT43/m9royQvNGXFkOtQGxUGyfhR29tKjzRJOxkkv6uApLxWQvzGLzRDqFJwypm
5Ut8/VJVcRQZi7ceLMLCbqi8gV2/q2W1VECuD1tW/cpiWGQ5W3ZYLig4dS3by/hL
ACgqGvJwlIW2htuAjEgFQgL13dsdywNeUElIqCePNcCrh3v/Crwq5iSpSngGdEi5
hJZw+h4j83jXy5zx/J4pDIpZopUwbSIOwGyAKyO0O1fVfS8FIOHaHGTOGEihq9l4
sEOKiMjCkOaq9VCm941z/NqpnFm6LmR9dSCZMCnNVAgK7Woxo3d4cNOp1fhF2uxo
4g3aQFZ/XQmkkhwiQQYlXAVc8E3IHg2e29X/4Oyk34XdtlygZ29+o4tBoswPlzrM
wqpiQM3CY+7malYhwyURIcIm0yCkCu/NarMXynjHWV6KL46Q3hHBgReYxc12INNY
xS+/AWYHMdXI3+PmB8Hsd/AlSz2Sqedkciypfz252ZWPmlJEjRMv4Yfzhn6miOwj
C1OCdBfxLZWZ7+JViMihoYYtQmJD/uoUuxf0SxZc8TBSc3BToRwkGOxNYaMRA/Pz
tFTz7fnKO5lNRTKcebk9Vt992TbdXo10zJ9KH/pEwkCRjqMyA5w3BlpDfcJbVMGf
vSBZ+xOzW4ihbExv6BfeEeZ0PrcF+0pY7KiJtPz4Lvjz5sJjjgrbAsb4jCAZzEqU
7JK+hp2g6fg5VLRzQmda+DijvXHMZ/B9IH2bi5t7M9u91k5jkwbuDgi/bLL0BWwV
+r9FFZijhLpxPOZLV+dFZsVqKv3cuEVexj+PmiGOmgYcFyWGr+Z97V7UO8bLsFjv
yFFcn4wpV+0N9JMc0fbnodRhR9dO1P0W/BKsOf8mv8OzdY6MHw9+UGzyitK/tZhX
ZbB3r289WB+crFIoVla4uJNKO/OpxKcYyjHI5nrvO2dqzAI2Zcl3F4HPfcEVz8VV
YCWNVL/6JJ1/9pu6xmQXkMQQOudnS18QlwF5n5R8EuLat0C5LMizypscMD8LN7SH
rKWGSSOdrKet6mzChGMD7NakAYh/gP6wkNkcoyKQP7qYpXmoBSTark2jmcAeVG13
nKDH38f4Ia7a3Y0V6sggJKTKIjX2n8e5/cHPClVWbDjXsrzD92YeafhoP+hQscEE
et+lBUo7T+hwOI13gq5cMx0ZpTb/HysB1jNoZfK/pJ9KV66pjgqtoD6miidtM+3r
sgr2uuvzqojQrOuvYr7hDAhTdmT8JPE6U/5k+lX1a/X2+mxQGr2d5YRp3rNmxTpt
jeUFaQO6pOZkyvKgr346pZluYGYBfZPu3Xs7fblFHROgMiRsMvqgeC6hUMx2JjwJ
shi1UpOCKRBl8MEJ57A4dgiG9JSnZwRyxH2/kKCXy5kwX7xEee1mI/2XkUPH7/Do
eTvcN/85peyO4JNNfFv4I0Z8K5H2/nrtuGD2dWueKN3iAp+rKyLmfi/b8IrVXMv7
+EaMb8FjSt9nEH9UJAMm/R3VgKkNK+V9GUidLAGPI5GT2gpGf9ovBxT7gbXAUgaQ
xjTvSVfbTkH1Bkd9fTtRxUt7NVyKijJZs8ok4kyCCXNz8RCyQnCf4cTn10U/EDoc
O5H15TcQre6XBiNkAjSr9aU2DWRp4TkWWbxi+bbqGbxWK/CWR9pMgoFiJeRQKfk9
4R0lnKpj617eAn6WMPOAR/BuPOS0VxIziA0IlNOqCmq0GHyVSktP+mXXPVj7XAY+
vRzbpoasa+5npMK+o4ymu2Zv7T4+qdWQDAbwGTtxFWyRAXwg49FlhuGpZT6+AHCU
RuAJViJjKkpnKyaKo9WzW8bjnwvwIvMx0kRvVvqRQGS2Bp6IITT+EtIakZoJ8gDv
ZAAOc9VgvdS3IBJSg61C60qzpJxY9WhR9GDqWQHqO7BzsZVhSP5WT59H8RcMkcyj
BUIINQVgt+RjINDSl7lGeXJpVEAAGr08lPO/xRtecFQJ5lN9UwvNdiyyR7iuKEOR
bwFCaNzfmM1X8mJOHdByGdYEzq48XpRypHNng1IPhG2MJFt8SRZY1DO5E2ky5TeV
S9CO6+OHcBbgvEHopaM6qYP5X7+/LEsSS0vZozGWWADvyfLbMpzFxU6hwglySCXk
dyDrzj4exE5z/wwOrhB/TnsJ2k5Aud7VaJkAqu1ewzrUVHql/voK56MSNsiEtXOy
9r8FSzEqt/BSStOtg+BmwCCaxH8fx2CoQxAao4HgTJ2XzNW2XYqbXFUIyGlx4vXL
mfv2S0PKom7PnNnC0EhwUnWmnBG4NlQ6SFk88MGFnlEaxM+QJmqXJSuLMk3shRpJ
O3sBt2KU6BHdvF2lXGzQNr+84aNAvvUbrmfX+F9qazI+udkWvUT8nZUu8rGrEvWz
9uwKQG1zT9egi7OnZBzZrJQFq6ANX4enDTN0em5ucUHfTPZmN32PCva9aP5axDTY
m8fYHwGu1fN/itzrZq0tc5WqrkWKIOxHmUsCBrmmWPmjtk3KQ/SFCRAVErH4UFtJ
fsZ7FOHQGrUxBH1xnKKf3LV/4EmOqT1hK3eN79Yjlz29T46cvawTJyj66zcIwelC
9ZoY5ozMRmxjbF6Frss5OhWQnxQ6yMyDaZ6guJO/eiZ+l5KYv4YfCYUJqcG3EyXz
Jf9V2hkKrVvWEQQPIZeJ3zZDrJVORiBOjDxujnPhDIOG47v2TwO2f6QRIRlSw8e7
Mh+JMvunRHHANdIhSbC/CT2URPeu8tXHZ2S8Lw3Db+Oe5kD479n4mU3fNMNQNRFj
XOqyOphFt8oiQOTONzcKowe5x4oSQ4Ci11Jd6yUd6B+7sWO3FLYc33Gcxzi68YBm
SEmQcqMW4Rpu/uFewiaqy9yUEp1N8cwvWBU/o5NL03M01zz9pWdFQXIwMBEhe4cS
1U+yaeh4l6DLj496lAEtEXeGYYMF1BQdqXakOgQfiFa/6vIzo3sQXbyXDuxTZGlA
gKi3N6xxEnasHHN6k5aqgZ8hu+DG+dAwlD0/33+yfrmgc8iAALZXAL7wl4q9ifOt
NyPndQqQQKkbdRfQDr83wV5cxmJ4+cMVNEKrUl4OIlzWGe/i6W+NH0KadK1m16tO
wUWZVkVOwkIXGjcV/Zx8aJoA5qcdIK6dsTqwnnWMijxVDmClRDnSucYMrZW13e+1
rya3fVLDM9kZHELV1wm2dn3OUOgcpKPnf2TbtTbPlqG57Qh7V/coriLkGl9td2OH
Z6s40SuUAUEhud+uE9CGn0qespYJnXZH49cwgynISOTHR98kwANJ8TqtjxNHu1Si
31Ejk9cMXC8L3oczASn7a0S20xCj5WOR9sEqy5VRlzF8J/tarqufhM0sWOraSLSY
iG36lcFDCc8wI6iQIbw8iCSl/SdmRb0qbI5lV+u2ttmXI3aNfVyvIUqjIvPkpHJO
fio9lUtvb1U6mp/1IFJZb8NtAiMV8mjTgZpSH1RGCFIh3VGwwftHwCxxmnYRB5Yi
VYihSJ6OoMG55fiheNP4pxhjNiBQGd9MnqNIe0H9bjBAPNDk/IWDObfbp6Dk0pd7
2yADxJL69Jy9Iw3MlsPpIrRMh8yEF12kDVL3xs+KTLrDSD26rzctLQcju7+0bARD
PC/V6Bl5HlO9XRSRZcopwBI/2sTm1rcLOgVOAT0j6R0iZMerNV0iKX02gNIa8Tc+
AXghN0ZazDVSZL6jHksqEKUGOSMkTGh6yAFuk+2KoG0h8E9f2UeXRGiqprSIf2pb
I4yoQWMZigyZR6n0C9H9mjsqHCQPCG5s8XpRPaiSeH68+MInKwhVLvEIfx/8Buu2
BByPng6ZO+8WxXCvVUEKwTqNO8DumeNYSowDg51crQ3LNG/SbeLOTfZ+mbdTCmu6
iAyNYqUeGXE0N1YQ4jpuGY+36FjpOAa9rYKus1e+uvm6s/ZM2HAyEPi7mTCkXjsj
ZSuAJxk9dg9KbAwks1L1H7Ct4ocLerTDYnRRRcECHYzLCPIVl8hPBe0rQP5dbeSX
Lcm3cVMjt/g01BccN6DJggWDGxlz4nfvyfVif6NcEiBh+HQvJB7D+CBvq/RjoSgQ
agujBKVsjRpNknonj5AjFPu6CHSTLUI5TSAVtNtlGSFOu0Hs6DwQs2F+/67yMYsC
Vz4e4Yjnnxa+2xkItTnq+StUacdPw7J1h91gE+jMoueIoKcKF53aozctqElZR8t8
cePReQZ4h81B2yjzgNjqNZIHhwSVjDTZsmfLcGRTpTpM1enOIkG0amwqip88LRpG
GXWcKejAmKesflCdvr0VDfBxxUz5EKTAL0rZu5rYZ1pj3qsj6/6rb+7XSI7l5Wib
ZKP+T0FPDoXZ0bVcigsTg+ZNT812dlEzgT6lUlBuaOzuochVZafnVt7SPlNdViDy
ZOinhLfRlICAzGLcTCd0/C6QLetmpodrmXLr95C4hB1HsWcrkKrxX9CIzzmWjFe/
Ops6j3zJpG0C3L90c57HHYHdF9n//sy1wypG27ADxbTlthvLQgMAHJPQXrGCBGDh
xFYHsd58ncZIa2nchisw8I0bRU003N+eqQ9lRXvA6HLN5O2YoOL83yNjVMrsabTJ
hfFbVhTgrYfbhiQA1O2IPoVNGngo0DY63cjuW6Zqt37EuW3Uzh7UPIbnvzbJyYOE
NAYV1JHsFe9Oj3O0hv+h5qARE3Ct8EWLB8bFfBMjbiPQ6OPOyyNwfR586nRup1JS
CbqV+O0fqSUaq2ntEjTGNn9YGYKZZouCKt8zjX6fg8FNrgv2Ojo6TPCrhvC/2Hll
/nJItcfdMDBdNX24DZDLD29wUL4vcjFYLY0bxueXGpo+2ozZbZ32wdJ5iDXFMvCc
OCi2Iwl/+f6ktWxXk30ZgaFG2CDFcmjVPCmovAO8uVoQZnMExB8RN/cr4WkawNy7
qhNkQ6AXUqLyS3HHWyDyrJtIYKZZj4k/D0imIB+57FMC0P/IXHY4BJZlR6lpZ8o6
CaIUhM4E2MuHbLENu2i6A9w6W80GxEIco5yr/Y2A/xRw0fxj+qm4hxe8P++wk57W
wLCwdcYTS1KI6iHohgOAZ46sA7WaeffSV85032Ie7POAyLEsyoOittd2jfImW4Ra
o9kwTFenQmevHQ+bNoYD83qUiJql37/NS1o+kb3BcuK7rcxd1lvPB8Cd6CzmDZUB
6g20XN2otRtP5+emFwG/Z03eGOrP85Zq9ZW7EqR9Oo2ziVrz78y0cPgzr3kCmvOg
rS2NsGZbu1wdjs0pIlubMl+OdAVybq1HceTWJ4E67BabeT497RqWRImEBwmS93gk
610hMRXAvlTUjgLBEetA5kGhiN3l4N+/5M2T6h/+YMzUT29iLKzWefIIxaEBLeKl
0c2sWkf5NLxaT6sXJVal9q5lXMG8aQ9ys61mc3jLczwQehVublyEbdZgR+BzPdaR
QmjLSFNHog5fSYzDoMWGWYcqaXa1QbAhtqbSL3y2p4PlQBw36YSkcFzbeqeOzU0e
NwGo86LtytRylCfGuqtIi522KgH04huTlT7qx9sduOWrPXIhlPlZBPRLmO05Ihj0
wd6+W/Y+3v5fMDQGEBy3bnM1dBMHiOYmMzQ4/JRircqn1s0ahAbFJZVT+ZFzp+2a
7XWWTgF0N0CbfWtOC/g6+60v8TY8bhAf9sbDy0I3RrgkIQPJ/KBaVi44UFHGb0k4
0GaUJ5F8zHnePojMtlFTQ/tUkm9OmfGHikO6+ID7FllYOL7qOU4YSXnP49w9nxBY
Q5KA2jVLNZBnOd7BcgNX0Mq0inU2n8hRyKtLi5SH+teLC/g724Jm3ddg+zGGL9Es
VQkfZVmrP65pgv4aCEDmuvUFxoUtLImBz+xEHLHJUhISLStAuaV628AWlNM3zA9J
8w+VuQhk2UAD+lTQg4QsVhzOLdx4jf4GZIgFQPLikpzdyb4gxEZAkgUlV07cIR3w
Mot6c2Y/MBRMl9yow0d9eAsC6KRhQlI5v/1zdQLr0vyEsaxhXOZ1nK7YaTsABJju
sKxtk4TyhSoEtCA8j2VtSbf3zddX8aGPZHIlJpXr5KcWa8Ky78cr622AnDtw4j/1
t3R7Z6z31/kIOulPW3WEi1Ib4Wroti3btEIjwxzljfJYEYzbvKhpue+2OghEYq6h
3zYXmIPucZOWko/RGCxz52J+2XbwsBsmTCrL5Um9O0hlM5iyvrq39isPPR/dWgiB
T1yLLC2qKYZqTzTo/PkdV08nDSFs8c0RkDQh5voGGVqnJH+vcJY7XqI4KWJH66GP
AbdfSgAQ3qPGNSCkAe319GDXpOZ/1KCmBbwWZPcgNVpv0C1Js8WcCMOcoALuT+hz
VEY4jV8xhuny6S4ujhydBJG/lfQ1zj/JE6oLzZgOczos4xInpWHdeIDLWFlKB9zT
0DHfh74UMbq7jaA4pjMFTuwuZtMHbQ/hkMKIwj4WnimKxtHNmkeuQ6NH9oxiKK9D
yDWle1U6XpOSKWI2Tix+RZiSx5So2nTj5fOmUlgtAfpplLcn0DPnylOEVVLmBep6
xbBbI2jcnqBojZGV88s+4EeIdAUVyny7yigE5M7vRWMLV/bD79A2dXTQeCBca3TY
w9X+s2O0M/UXc5gzs9Pj2aFJQjry1DruF2o3s3tL7OOaxSpuqoAhgcMEDXKW0MF3
9l34Bze+rHCtZSg/PKQDEPaZS5/z40vjvBsZ02z+AsxkV9KUUJKmLGj6eFAJtSRK
Ndt18SJSiPTt7KcMiZjsrOkUyR/hTwdH5aDLMjmfC/59NdctWsTfu/oHdYX39xhO
SKY8rqmleAEo63UZATL78qYSXDM7B/XVpcTndjwSylXJiTof3KzleXWtgtDQ2Kcx
IntBXCnrckNvPGc22AUFM6kKUGc0XwqSYQnF4Suw4pWDO3w1TdZwxlDRbuf8rjeu
cvCNUGl7uFO+m3sn67KKbfQwjoWmAhSuEtQX2yLEf91A3WBTYP9uPxQkYmfCaxtn
Viijmabn7tzIKJwdd7pZykYiKUXPe13wcHTU+eyzDMsFibu8totAXYQDi8Ye+SKX
2mfdsuuOqyenQdf/tK/Mddp2ig2QR14gXA2E9D4rVDahD2qWca4Ptjuomnqe5f16
JE5xqYGZkxqaBCnrxGa7CoPbflReysNMDHpxs+bDm7BgRWmpTfo6vzRZsxqQD4+m
TkxBKaCh/21Cv+dSbcsrb9KnVzlYK39xl+uL0BTYGrmwT132LAMOMffJ2smrT3/G
w3LkjmL4XBhP08AGoPhac2JsqgnzWRb7KdFHIDWRvXjk7VJjgy3fRSOdSzaEMidd
8ave64kJxmtQfMAVLqSm+TjpRku4L48E9XBZhITN1tXXzF4XJKocuOmxkyf6FGAg
eTYHJZ1bPUm5SbaVKJQXXoMIolbugS+/4mWmcG9N/oYPeIZe1b5JBF75HNg+PZ1n
6zBBhe2WmHyas/TVqDEM3T+VY5kf1E8fqLkpNaX6AAuc31igjNj7n04XZgVS7Noy
SPqNbxIYONB4e7b2rN7hMtIuCm9Tpg5VXsvRcUy9e8eqDtu+VfeSXzkS/OIE2+fQ
1ukjnbR8JwA48sy9ZLl0U2DBzUN2pOYsNVfECqU76BOlQ4Zbay/vE0Pklc67wRzQ
wTdO1ltA6c0hJgvwPZovjsnPFRDCB6QO9WcdJrx5Ouln5J0QRFa05xQnbDeRVtcd
66MHcEFCd0q369YlEU2AjLhOGVoEStkIYz8nJ2Tfe4JAEJ+9nD/0W3SPQ4kgWCl9
nxBlncM0KpZFoHSgUSls3XBW9zuawBk8uYmzbnPPvNcOxYAprlZTc0mCnqvfC6zz
HpWXI5DxW+e95eeTcAegQIu+iAtZMjdsP2+k/fPf7tvc4mCStelbJE5tjtpLnXCo
PgSwNKkZlEX+xm6sLGR22TcNk5NwgNSNx0EcVrmKpBNVjPN41Tfv7I6R25ur21Ta
nUTnlXiT7h2nuyvkdLP/u2CoUnz7usWsYWgQ4cub4vdCg7wW/06+67IcCkwWdvsS
8TRHBaokoFL8rq53hFTKKYL1VNAP/f3u9PiPQlt/diYNRVWPxLh6jyWzNqTwBmcZ
0LwpgjXa/hpeJD6Q8eaouFa4a8adXi4XBOoudBHmu89nhAS0gUmtyvu8RGZ3hB52
L8AruQfqKjLmlEvAriwZUKX/oRqhXe9UJOVkOoZHj5a4GJVSiXI3uVa34gmJe4tX
hfKPKWVv+aAoH2euMDS2OQOFU6N+J0Absv+hLyWAHicedjih5An7YUE199UG5/dy
pzSYlUAniUVv9ZYs6awCDpGTEmhOCn3teos51R2KgJIANQVFvspS8nbWEu9aHmD/
Q4TLOw1mMuWvQF9wB15tP9ZKV4qjMQR4z+XwoI+AfNmLX0srsJ3m1SEjnuSu8XlW
LNBMfLl0HE96/EdHZwJirbhFFzupN3QulmF2RtgowOB8kDTUjyy1/Z60f9DNNl9i
wcPYfmi2Y4tfydfYHxM5G2UCDNMaNEv6eiQR6JNS95EZCGdGfJCUA4rkewQcveG4
+d3kZ7sd8neWzWiT8wLa/l+4MpNYUYxOqM0ddbyh/yaOBdnZIiipndGAiRU7O5Qn
AlXoEixC5JQeKXFS6zIGuVW3tSX8SOr54/Oucrjk3nIm3MWvceBsNJ2RTlwEUvx+
3QL3KXKl2pxWYKC6elGA5iRLKLwnPds8xUu32Z3pNFKg1ZQyV8+kTFeoZaM5IGj+
7U4a7NVwFJ84kdFZRkdR3Pp7+sZw/M02AOMA5t3luRzaRdTm4xhx4/KE/roVHfD6
4h4JTOCrFDsgS9Xpn39oSJabavM/E7BPoW37yMlhihVQNQ2jbIIbUUJFkXbME0ok
5VeE55J9t3BaL4ITMMbaj5BOHQCnbFkOiXOm4L/DMitF6XRxMPBs9Cs1eRxI4BE7
XWpFjHlF2dPzl2ZIVAr9hCRnC2NUqzTwzgkkfod6GLkWnPeApdwEY5KLHmH7Sqir
SW7molv6TAO+beRkjtZp/L8GPW12+JbFC0erq7/hRNydgDp8sFJh3gffsdroJG1n
x+EIO0GzaUyYiFMDb3s2KQZMV/ulQ7XIL13WJ2Y8SFXn5Baepffbhm99GDxi2ReA
6UxZ+G6ro9jU7e29gUAK+n09IDzjCEDD7HuQCn9TLbMN65k/H1PXV9lcZlIxYvxk
NmqluKxHryAAfspaiPG76kUocDO7qF51Atc12m+VwJGglr4Wygc7+xClEMVYo5Zh
oJWscW44RddkLiMfk3aOyq41cHzKgtbF/tQKf8iNpy0RjiDbWo4pV1sw34nlNf8h
nAuBRQ8iYD8dS5s1nYVOQAQSpD42y7pxjYvrDTqCBdXFLcEjBIezDpZlWnweojwk
hvDUcWMAy4aYcgU1ffpDWjQyMPldFPfcd7oElHcX0rHj4Xf/i49SCrEZ57KSSV/Z
FMI6UDZ3ZDNkg5tqQL97pwKgGUVfaQZTbo2YUBv9fBULz8DVnjz3kRpM6rmREdut
NLojA4yqSg8/53ofVxyPfuGWlxuT3/5jT2UEU9MPnT1SGM2IXt/sJJ8ofxrrcuiq
LBb088hMZE+//OK1lL7DHT/sqb2/4HqZu8L6eOdlIlnT4RsVhZ0kFmzCm8qfdxkB
UFOoncwuaAGUg18PmMSPADUhe+uuzJiAsxBV/u6oOCZchV9aLQSOJDnpOtC5tIlv
pxILxPIh5kLIfAtmGTrca7hRM6uDNHMkAuKrtYnUXVlRQ0n972U/YehMYWH9ZGNB
PgrqtaOdzxdg34W9DugvUNjo70HuOfqHFC5qNtc1TNkfQCPsaVPNHd40qDC5BV2b
iNj5DfCzaCEhjBTSpiOqYe83Ogzw5+izEKINmUwAOMGf8At25OoPZ2+n3P104qLw
X8H7EMVt2UtoyOVmG20zhw+qR7lmnZ7j/FOGT4hL94ZdgItcSC7wvPGuvrCgYowQ
l6xlApYcxb7kOZ3HPmwAjkmE8fMkulXI3ZWB14sek4GPVOLQreCTesLe+GGVjANV
pw/87c0QTfwk2kequpwtOb71fzIMLQtsSazES+wRlYe5dVzHmCyMPDjREau3uw3k
SQwpnIx5swpU4Oi5TBAHGWXfXyHGIz3CgNYlSUup1S6Bg3r2efy9jSyiFFCWcDFr
c0lc6Rl8Ciqt4j+J5YiSVmoT1vQtxGkUvt89xa0tU3csSZLUvMGq9dXT+KgIgTH8
M2QvGMwcPBVit8dtYlK+4So+qXMxfyDBRSt7AMV2s564GRQ9HKE2RKoUFeinLHKJ
CWzN+ulRga185Vi+HFiyGYPO1dN7NfPU1rXhbGtCRdrCh3iU6/PFY1DD2zJ+XyGp
NoGEXlrb9gIAukbVxoBZ2MoJ/T64dSLDYjHSgZpHlbEPwnL1ChEwg8Cak5IcOyjm
FiVjNxqmSqhvdbJZd2CQy7UFhLc7nt0fThrcuaEbksFmWews+iLww8CXdYMWylWw
ylpYJH/h9pUQtmsOSWZmQw0MJGZuuYOvjwaoIkvHzmKegN/Vs5ZIKtcDg591MyRD
UWpdMxSyZ4zFRFk8wEMQWYB9aV/KjsGa3P8tdHxqCEHRSH4P+m66dHNIUsECqqTD
0J1wBP3F8Ugw6+r5noXHKqxE8weWlQ2VWjAxQ02+w498hn/hJ5p9xE5nFZJYnoNJ
c8cO9nypneZldwdzBYSAvgqlmQxuUw2yB7SSqCVuQ9aQEPoYwaUv60riFpQXqcKH
/itZe4II4p4SuCxURKS71imZYyyHzxY/XD4l6MDBKXqWemujQud/kLgfTXGAL2bC
/ga2mPy8zyrXEXTxyUV88FtKHVGSNpE/SYkigzQmTwLMsZWAEiW+JqOSmLhW5o/c
pL02yjk3zkEDjHON816/CxXcm6XLCK1ICpoaIk5Cy5ZaDZdvGeGo3HRIHN+YiJqo
Ubwh3PcYqAe/7p+hHzyaNLHcxAA3EsXkch6t1Sp4+HJ50V1gGdxCK5Pjc7Vke9Ot
4hIazeP6t5GYYMpXZOKLTBnBpmbWx3kea5nItKShOSZt3Mu3U+aoHZNB4JDurdie
tFxEG3IoaA5tUrd0QG1D7z0UL9C0Y6JxkYbURongKtqPg71Ww5kRKEXiMxC+oVjm
A3rSzWEnaLoOhBDP6Ii8aY02GsiIuUpP5Kri92OyuI/BNtgndqRGuXKeC6a/AbzG
4Dg+vUN46jtRwQU9at6fmA/5kXuQwbFxgHegSK/Dt7adnwd0dDic+LQUH15uphFP
uOmX6Wsrbv/7friY8+ym5ctjeON3XUQrIxianCwPF5sCajeWXP0oBWHZvjqkcjK2
sRAZuoNTJtK3wMPCaaDEL9RfYL/LHqQXcqAXcmyc89DQmF2JwzUQfj06Z+ZN+Kxb
5GtCiVHEe3FGn0SNievSVlrwDMucuh1xmufaLVpSaD/K+AgAb/h4NI5LUofjEt70
3iwPOeGdyOT2g/VuNtDPlfgopivlXx4S7Hh2ag2bqnCsO3DHUdUrru+XJiumDqeF
PVrydCSX6XLRHthBo6SpOAbi+59pHEljyX/rWRiCxvqlkSyvdnTgG0mJNlbSomlL
TlQY8dFtsDD8nAW3Rs9D4iBOMCEMgNRDJfq3+X6mAnwJJZf1+/NTL8OBuicXas1r
IKqF8hgfaIMcXLHyAyKGgeuBUX1rZFzbkZLpnoWIF+M9qcjrgXqVNfumCodTn9hq
GnUPI2mMzAb+pJXQ5g5LNGTWS+dTGKxFizR//In0zXLpoVtsWEQBFWHZQXwUCSRd
idK5yzqOYyXSkWWCLlU8XmU5UnNz0UU9Rl2ZyqnwfTsuboI/uTu1uKaWc+gNkscM
XWbPjh9eJqNfq51Ugnkz7e2Ny4VlzEYn5enwniUv5z33Z0dJCk7FzXTc/LfL0dDF
WMXAggRgbNML71qeLj24a597UpUmSMobsmM/WvvtJngbnelNjpfzNCwRwU6/WK2c
7j3Jl76a2tcQ3Osy5otsy41rnQWEd4aYwqKobj6rybj7hqKMXOg76SU8JzrAliMM
NK8BYjaTdFTCQVU5hM6eB3P0nGqwQFqfjbMzyAyCmcbxkVKx6j1t63V1J+QHu6nF
oRR6ePq1p5g45u4IpX+G6viZ/0sVsy26lyDbKL8tqEFT2arSa7zxD7PGoktdo/Au
LchCtlLFeLThdi0j82LL1Nsm/RbhOGRo7oarrXTmB30u0jyyN8j9tZp9oVZQgqT0
26w399c9tSZX4RWVqb9e8QXz9wIcFOfD9FLkyIWpPWGdCaSQxOMBo3LnaH4YCjZv
TJA7x/JhCTd6ydEAbbiDM1LgiaAjE1FM8HkAKq96Aor5Jj4WiaOffyLUI0h3QpHe
WqUstunMvTsnhFOwDrD/enGDvdypepqL8uvKceVYlQ5FFWOkPqOwlqYaTtiZagi8
RKyf2EWix3y7Yj5YMJXPjj4F9R3P6YTRQx16ZaIKZ0MkS5bjukAoGJyScgvsx8ef
qOa1qzjNPX9s4lEW7VjhcjqlbwLywlU/t5LiS0Hs/QEWcP0lbLavHiclNG/qKEmj
Ve9W6167I3vlyDqGtQgigqNRRxvT+xqCo0EmseADy0Kd810wU1ywDv1jLTUoqAN9
9LuZURQi2xwXI46hDv+KE5PaMlj2smrpAhU8BSLhWDWaG57cDVBLsqlUPH+WXK2U
dsSRYkf0ar4DK8nk3Y2PIOtUm2Ky0frfI2Ib0v/h2uvlGq298WWZaiMSxhB17O2u
4QmScnE8jp9gCDoEdL0kuXfuF4NQtSfpkhfBfCJRgWFjhrk35kAO4rF2m8s8aQfq
yPzahM29WSRpk1flXHZuI24RUPJJfsvlxnsLddbCuXEAjHaL5SXqGT2VjlzuyZbo
I/UZU8+OIyHw6HRpQf/OFWFCs2lQxVKgQUJ4lJm6ugRDwk2eJ/0VDdqV3fqLw+xC
IiQW1HoUp25cqfVFMr8/y4DnUpO8UBGKIeShLIplp9xHGzjghZAAd/Tl9pIXUjUy
gmGprWIWmoTHWKvlg4i9Xr43cveC33ygniXZ7QxwKNoKpK0JKWH48TkdA7nlyOm5
NLzZhecscCHfR8gS3Ua52K7uzUzmSe9OP/DS8PIWdoHuyxXOOLhxR9hXbd/1eBkC
KAG5HkIdmhHRIuiLj5/6+g6Q0Fx9fbPdtyoHTL6VAW2Wiiof1rS4HLNAuXfxSfjH
UipG5c6s0f6y3PIhcyRJLUT/8cOwhhb1NDFrHOjRAeW9qWfq0HpXNKAnwYY29zSM
LfZ0NyUgwA/sgJAjgxflck5Cs5r1rfYjWFbqwuhJP6/wc6y/qkjNFPkgIW91lU/M
5YG6SUjWjhXVWV3GbFprpRcLxJ1X5p5+JDwQ4qtmgQ5vscyCkS+OUwf4PPPoF/KI
tq9BE5B7sBeR8sHmlSC1D4Uh9DXRnnm9jOEGhDrXIe9dYK+Ds1rFSllhmD/yoeE2
/27Q6rL3he0jzKIa00y2JnHIOzcJl3pAeVObZKmoGzv74OM+1KfYxIjzj9vl+zjI
3J8a4G2vUlNiV81egjxbTTxoR3b3XnYTUvL3SN0hyl9Uo/8kvJ3/1B6SKRcOHJ0b
FGaBkLajWvm5Pyb6f2DTjeun3WcUFF27YMGtC0BpvaYA5TVbJJM0jML4ezWTPZA0
/dlMzv7pA12KmbdGcW+WgAIZKjTYCDLFHR5XHCa1mriDsO8+Z/pCyVglsw1xih2K
LH6GVSlyxWBtrAGga8KdFvZdfMXGgJBsKNJAyKE7cGJzX7qKHTcp3l9kHhOjmOHH
VonZsihknqKZYd20HNqkMKQKaqktna5njOPTf3jhom/7IbH2ZzMssoZpZzMYh6BT
QWRjiAI+Fes4oZer8NdrWegyiQc/jJ9p6l03ODDdCbJDOG1sx4H/EgGOXLngphud
l/ztpulPdBnrXue0n2IT4H9gNlgQd6Kp0u/X/+dhn55GGAeGplI1Uj8T+moCxpEN
W9IDAJx1klnfaCNuWZS4bbRq3rYplR/PAtdGZcjmCTlSPJH+bmgbXRFr2vaF2pST
Ank1sOnrZQgPH2hmcbT0mETOBXBKdHbKuBMNiTxRsTF9N2fUc0ArnFwJXkL8eAmF
fgyKC599jwTrQ4IV7pR3ais5HOey9BABH8HPi7B9PDm108GH+7LVJqsaHvejjGSD
bDmdrdXZE8xAjyOvhCauwLJo8WK/4Ul6AdjNwlLnjGjNChafpcIwcTgPYMagQ4OS
PL6CH5dQjh1rvqBKvkyD4q4D23kPa3TJ2JwZFof5XLNxm1crvBHqqXG9j7z1g97/
ohrJ91bcXcq+Cfy8gGAoxMMr4wm+2ZRwvNRuCa7JtxmjICrc7UhvqUgXR/wnvOTn
gZPZc4SqlztGqzwXSqcQnCbsfb9pvA4C1haXZ+4C2skAf/5/4uAFPgzRq4ifXEch
gGWXPhTJOgXzharbsw2pqDyn9HC+gHKbWx/7ZHyeb3ydzdSsyKaYCZgqz1KWf9Fo
ie5UWpTXZlj2K6bQBs5p/E2HTjQphNTdCAd/Vx43ZmVuVqis7QjHfUgg3gpwt9Dd
L2zeaGqYhY09bbcDezNbTmg/VAIRIv3vFnw6FTKkl6AgqmzqkPBWJOufyztEor2i
tiW80wmz5lWLSU9VnO9cyKCfUa2wTPKvzYgOenkzLaw6qy09ek4ZAaj1AArraYEM
xfXPS4OAiqHIcdwrT9MIHxlEYMoyx787UBoMhex0zNAS/GacNvd68yGxS344bJx2
Bzocn5fbhdUmXYT1Pw1PBpIEdstDKIuCejBN39fRQH8J6DAGygMLF+iXWvxzjgHn
8xK5iEFXx6GlpQGpmw/Dn+gNPFGJEGpyiNAiPPYh7Hy/xgbBZMSL3CX46ot6WVTL
OMJffotlW9ngZ8EJId8Cs63uMA0/KQN109/37HitU3E463VS5t3+DgdHFS2jb/UI
RTA6Bz25VA+uoWMhRRvtBG6sz3sDt6MLjdJ/pGqo2zfyHuelKoZl9V6V6kgscbHM
LfBNvPIiN7VLuwbrSaCxBt4Strjeayc+cqfhbvaiZNWKwWw4lEyP3qVu6NJYwIDo
V4eEIKpXwdZ8DzZCvgIxn5zTj2IlO3WVW56RZ3HYiASqcEhXJKnKhaWuk5TU19xo
VJdbvP2I6or2CuphyjdqLVl3FlaLS/JbB9GIkBv1NEcrRIdFO1gYCy2Bq1closDf
W708dKUD/inYrvWSYptUpqx+A9Hu1kfP794wCq6iE8FMEt3jAvpQ0nSYP8E1lHn7
feXBNysw/E4lFWr3RAcaX5u8nTcQxh9oqCrPc+NReMXSNirPe3L463AFqsX9e2EP
lcWC+4yr7ZX3E5WXiTuquNFHuCjnjX+5qgWGSZZjTCuIdr8Bj+MW/nkt8Nj15v8y
nUL4G74sakb1CgMYfPO9nMRVkDGmfpY66ulA7hNMyD1vXKwGQfTJujeaUa2BcETG
WhX56EsKsN9bp8UCoOPVBRVfNbept7B8w/sudNKs2aTLMu06QWqp6N9//IYm270G
fYH9nzQeSq+ra8AtAszOD+CJS92bhN3M57SAM7LmvjGoi4FysullRmskn2fjekCm
PXUoVvQSMvVPNbbnrc/vrjlEitkztcqot+XJ0LzcFKVpsiYl1MfbhwFvJNErrjbg
MVukd83zYDWsiSdldWMfVl+lxTG7CWXex/HtGclE4KZr3O/oY4k20oLw9r0Tjw5c
zeXVAVY6z/LP//MiMfps2WFneTVGG4pMWNv4usTSl6H9jGK/ymXJGSkANYqPQWsf
K68PZrP3ysH7D3ltO+Awlp+9HI+r52BJb50ea9FSXfzZdgIYqk00gqJPgEY4CMfx
0md9QWXcT7RcHtNVCSUUGxUK9+g/tHp7UIPU00aVkOHcMCrFQnXgXzmuON2u5Xf+
XLTZDE0wslQ2wnLhmKG1jsnCKLkF4PG9tge1brSorwvzpr+ZJIxefUqBIoGPBj7q
GKwpAO6cvBAL2Ri/ULUdHQqFyaQ9ykN9u1eAdHmHze21635v2/vwgq5uf3s9LiZt
A6riNyLKVNFCSp6wVrBXLwuWH8xc2iFTOe1WvgHqPwifzoDTU3fCaeWUM8FUNt3H
lhM/MNFLeoWfdJElGwR9gsnVCMAp8VVmMISwF6o6GjEUWPQelnIWSO4bh7skKrKL
QpSEHMhqJ3XK9y3ON6QYSCyrUHuJRUC4KXpbQwThHVEhXS7gsPSKpfUXYMVrBH/M
s1+6P4HXJbkBKDf9g3XyDj3K3+sdMuX+8JXE5COc+rxojzw+8we+VH9ve9KRVGzg
iBdK5vn4IeQebxYYZVgpcQtRszqW1dVIw47ymEkWHSlaDhHekQEdVF9iv/IAmpLu
tvRypBUnnBcSfrN35Vps4FYKNVLynH2Xo9Pt5/igSo07+BtSwjZIzkrffeSsfq1e
llzjiFRN6PhikYcHjNhKObBfj9lnDlWiL2e0ml7YWoMkiV2YmAtnFGYPl+YN4qZz
bt4GhmXiPCWbKnxVPEhRLSwY9XprgcoM1yrB/BSy7Z02v7cjetwnHHG9SBZ6fZz5
rjyJAm/nsOM0jUPK23rDdtD+djYirdkjMFdZlw1qPmskbzyYYeoaTxgLJbzGtUS5
f9CF4/aAyRTYqL5Ua9qYFCSFncw0wSkY9iRCwp2DZO3UyGWB0IVXefj1O8BsadW7
4OMt/wo/HwqPapDXVxG1fVrLVyq5AUiFXgfwVGL0AXhdOjG4eD96Z8nEDyQpQZVx
iy3Eh6KAbxud4X2NLhM3J57zIkk7wxUOMdbhyMUiYNC3TKuqLOagVcWEh6QcC70L
e4hubV0m0HVjJEHOS0a34k7FMGUk+IiTL/n1ZpQz5jt1p6VWR8OZjB/haPVWq+qV
qfJUiQ0QBsDXraKFCnznskCiFBGE7rkykZQfJKk/4R94mDhXwfPoJDaJnajK/93z
dYmelxrgL5t3cZZCKL2E0kTxcopJ1bBihcHLr/txdkYwSN8qfjBGpuO8uaecOtZ4
Qq8Ke0Xi4BbzRfl7BAFmA+5zsV/3Q6KF7pwVqiA8wMuEjpDD3bYb75MZLyFErDhZ
KNEFLjGPxyKnpyOfxqBSHjkodQbZPK6MWWGHQ+XexnP5Mh2AHxXk0O1UVckikMTP
ZwEuZBCiGFtdHG8qDQ4F3dZFrH/YWILcbwl3UXguh8YB70YO7keFyJ2aF4bdslXU
gVzhWEEItllDoUyIkMQrXkJ4ugK5PbLOZ30HKKTzzGI/UzYlfFGVGvRMB94HTuBK
uCYWfBPADcJBqytGW55mVaGnBygmcxt7E3FMVtodYafaFzDGZvj6yTv7ONngYT4A
ZrL8cSYPiune5bCaWWoyEqkpwd7z2wYi+L5HHhYWvJK1cAd3qu6nAUxYWg6ot3KI
IUIs3P9iXd3kH4aKdIeuq++IyvSjNSPAZle13k7RhnsxgcULGGvldpMfFYB0ZcJ8
SA90mSvb3rMgqtXvotP/vefBBKyHMImG/SyAWiEEvlpDNl5ZnqXiRBNwJ8jGNkQc
Ee4XfETp8I5wcP8IaJEIzEZIUCwkNnYaGGyR5RVTGxcsP8RYMjBxvJr3fVpvDM3N
fydJJQDg7DJ/SIpZ7f+MudWbwRIKMfKX26hK0TtGHHs+auqvJD3vSOpTi+nGKSip
myKm7x9bb2aVTiQfDkiDI2AjmObQj/HBlATnP1X0bbppcBU6XKDOMsRxjJGAAoS+
75qQUucGcnhifUSA2x2BWis7tyy2Fzq1UP/lJ1gptQltAX7/G/HkWagjQ+3mxJd4
0GujDaH5zMygokzREzsKEEIiLAxW1FaBlhRPhckWGyXASAjbRiWqxa+B6wjuFKG0
8m8mDApfISpaD1g3STF9PebYRvmKqDDpON/Ru0ZRY2hy8VxPULazhFHd4mTgpvFt
eOPxIdC9j4Mg04j/IMQdlszTi5FLgd44rHdoGu04tYDFBurV3CGZ9TpUtwz2P0PW
FopGcpQ0KK4fUL3jAMqDMpxArLqFPqerh4yZa2gYpkpxq1mqI7NqevAJ/TwpebLg
KeyYMfBgLC/b+wY381arddypgmvRGBICkt3P+12ZIZvctNM0mJoRaEQv4sSw79uu
gZnpNqEt+aTiCP2lg7QBG+rD55h7P6k+7lbHYa6sFkn4SWjKDGSsPEEGQjyGifA5
WMU3Ryo+ts6y9J13liXrU6O73/Ov3+/movFkJD2PLsyyhLB57J5yn0DzYQeQgpe2
kd8/GLv4XJ9bY8FQzx1y/Ueqi0W5qV4U0Qic1OwhZuF1UFEauqnSr7f1204tkmK2
ng3a7U1jI7RzcC9yAFDYjEPfd5BsG6EhHn8n60xF6vwWLl/ikQ4JGloH4N45G+RT
8BL/n+wdv2o0P1AEPIorJyl9YfoZmTQKDWcL4xUyqWXSTEXGBk161bFOvarvEefd
GdMazFxToq2jyuxPftRMXj9h3fj+uCYxSwXY1ZJESKf3QHWeVyQmuY1J+DJxOwTm
SizRRDkH0VxVfb0xfeDdMqgwh1Su9O/qUB6j1fMlfhDKdB0FEYpw0Zp/mLGCJ4cd
ltbvNbS+Hq0n3UCzqLiGQdegnCINlRLl6fu2Ozk9Ufv+5oImtnATUHWneSRudOnc
T+K2JyjxxOV4zWbSR2fY2YmbGkj7mLyCEDieoPwTdwozxrSfLOI939op21BuCysB
CQOsyS1OgyhDHL4hWcg2uTTZsan9ddtj6siwB50kIlmX0WlRz9JFx70NKGZjs129
HK57e5bBIXd4irlMPC6NlxPxeqFwMdWFmlrPvOe/h+yIF4ya9GHs2ZakqO/aPes+
BNPV/s6f3PVt2ze41hzkrLVznIPZlG1I6WPqC5odobat1dfpJIgR3kSC/pukQnhA
sHOk6FJ+nspyCu1S0EtFNWb4kSTIhBTBhLDPHCWBi0nBZQ0iXXu/YsZkHISJKRkY
FcZE7IvdZE/Xg7m9KuwoZq4j6g642H0ivMNXhXPKGwxVoRnfF/BYOEnGlo3RXSaT
PmiwkajvnlwZfATVrpqX0BzPcR7uUhmKCZVhe5uHETJZ13FD2quPvTMeKcngMwXo
K46dfZsHR/+7pTOteFy5KA3ny8bC05Vsj95SVgcpMqz0ainaeoZx1kC9DqNUCMN6
SrLaeg9t31uT1rZU8hRfHfAmUCg+PQfleCRmRFKeh9Wy759o7NRPdvcpu0hb+RQG
rhPRgFSSQI13LVFxkpnYAyXkYLDtU0NHvk7/ivBcFPJYwSErV8/QSHZTNukLLLdX
D3SW8tYk+SI+QhG31DVh5z41qbOvJTwaNlMhvnRnmEJJ0HAKvY1R+/rsA7xtfsCz
poqq5zQZE/ezEySkxwQPIw2DLeb54KcRVp5k4F+Jq9b0tfDsQDmITiNoqTyNiZD+
1tRSek23+hfFPJsqj90zkGLi986q9lPcZFSvpw58kRI806eOwogM4bnDiL3XwRHi
K/aVwHBBbY8p5XvObCjMrisw9grDu3LAjxrILpBUP6qaSxHkSBvdTLN+4TrKmfJT
8289Q+SS8SKxJ6UeyNhAebv2RMhv+++YiXZ+rnxP39DBJlUtxe70j1MEXpRFl4Aq
fsuGYpcMDamC1HIdFZhE+qqLS/2Hf43r0pKFHxuozg9trc0/IueudWhx6C9b6k33
jHOPWUgKTHK4fJo4uWInaHX0mI36XJDZbRVMoLW6mJFLBXhkg2EW3A4fYu2ceI9Q
MSZ65FAXnh9MTVfDJwkC5eAXUmR+wutcTh+MxAwgbPuwQ/9+GAuygImsrqvwfk5H
OmzOSgf0w3IlOfd620NtcBLGbAgULWEYh7H8uWCgrsPa0R7ZQPt95bOtBeSjCnLr
gXEgEll3tYGgHioAjt/VresEg5hMkwWT6vasDsuoAUvIehiWV6WS8egjMe6A+8HT
79XQ0spXzJ9i42x4K3unGnqQ7skhGF4FDfMLewD9VZEy6Z7JiMG7HSu8Q7JKMq7f
eGi7W/yc8UXMsj5c2gcgelF6UeinkTHChsiprMzWw2CGXR39nhGZHaDtoLUC3ywk
bi0b/yWcuYBlfl7gIszLJU/bLNep4VWWARFwx4YyK2e8yqH4ctXEUd4Wl5tZyywU
PCB1ZhPEo2honEJJ5/i1B7x52iSl0LqrmyIxO//PoAOU1vEu8VdEqPZxruESEtFY
s7h+g9+xKeFk/cZ4LJ+Wn9M/JYFJ/hjTuZgF79ApordgAmzRziJyIL4+t47+pAw0
JtBUvUBDwqNryusvRE8THz9u2hMQF6NuZAquw3BsoiDOwRieEBi3jAByFGxTA7aQ
OYSyqgEQfLtX/MnFxnk/ipYY011tDMZwCBd+AD7NTgpYtzQhgJDFC4EFNHOMfoyg
geoHqIIBsjZJ0gUHVG89iF8kP/zW30h+Rfeb/s5VPvBSj4c82WUar4aPaLAgb72L
eS1shdjLDdBRMH116YpNg5YFx+WwYcDVlGoDxuiALvw1cucS3DYl5+rYI83S4WQc
t1Svn2XsbcNEUX9DDxN1vQTIoqmjpv2uK2GIxiB4gesdFCUlZqyLB36P3466RAye
fUBTEEnnLj5t5WaB2wgCFhTJy+d4hCeOPtQyIzmAqRyofRjvKBDzJwgm6IeJqMK0
as9Jx3pTXGCLZ8o0fzxEErOgoJnIaDp2pchSGOeIbarwX1CtxjX1u8Op7NpuVNR1
VYFOHj5ToRfxQPl59PGJkddozh6tYK3KDo56M+PSncjyi/6fGQqVTykOYqD0KJ51
HpmbYGMTGJesqson6T3QUrv1JjMYVlc9nV37RK7IiOMGFjecjRZO+gtzV996tZpw
EyXAGyJhfV53Y0XXhcGb6eq0kjpxPiMcvFCx2hICtWURKP5d7ZpASxONAm/1BaHc
pcCcd3Yq6+vPuCg6haXaWZIiyx3i1S8qZWZQsD07R2twJcZ2hIjWnwIY/Ef0VvRe
D7b8IdrYkUf5uvOnbDYiCZiFAkmIYaXpALUNpX3kCfJW4/TxLyn4cW+rOaYMYuna
exSmwSoC78Dc4lk/HaqV5qqZEMd+o/uk26OR2sKtYgrkwHXTn1KEsYEzf6EuBdHC
Lz/3vA7o5LCeSXE8jca8W5/yW50JyeN5Fkp3sT3RN6/UIIUIvnoT2nPODXM+TQ73
peW8R7yM5g+NLPnlxsvgUTH8/ThRuV6NaukVzJqgQDEvibzZITRweADLC+VEYqec
Je1y+U+6Re2/J5/TTQgNCJG9KNLrJDzzQzNYgknOjDXOk7HuhVaEsOjK1mkQKXwa
I0MdK0QkkioiQHtTXfxFZPmHjJLpwMkhpOYD1rLlgmuNGuOKm1u5MPic4hIBHb/p
tgBbk5JlF4+v0q4KX++eYPxSHmISaxYIgAyfCKy5YUuCuxc9AQM19ZaruSAo0cQ7
BzYmZWTEBxb934i6avdrRQ9BU8wxWJLEqdVkvfpZSVmYY6T7XeBFEeCyUuynmP4h
OW7vjhFrr4+QA/HZjR+lWTxjw6FMsNgKsPgFNnEg6XqHbh6JZEQFjwhUq+Y7tcK3
OyjHIA6PJW+ybTv26HLxGwHyqDN9nwpHzR5B76yQZJ4zylaxc9N3MeM47Uy+t9Tc
3hSdB4v+YV8LuwTXIk6L13FsJ+mSk5jHbKZJqTePJBp6bULg3sG7BnwmCMXxp8ei
XhKgTTyWxwzl0XvhkaQGJ/7zfTyyguesNdsRyJG+0ZKbypwDxkbcWdWhd66ifKdL
3i9eoPy5L0pc20IncooAxDKBmg8MXaDFaeX4Im+vG+PZa7dgKBWPZG6U5F9IPlLO
wzODot4uX1YG26esLWfoGdU98WgT/Q6HrAbneicNAY7Ry6+5sMnvR0tAEwUgjNeg
/sU5+B71aioNMXoWHuTU8FVgKA3FK/zsdBt9XIGT0AGp+g17VE4EAmxP9bjj8k6v
tlQXcVIytbXebEbdQLxJAHYoaTRW3F+QR0oY+15BrilEhaSoekpNNuEZDapD/O2x
Pze5prtiY+u1ajKzYatPrGflfpOItb9AZQjuiqHy9lWsgr4fTea0FkRbG6SE9nKd
aikNMVlIrpsxyCRJOspZbrk7EXcu+ekPDCfMgmBA3eOePIiTJotUL7+XF/GtSAJm
O1CFeQXunSbyYDgKBABXwnBgjcZtzCXHhwuWRFzvoN+uQmGKimLW7zuX/v2qezKq
l45KlPxYcXeRtkWmdgCPAZfCdXJySC5VD2s/OZylo3YsP5vjhX6YChRIMi9BB1Ez
dg/7xUbzHytgjyr3Qpls1BgZfrG4lyujqcPtdsdRAq7UlxzNhPUSlqR5He4GRpif
azygD/fAX5Y2Mr46yK9IeHCF3+56KXQsAVmb6vSVms9vxhc1iglyTQdYK650mECW
8WHMW09SH6qdhC8RFUjLm9zWL9uqn+vEndU+5o8G22Zv4yor6XHB0UIKR2runR0E
1q8JdPjQ0G5sQ89v7uXjFdlLe3OLr1rRzzAqLQ1K5qPh+e8yzv0ePEzJGTh10tZb
V4WJMCiYjahP4JTrsItsLymPgE4fRnalgCVlbKzgs1Hcap5/pXJBZ4cK8yJguQv8
Gov2Lcu/uJqx0VPVCj0qwZzN2P0bQk0TSgQcxZuyl70ez5+Pjzj+j/d8BLvDXvVe
ljkpOYP7FTIYKGGWArpWS901Iv+EruDujjUiZ/2S+aaoUYgOX/3N8/V5iMyPuIEY
ocSXC/Ty1AKvoItO4zmQsDyfQYj/4bpGUR0luIFqko38fppCdldyTH6XFnFw7x+q
RvwFBeCwPR+xfsPoGPyXIuwIxo+H4KVPvtQaNh7bSAzxhz/S+mwL9yAZ0AXrNE7E
CEFnlRQvI1H0ndd5JIuhKu4g2KUuMbIyzGbPeWuyCrbjdn0q9ELFCLNCNCPYBeZK
UGxKLxaoRP4SmPb4o66UM8ks32TH1mE3p5lVWeF/GpHlhlMgFRR7iuwze8Y2lDeC
av5H5PXWhS8KMvuBLcDWxc5HjCoGex45OzOXoVZri1wNkq6SYd+uaY7cyiebw4N0
BC5pdAxAtoHTo104iRNmNQjZEulGaNQrOiKSmrymK39AtVyIAmIcoSeKwtwX/BbG
mjtC5KzGU1Zz62SijaqouE6ifSKl0bKAIpKlw3yHa1pXSQyEbP2+byQVnNpqqxzr
mAM5Y5GDk04ZJxCoxC5pmoxtTz/g+LvaatI0Uuj4fK1WO9ueOgNFHeMr2R0MGoi1
BuERw5S0aN/TDcdqa6Ju1F7EozvRk4Rb/quu0vivUbqHDAl4OIfQharGaE8s9q76
/haG1JhWcfSAapc+ghOcEmmJC02ha/nN1GgixvY65fvscjnVsGb8prNz+19w+WF9
qh6X6+USKnZYL3tiw8zq/B2lipkO3EqHoIL4PJgHtopSeIux560JZrij3ihxsyPo
2nvSlW/nfMI9Jejr2xNFO3pwtKC4HF1YGIOqLVjtKgQVQv6WFQsRmHOk9ws3CsdA
96ysNJOnpiOPsKhAzwnBLVdCpKIukMRT0YpmPEaSSKxk29AkglYW+QgDWv66BT4I
rV4005RVCHhb3DGW3RY8/8h9Z0zmWI9KhSOro5sins+zQhoEtCEP1cvCfxAeYbk1
idEpQDNjS3hAELMFiWCW0JIa5oq0hrZqa6eqNxrH/WtHSf5wfwqP/hj9uCSZK5kM
CF9P0+WwVu7lHqImj00XZ6YTn9gkFMUmB5yzwFGflV7/7/7XqVXYkHcStZqrAhes
evmiuUop5DYRT2dvRQnT2ka3qKVLuKavGI1RHt1aSoy6P3j80/4mQufy2xnsyE8a
dH/ifj7vLb9Gmm3Bz/wv2utCWld56hZZpIv+JjcBso2ifcnqY/mHvWOl49WKXDNv
Mzgd4yLlY0p7dAtay44sS+GjEKRlse2kQF6tuOvFCmUnIhioupwWebktzdl5KphZ
K5B17Fphpucyxl39uDUqOgd1jaceCcxaCOzuUzF8IHYMb8PWEa+FpvBWunY8+FCL
VuL0UlDm/1qiA0VSarKZqTZphUnAnA+KUT9bBFPm/lRXIzg0S0I02LSfDnp3ucqA
WQMscukmnlDINqnXHO5Li+4Z/R+qhxDTspMLTVVGDgMJSwtYzHFCRRdJrEo9glLp
GfRVyE0sve5gOROS3fFPHQmRlJqwjbIRTnb2U4ca3bZ7aQsX7PGeBUvCF/bWUpY4
Kc7JtCIBbhqJo3002YHyLs9PyY4cJnL6za3hhwbHCfpaRya/d13XiAzVlRhnODmc
EaS8e5Vt7itmfSFRMDdVcLywhO5W/8JD0UTTEruxuMXz56YdqxdhwEm4CTxQprqr
PGAgu2LMBSp+t/ZNhF2xsjV4cZPUuF4ghm2v5loQm7rJnwwFZ4KrIH4DEKTlnjsn
Ev6Kwbz80O53MFPt4gfHgucxD2AUZ5A709KEp0xjAgOqG0J40WBCDGxsHVbZmj6k
rRaeP/F5t5th8yLD/uzMd8fS/NyYCA8ZOcGks/uFoN1UTY5IGlRgV5I8TAX7pMSZ
U+PolN67hVHGqg1Zo0OuEaQCAfYjWDDCQuBiOfefG0L2vlvbv4DFFCWNZcCgLwS2
Rl6j/KMM2RRZIQAH4OtG4qF/IyxJ9Q+ElWHQKSGeOWNXa2Of6EWIByFH8sNMmfjk
Nne3EwxdUA2+M90qAaQWH43WKRfLwEULJUIoajD1ilWFrSKCvdWnOKxu+HKYLTqf
2x5lGhMrcEqeRloR4K0sepVPGaKIY3f2uejfTQUE0SI+M0S351v6Pwkpb/OCFzFm
5YiXZYdGVVQsypAWWG8u2A/6eo6ukCa2t7NaxjpBI26okRkLpc9KF9var/6Oh06a
jEGnsY8ni6zIVgaqm2XJ/9LwxBtabfWr1a6mo9CKmD4TEJ6AdlUIP7Tvs+y1Q9jW
VuGvzhhDWNqduwP+4dL+Wx8onI4/zTrvfGDtOeqbmV70UnOZJmNrc/u+A1geArZ+
1ZVBJreE88NaZfYzM/m1jHN1MnBtSgQXz+OjGxdQ57p0yqDjCX3TdRMXaCU0dtwE
pIlVR+mfZcFrG0p3Za3eYrhLDagEtnWNANKQi98LKw3h0f4B6XMW3jAEUDue2OMb
jLPRxCTxNrOj3rWc2Dh1HPTLAwneqNEWfrxBCfU7Hg9TnJ34Eiek36xkjpUaX4pE
t9M+TaoSKX38ubfQq278U+MZGsuvZsae8NALM+7BWfISxi8rmVkoQvhEXzS6MhhP
BW84GCreSVNxBcz86gJg5EJf5cIs4kr4KfXY/T4J2NxXCtcTEALIv3avGEnFHk/0
clB5CGxTh57WjpWnYJZucvK2HYzImEI75entsc+hccGIQUkvi/QoVmUDElm/iQEs
bU0jS4M9aQvaS5lTCCSJxksIC8+d7HF+XF9TzAqe8gPtYwW4X8CC6w9+HdpjfsWx
Y+kkibDKgemaZqf0YNYH+Kex2Lfxyuzp6vnmrrxGio//OLswSCItNEU5ESscc8jU
qZIaEN6ePDjFA19vgXfLViwrZ/HUqVjY82dsJOA7DGp+DztSv9tXvZSEc329x1yG
h0Q20nDQWfZm7M1r5SunUzPcQtHFJlpbNt/Y2G8BWwuF9pW4r/Vmb0GaybB3Cfsm
QFj9YR364eAETF/YLqNsqd09rf9Sj+6aALdLpGsK+cupNKkMzo7c7ogXWS5h0e92
9vwVHiP2XJfcqb1dSPAIJcZMcsnqoZdR9g4pqW/Ec4du0YDdulIpPlZCWmMjxbbv
RB58z66sCB5Jha1QAsO7PLU2W9v7G5HI47RR9nQkBjUSqr64IBRRPeJYHrW0iLIK
q+UqsIL+/p+SkWIN4KIzheuQmTL/1gngFvNvQDEaeIDfbJV5SQldklNM+DEXScEO
0uR25P8WmSR9lM+j7qCNzIewW5IUKB2NyFhD1Ht08vHnspN/SNmFY8mw+L2jZlNV
z6pyva/LrD4kWj2aqlqz5fFkP7ZM7cvwNMgSJGIjm4zYKg8YQF2MT0INo7dgV174
AJwhHGaFRCxGbxV26TSjEeY7990oliUGZk0mbADq1DRqZxPxuIOltPtJesFeWHMJ
bcwMmtw0X1omjTld6FdqQB0Fxq66Od60n3yB6WBTSH2s46MW0tusw5ATFkJrIyBd
Fl1PBwB5NpUf6+o7Ztygin2RJu02R9f4fxRs7gk/NYSHvUbBHb5txsFyJmVM+Lu7
6eZUDnfc+4dyhK+nDb2u4d9DIOw4+At9pPcdArHEEOm7RPRCYiM5mxC6HubFjI2T
eLXooPjaKPCuY6j5QBkh0YoNeMOMj1+mbJqHYo/XZFRXzyGbMOJa1CbBmEXanwVo
PeZWKVHoSRyeNYVe3zb7jO0E/gsSl2rr021vWFV8zYtCnNjtnRrX7bFrn5H7PA8+
81UP0RxD+aLccgcpA4ZliCC2qBkQsSl4ADuNSc6u2NKaiR2+u+kEZXaAshY90j2k
TBxqEy/TAss7z0Eg9Issw8eWw7GUWfiq35k/qIe6jytfA78bvMPlAPvlsTNkOsUC
Bn8eQo1ei/PQ93/5ywHIYCeEBjtB6daY6W4WsCp9krQnnmMoTYXx0MQ9GRvpCuZV
n6wok4FRoq7cwnlo47wAUFtDkHa7ltMbo2uSFUBIMu1/waom1uZ2t6wXHYot0mF8
MWpLwLh/C0Qb1Ru+81tMJVOI6qbnTzFgc/Hh6uHow02zLpBzxAe3GfsxQrVZutr+
eehJht9NxlI7hbPdTYYOP3OVzGaVbmywnhRNmK7KEJaIbnuvf061kiId1j5ixooR
EpxGLJcSRKQXhwrxtqGV29AMefyfSyI3TODg8oAd65xLNkhm2Sc8kkVWVrm7+053
kUIP8Z3qPnWB9rEdV0As5sOIqYsbKB9b8c1x9gCgij8eYwF1AfzSiRxNRq2FewMh
ZpixpcVkviK7jHBq3Burx5m1LIZETpszmlsZDmsABJHrY6p+O+qCiOsDcIjoKsqY
pL1jni6Z1nq5l0v+/Hb5tCk400f01D56BB4nRm4tLC04JAtL7jDt/dqYaKpCXNYA
YYrskNIOk1WtBqyQSGRDBAT0ao7UXNjZ+Gm8ioCGCPTQikkkA2tOqzoLKnPPskh6
oycbzGMzK1G8aefOVSDiIdQlDdX9G78spbKruc2vPRrU6KdE3EJJmAS1gyPn3REk
oAi42fP13pGHhbNye037FgNcK+mGz07pQncCHvPwb3fT1Oqd5wZyBCh3MstMg47N
kE2lusXNpOnrQQnKOGH4hhAFOmEqRNeniIkkBwTH4iU6k0TWuy7hQoJPIZZsnOf9
sI4IdXPNIbxocrzIVbVnqalHfxHNIPKlV7tH/aWsQLNRmPtYFySaH6XeDv+i5Np8
akluaSNzYsJff5lVzIcwoJeNgyn1Boe3LQyrrZKaJPDeHmqVRVuOkC0ccMy+wc9r
UnhoirTGK/h9eD1U57+5HWm9TQD6vFGc1xTzDyADczx+3LngDzZ8onFi4eXtPEOG
WhV7Txktm/Gv6I9cGpYvFixoeDiaZYsW1EmcJAg/ExLu24HnXvTzvOOjYWjgbXkS
MuP73Y7jIy7FZjg3vdQupZ/sFiabI6H8aaiA6/199v9KwEx3en6UnChOPTCqfPb5
lDRH8k2vLNibYCUhRKUZaib16FQNkQGqBkGTAWeB5xrsMctG+umRyvmVo7/LR1BA
CG2ngCiEDxI0unmxkeBXsZBCgNN9pVUI87Lymn9vZmMrHJwmBrUCo/wueluD/fkX
Dm9pvO0dl+DPuHDJVW9fx8FjKDpjrRBautHQnEnlW3OzXW9wazJlT283pkfVytYv
jwRnjUWlXDSzeyOEc3IudGCy5pl9GNifZxOxIzudKPSAP3SjFJPpY32PuKbUBW8A
4D5SQHjGXz8EYQ/r8Q0Sbqx5P2DEZ5saOMwt8MLTovDqS6C8W6v61Fz6W55NgQXt
x6rNp7LAu0A2EPI6O5flEeG7rZ+yOZOGGIGKn6VzbeiwAfRjoxuWfzVWMwXRsmq0
ZjnMZnl0Y87fPM19m/R+6We8LDrOsimtHsxpfkZV9KFMl60WRu6+1KEfgcgZk8ek
qhIqM1vIq3jk4V7dnz4kqNZryn0D7/s9K5H8fsfIw5gzVhbxVLgMfYGC3NTATq9i
KaqFvrMXC1rLvXkrgx/r2PvkBGbn+fcVC1vRWHsdflFz6/FOckXG3FuRn9hopeQ2
GvuHcLR++l+d7qTDglpl4XpoxV9/m5+qJPt3fALffuvN4Hdc4fmwziho0d2OgtVT
LYGQVtT6yfeDehm45l9b88g62ldMLQ4FzJ+rkSxMhYCUr/TjPNn6Ho6T7fPctntv
EUSIBaddeQs4Bs8cpJwtsTzfGXd/jepGrcnQJE/Ms4iy1l1JbCTIOacPUBY96vVn
ZJRkRGgNm02Uicp82CZDXZMTo9dGvfGB8DuCNjoGzVp0pv5H4eUcKGKtew4kHhj3
5WnbpM0581VJZ7CvmE07pQU+mLc8qEcYpNDX2Exv/GODUzE+RNWIeKG2dtt4FkuS
5DcehwxY5wvCoCYUF0TPHzE3LjMMr7yFXR2TuPX+xpUYVQRaPaqYGLrD5IaVC3jF
`pragma protect end_protected
