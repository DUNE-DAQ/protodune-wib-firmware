// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1gcre7JrHc+Y8vOJUMep0TDEgYMrUQlsv3CRT9mmdQ+I+tgsB8PpVX+4stJ4XQGVZuKKGu2YPNmc
TGCDF+kyyYqt4o9gYnYW4vGAI1uxtNl1G+h/YnFjjVUk7tN8LdEfN/P9pEg4Pr5ue9/Md47BRHA4
/GI2Qm4GLpXpfPUYMyOx4V0d5cC3ADqXYNiEGnvjloCqT5O7If6vq7VHDU8r0USIWlguUoidXRcW
yjGguMdDIqynRozaFf2cYoCfKw4QBkKBxdCGZR+lbT0qGWU4Nv7n5Q4Lc7pBX56Qmtkg2xeSd1Su
q1kTSZU+cItFfWT3OgPUGTXXLW1x3pruaA7G5A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10688)
1BPaAZYBPzwqkvbTLwQkFMaGjwQp0XFPxsEYP9zohH8/9OwxBv7BL6jZ/ijXSGtr3fnCoqkdEDqi
LdzlWayEjEWulmqJFMZygxu9bmnL+B/dcbWrY4Wz2ODWuGS0iSZK0zZcxx/dM3ic7cOxVm9QGD3r
wLVZp4+aZJ88adhU54dQNi+6rhxrvARN2oRLhwc6TxoUlU5mi7D0wtT02SQPni6QGRrbfJHtyxs4
pBHJIC0FOkEFiM0rimL7o8XE3nD27pEYVrP0gBf3US6KgEQ8kRtj40ksS3PwYLLXj9nkg5GW+jTR
+aRl6zyo/L91xiPurNmgxC86r9PfN0pzoqXXCxRDs7dvYjMO0kZtDipyY8bAjgKYKR66zekb1PTk
NeJPNQATQCh3O2mPPCv/zDqaRzzilMpeBvaBAww+oIYxUY4VA4ILvDxGCbhAlbfc5t/9xpgw/bd/
dq0JLArOAuZXDlLjsSRbMgeL32pSmRu3DDgm3QP5s0opZpzZzxOcry+ZJxUgW5IMUz70veP6V7ZT
aDMnCpAOP98E3FsODThlje81EUHOMLZ1u+Ucqp+/8OIAwpJO2/Qp4Mtq4NUBaoWEDpxPPDnOj/vs
y0pMw5ZBOMzOZGeftOnl5RFIYXmjg+BLKC1wJPGl6wk+Gld8eXiASypksf50O3QV3useiaZrtSNO
R0mTnS1/nPM1KKcIpq0xxGuCb5/u+4gghaSmlXx1vpXwTzj7+SWeOp2TTiXcbSvRH+iFJTFI5eWB
dB3KigM/6djEDQiWr2B/me5QFZG9fHWNW1YyJLO86JIz8wwYLHExLOuXQU86GlnWw7BrBtTJXY42
aHRj4x9Pr6ZaSTw2yTor8dCJD8Zza7+vLZkByU3hggmeNxncSavmITYs9MzyDfZqCV76C0sjba+D
dDeCaR3kjLZ2L2B5UtSzBMKxRmOin/1yKWgyy+XvQ6QDSi1tGzjC/oQ+ZM9/tS/3DBQUW3jt5WPa
vxrwnVIRZWV3vdvVaiMtjbEpN1/81/QHYBA90WF1cqllvn47bnRJ/SbZfTVoEtavIGqH+5i29IJL
L/y32LyYzrrYPRLXhCQh/p2+dCTfmL2o5CJpmFP4tyKpzZrp1TEtjjd4F5Ujim8bVJAjSw5hoY+y
TsQGBSP87+g2nZSwsy3sU9QeqNBJAH1MzYnporgdsBF15zB8SeSi1KrzU1QVFcLu/7T22TXf3RlG
9VaZiiKl1v02RNXjIzT4mH5oEA01H6/B+X7uOa+w4A40DprN2gkgTiyfa+F02OjZU3lXwT5zoNx6
7vbFaE/Fyn8hOt7iHHI3ymLWBYH3igo6g3ENJ+wR+hVrLSGo/OpbvPBNmLH2u17yyOib2miimVeM
ln2NQqDC7oo4fnOsuURFYiYW8yhTSnQMI3vs19Nirg9tqNXWk8f3o+zxOUFMi3o8toHolWqcRmQK
7sbFrSRd7kYRX2ClnQya8EU1rj3cWhfNTcvqs2P7ofEi+qP+ErlweGUW7csbi4SLhFMOyJCWAzyh
zoch6b0a22x7R+uX1RtX9an34LkP2dkXVpZHQ0jJXxW41IdXF+QRrLOy9T0DCM1jzecY08FRpz9A
g9ak8EpXXoJpqao6Si3TlUvMRExzipWT+9rhP1geLN9V2+Sh85BhdiaEt6wZJGwgFA4k9144ZxJ/
tJ5KXjg2lTiLAUN1vaG3FVZTplhLFSfyhj6kztv83XABEOxh0HVrXu9g0Prp5Eh4DmeaV7/HcbzX
j0Tg5Qa6JLN10PAZUCow9pb+NDLW+LPNutGlt+S8FW3bCNlc+m2MqIAWvLCYpfXBZRtI4TsjFDNk
HpXTh5TzGDQnJORhXBW82f4E7qfz5/VM+7zPiiTwoGzCHBLipfzREwuyu6qd4B2wkkHQX7OpILTS
Rv8Bc9730Zbs+zphbb2TgohahuuWbYmmmZSD8eLexOMmmuoeGCqg9rJSU0XCNU/A4zUhbzP1SVv5
XTmHYO02uMIJAIgqg6PoHwibn1hvvWrBlqcQn1d/J8UXrM1qf1+q/jbHQureVRmxFUCCUf4gm4fl
fiQj9h43eWvODJJ0BKqYLROmBu70NaCuuZleYd7+Y2FOo6LvvyainqlMUyn4cCCaFgdfE71qb3F3
VFHbIDWdgdxcsRyNpHxIiw5gEWqQ3FlG83iBNBXPvi1su5LIl9fzDht5UzPsFOXKH9TdnOFTl7Z+
h1XWT/qJyUy42DUzcY7mkKj6sLppXT1vKPqlTt4EMPPnj5Ux70svuwj6avezUZBu4zVklL6nCrYV
wkc5MNYXLci7g/Zift6ZJWkAqb6CKfQ1m+3IaDmuUyJmK5Rin58p5pOzCQey9Dl6j42uhOnHaw/W
zHf5XcHCsYvdfBVg/xXkiIdwPDECEOgNedFs92CN4jFaiRT65NUgPGSdfsJVeGZo/abu0uzDZEnk
0ycg5HQEyvdngAjMdw18eXhDEPx4EOFTa1RRXMe0cn15nqxjynD5PrSwGp0irS7uKtQNaeGnZgPB
oqa0tYUBmv+JLXt4ZIJa0sGbdoi7HD+USmH0b9eFNVyEBke4XD8w6rsu7M/huQ+kPGOzOOiRkY2R
UqHAn1yAE+iyW7VXeMoW0Eh7/TdedtvEVXGixehCD+ra1nBiAdG1HcKT68+f73qVWXLRtt4Ojb+p
/f2LhirBvnfCtcQxxkkNjBJCQV/XB8f54Q3uCWFQ7aOMFBXZ3oTw38Luxs3dBiGjsF0sePoCO4ch
am+b4qNThEv7zDCalKFRK4panImATeoYAYW97bFvutyUBXWlY31ORzyRRXah5NCBvZHSa4ycS1dL
EMmxe4ZorVlqo8Gajm3xZ3zZxTFkdYRTOVSgP6Bq9T7gRtTtZsTSOwZM1KhA7w4J506QrFsjKNpv
M1+/v1zMuBr6zAwz8m31TLQZbaCivLMtqR+E+AOmAB8qAIxq9CtoFkc+VooQvVlqs+Ln93/gfwU0
pe3dVnvqhRNAXyNsxWsrNCXGmvZVrH2cfWU1C3Yi3O/G8zTrg8WZhoNF5UGt6REcs6R8duT1m/Y7
cadX3wCmku71YYyY9htgNLeI3C2TmsxCadrT+2gxBDxzREuMdEpRi5QQZbwSS8+GnIacMF4/zgL2
4ScZa9rdLL0t1c7/fZRj4cLZUFTwfC7qmRDINfNxKZRvNKRzy368Qyd6+ptThnQ8ScaNgh0q38rR
vlXHIHv5i4ohFCcrEruvdsXEKjJWiXT2d7WMts2xZMkvQ/4cK8T+HbZ1BqfBOuJpMCVdNJSWFvz1
gd77dQc9xUxN0FTjDu5v9gqRbz/Icb4Hpz38mV1yuP8BZ57n0Lpca8dPrOn42Afy8qEgyxFww9V9
ZaS1vPKQiisaMgmMWEy5NsdII8Ayk6rh+jhjVVVosphc/RbE4V6jbJCTngWLPmBQ15fgIAYLxEP0
EQHZwYH3t8oVOjWK0UBBv/zBgEiyddJTOptFnDXj+bHh31fZX9C4ty21iahGo0vMDj89+KYecYph
M+317d/FC5bnS1bIDE9JhFulcPDXYHO2maFrKlxKs4mE3bEg1TZZzDd+QWA/BvB3JnaetPY28kOC
RFuGDHCxtuD+1wajnlbF7NP+kYXD56CQNDbuI4Eq8X3+7CN1XnZS55HiDC4zc9QmwR5vFR2MLXPS
udIPk3kC5OFhRoiKJlxQd7K8Zr9A/9Y+mEg8RAGeNQECcObnyC4ti6kW8b824YJLOHtXvR44kf9M
em5cWXQz7kV50zpw6JMIUJ7ifsFPr6aNNHICICTZOPW2uQ0W0g4o667p4RNWgZ8kTCQEeV1Xmzk+
7CXRbAFezyJssTGxXo2xBlrjN4c8wiaeozgM8P2FZEHAAo22PbN4IXmyJvdeK5UIIZsAbkpScVFp
rWtZlTmKOR910EuSvE/Tz6xePjU1aqxG4gpo1M2gTPUsxqsttOeBZSWIEOzHyvYMn22hpHVvkFGw
O89cDtHiY1bG9chDRdPk5KQaK2g49qkvs9zISzkTjcZGkxyuvyajSHIxfX0NBB+08A08WJqCxIjp
kFDpEM8jX3yyNN7xKowz8RC3MPggT597LGcmfvGsJH4RqADfUo0iJ7nPngtVEWanuVJtXxpPS/sV
i4fv5UOyDTvRvpyvlBAIJk5VWUW2UiHgNVHqUNPc5sY0tyOncGLUrKofewewUUhcB5hWthhGBZo5
PoThqJTZA5YSz68we2WGDK6/BotqdJy8DaAlx2NAtOXTiYnXqAB6+2zyFP29ClbVG723/dRQwiME
6onHHFMFflXzpZs4PIORvg1dNSe20cPK9Knm8n2JrAhHUupHtYKC+l/z07E/sML23ztS/nhKEN3C
TY6gklRMbU02m9l1Io/GgQlz3Y+yNXPyQvR5zcFPH5geYzKVDDp1GBsVeoxRM45pIMyv0cXyzqLb
R/oJsCUSzoqV5HzbOsRAsPI2fL27E8CjiSyZnJREGHR3MbQF2Xf5yOmmSAD3YrYHSINfyL0hToHN
kRf7UBZDKuK4PbSqjcJI3Nh96+bdnuyxjhfQEiHpsbMGP+0FTPxPLP6mOa7rngCsEm0qZA15YNpD
kWWa7Q0P1plBoj5T2Lk07OP1ysi/AjPvAstxhA103HPfb37I1dF/SAKOEKf2s9aHFYPNGVNd11re
LNS+3dFx/99cmXpn6fqeP5kGzwzqdSpNQ7TSjrVPcYxxL8rQwZGL7uU0DHKXMCStDhUME1m532ff
znkQMODshTj5A1CFVwRJ8t/q1ybKSn/V5Pn6L3fT1mLCa78Cf/TYQvJmI1CkrqS8MzFqQEJusCjE
EpX1sg9D+XuyxEP3EG8R6X12CRPGTRoYCeHL66s3UyS0/K5aQOv1x7xa+lo6UomPTErjPAN7PcTx
e/nUdTpfAEztXN//WwECGwgoMrkvAbKrOmfR1rciSWYooMx7Qa2fJcRmF/Z5+BPw8fVzgrLKkmRy
y8Rflfdbzr23rRwjSSVKbj78QIksek00CfOjiGBinSLCMvqlc0aZ52/kYvl+7iV7cKl2UTZJYpKk
UQoTZH6x8w5d5NNseEBj5i8sI+L6ELX4kA/LRFystkVb5s3pU945VWMhmCPBQ5arU4EQFpLgWLxx
vO+naRLhM09B18VTafMkHUyUWf6r+2RTcJBNhabREIUjiHbOwwTI0U1C6m74RdedXc6OjCHBIc6T
CisjNLXwhb19PLXm/YdjbkoCXo409HeaCIA7I/wcW074aBvVKCYGGgYfXqClh5ENcBk2+xtbt4xT
dFPVIJ//sy5viq9b/ZFU1PRC7Z6H1klOPARneFu/w761FNgsx44YXGd/XDRvOREBroiPmey31iFr
9pTKPW+9CV18Xu1xpP3dUf26zkL0/7oUAnOkfCkBtddCdRkFfcVmKGrP6/09bKkRnfWlM4UHUiPP
uUpgP9I4UmXA3vjwUBLsyvx1qs0GqSj4Zo9ha+gEiyIzAVRtrsJTsWppGHvoZFPYnq5Wmsp+2QKk
IjhFFmCXCIbSzzePtFAYCVPul8PmCe1kbLmOMPBsv00NMkUTQqY7TI0ruMKkD++mib300taozX90
CWPZ115zRyEj6aQ1JxogItREgWRzvGZ97/B8T/YK8t6DIHjQedrhwaWJuclrt5+Fpd6R5ivlDIan
nBs4GqZGBHEuFF9FcunW/zlxznIWtxI1+EOhhAj6JwA6UFHw6X+6YY1GfbmmKkN2Q6vlGTkovfHz
ZFKxqIOOlbtuDWTsbj9Nykg6ymQWM5CdqtSid9WHO7XNj6ydzwNQToNd6hB/Tz8GQJfdFlz9SmHW
pCI7N0V+OxUOVeqcUC2c2ChkIAe9mvnfaObaCDJerDvBKt/xiH+bjivxUd3kF2CZX/88VZmmONkL
Ol3QUS5Gy41nPI96XLMewkaknPmdfxAOefEIhyk/V/BPB6oltB/AJ9PkJ4JmymOhK/RUky3SsMo+
UsVP+YJtpWJno+QcZAQt/eOg2iCqdeTEapJrAtbyulUmim+wsXCDhLK6cCFzKpPcF3L8Un2Vnmgy
y2KQ2p6YLIuAPSKiQ6uEsW+p04kHs4u9KFvuhNdtgKHBbuPE0iYw+Q9rI2lyZV+T+ZN9KsA9x+kJ
LbITXAE40JWFLMxFIrSTXAi3/og1Lrcw4orr+/eKCIqsXDGUTHCnefawHuTGbNntkrIjM607Dmoo
oanAQc/IEu7/k9rW6RTmMAr1G2QMnQFvhSnKjNFJZ/F4xyjQM0Iq1s/XDQjcylesQPQJJjcEQmCV
Kg97v2CgxPOPXd1LxecVt9tkvxspVKeVeJ4u3PGxyJ/EjOF+xgdOh/CAO1pcxfSxB0v4eowG5xTe
mPjoNXVT3MTUVH5pfrS+hk8WqVy+VgA9VoTJ1ycLHAMYq4EdNfu+fkGZvtICXVm7cMxId+S5DGxV
reF6Wm4bnfPuvBRDJF3KAgWi8ZUqBb+d6tvShSKe9m68ohIDsA8w5zduiSNLeV69+EOumElM1i3K
SEKM7r7wvUE3s7zyvXYa2vWRNzOUofMTLZujUqNZJdcGb7cRuJov7rb4qUu36L4hHlXHa82+6Phv
C13pdJWjWsOMWrYwgfq3ScH557goQq4KrQBQr1OJ0FpYVLkZkIcszh7J5KO9fMgCTGJ7bKi1Toq3
NOThZFtNsxUH8yU/yZZGZ4y8xG0MxuHfi74BwJ9sfuWOcQBurdslDbpBgM+1oRVqft0Ek8HK5zV3
PrCgbJrVqzTwqMQZ1P/Ek/TOuQu9CCpgQ4SVK1BbqJ2ZipbbzYmlJ5S5cnyNfm1dA+p0XV6CqtLL
izU21yqK39prBdqEmOFuitcR+GgP7rroc6GZEEbf0k3w36nDCvseg4No07c2ens+tfipuo0NxYwN
5jl72GI1mM4aehWwsJURYbB7Xjj7AXfS2acSpeJ0RFEMMbOwmo2g7ajHItIZW+k6vPftS4ZffV4A
PizaZ5Y6ZFEIzyxFJxbvP2GBSrDtED1i+HHHJvjq2KBCw/FUbGlqnJ/BXWmva8EzDerGfTJRJn7/
Qr5vi3zv2tpdPc3ooHSpvYBXORnBSTjJ/qsTjWoa1FnPyL3DVdK2xtI0tmvG1du7BRzJxoe0JxfK
YvmL3ojpvhxjPaPjkKf6p3kof45O0JKc1Ecp7Cg3wK3lt0/EFhBJ7DjfHtZgPNAFX+dXRgt4+ZeT
CB+CQbHAIO5cAzTJbQhubwk6Rs4Cm7GM8mCeE28visHrbxH9eo4jdtW6SuAdbjKO4+Y2hlSeaIjy
0JnitxOiTuEJt/GfP6H2iF5853wsIdew5w8yFNatywrd9G7XMyOnSQcP4uL8d4UQcd1/yRTbwTpv
31LhfLqn2TrEcEes6lC+GNVIS614QuN6UuFyN0Ay6bqOyo/LVQlE0oqq7bG/VrAxS1ytS7ayiQAE
pWl/S0XbIDPTKKGNs5oGFdwbo2r3sM2l2MVmXi1y9RrF7IW1aQaKFsl1movlgKvLsE4fXDDtIVSS
XZ3p6kGvwa1VltWaVstDZKSn03ZgbKq5yawmfhdtNjf2/cwORreV2+GUW6h200o7b3wKrgifApfw
eaI+L8fTq0WEfEQkHqpzFb1eeMmrPeZzld/xhOJONYu152EWl+ny0xMrVHoeEmH97LyErZRPAQuL
Mqm1Skp9ENOBV0TCKLqmb8xOUzG8p4Qxk7ll9swxPVjyguH29nNSBrvR7b/nfyHtaxXt4VQmzeye
VJFuihDbJyuqYuw2/zYx05afm/GRoJiYlHzW3Lj5F5K6DwFWXqezexxGesK/GS63dB67Y0poRgjx
+iMbeqU2JXDGP5tancOZJ329B852O077Uirbuv6Gmsq/Or9XgzyHTX+O9yiXSdZnu71UMdHnNQf+
GFPs3Q1IPBxFyVWBIXkg7vBenB4oNBTSlQTBomHuh+DrlsoeCM8RxveEbCVMoHqPoj8dqdO1MZ5S
KlzMn2F3u62MO8++h1JzDw+ehPcIdKgcO8drBypM+B/bjkMs/HL1yz++TNMJSjBx29Fskaiv39RP
9gu65b2bq/BnzYfGqDgHH51foRKQhrlON3a2gt2DsxsoAl86KbZyBb0xzpOoFb4SeIt5MH63l5qp
zjC0RZfNTmomspOyQufpyXdSSUb112a5iJQmfCQFzEvgi60++B2PTfiCfZbUb4wzbSe1MgO1v+aR
aoeIetEyLHpMPbhjDydaP6N58OKJEnMpZP6vGvl18CSqsiuU2kGQ9XYLp/4kxg6F2MhoQzUDGyZO
niQm1AZAfnr2FgoPmaXcbiZl4BwOrzz6CO8CRabCnKb+ul8Se11RwrFuUVmOW5gtb8UntlSNcQeJ
BxAcScKbfLDN0sHYZ7YaxMFJ1kCdNFDp04n/Cu1lam5xxmlfUXHsRe7pnzliF7N6ksn1KGdYH7cc
s+XL6kx/UGVBFy9fMQF5vqK6zBbshIFliNhVNCZtTLWWo6vmE5+M5Ie+AM2huIV5vQ7Hbzy2+UvK
nCZIPrCnghLkw96FxkyQZ+4AgMu2fN5OKmec6Ox5eywvELxJ2VHIWa2r3KdquOnHPM0iOUnNMhED
q05nqAWQXNCRutU3UYNYWJeUtdvFzBIx6Ynmw8OI7FsyBLHAhcfleOOsR7n9JFtzt0zfFYGnyxnr
ws5lN9l95SiKAJtOTWvODBMu47FvJJroT0bkoLWK8v7LN8clCaKqWK4c+WgMuAIiuaLM4DXjVMKo
3DBKlB9GRZfb74oM2boi/DNtCy5xshv14Ucx+SPluRJr54pCGLB0Mlx6ZUdR5blR83l6YVETwuhp
vRvuGst6j4g+v8blmNat+XWCcCuTWpw/9ddWTgJnsPkMnwWD1/o9k/cmUwjIrEcbELzWX3D0AdWE
ZqJMEHnowf8PIyWblmi6To9ZGRbuF2ad3Hhg9DxFieXGjV60mCp7s3M1+CZNS7YXORc6wR3AHwa+
QIgeLrZOR6Z/HgyA6wjMWt3CQIP0L3WP4eGMcEl/APSEP9wa0xhEWeWrneksofeaiR170cOcfxMj
VFWWviU880j/P8uWz3xIEcN5FM2bGV1Oh8dRBvp2ZkIdP22McwHLkTKrGLOcRaYUfuaanuu1d7EE
7sgqoioEKGgCdz7TCojqR4VQ88Waq3Gvk73IJ2MuEsxGQyCpW9oOTdGW9DTGMW0qL+KZ9cjdZq9+
dSwqM9qCT4Mla6eCbUBMRR+0vxn0nqjuTi3N2zfCBu6jZGcqsj/Zag8Epd0CfjNWCodLbANOLOlk
x6b5BFfya2lFcGJQvDihgAvoN8EgH2U9DHgfGph6gt70ES3D/G1YkCKFaLo+6sXkhq9EAWYk4ZS9
HngnKMbG9+u1JLxBv8T0FJPC+rJsYaBoB1cMCXsLAnPRj+6oTm266p87AWp2STxFOyd4u0+TsD/u
E2+QXDgR/dSr0ddkXHZG0lutX9iV9HxFMWrUxVLRBl4ThBOMWtSYMFFrHqnok1JcYoyVoUkPq3PD
xVk7+S8TcLXbAmH+B+7KB3UWHJilfv7WXB/EoomlufjYMllFgrnXpnggOIpCgi5WLP8I78VOYM/R
VxWcfh509YT7415cK62ahQ3nDGx3ey+kJ1rDvZxhQPWKYZEtyFPQbVkuSzVrnGNPhdGzMVpKNADS
4lkZOhzNbJjTAg5vzWfSFlNBb8Esen/Nkbi+lmvpHKNbS/RGeXksis1geBQL1g2MKQ6eEYgv1owu
exBtQ2MhLuH83MGgAkC5veLGBKPe37hBQKjFeqT04SQHwRZgxytnWo9d/2flTUkgUWdIW4eMFQqz
D14e/U8xT6eIbs36ETFUzROgsIp1CNQv6xat13IsGbkvyXzQ6JFS7Pbh1mIssLEEZWDDa1JSTbsX
30ygkSW2a80770HwjTKXdB87YkKc0TJ18ZnqSFnf3wfvRC2XB0a2w3wdvJRQwDIyyzSig12tkfHh
rI5FlIQZId6PrgLMkKounRLn67mzaUdst1tPLuJ6Y6I+OTe+jNTJ/4o/Ne9eobm7eBO7bjzAkOqn
DAQhDh7lPf+N139Q/TyaY1foRwMwRexzcmz+KX4FBNj8k8KM9/Bgh3ZMpApEpR5AZjngSMF5t0Fc
n34AnkCmnBfiwiY9TQXj3O/HBGBs75T72UB46BJoWk9z1Ldu+3g0QAzoS3LJUgJyy3UkS5tEwC75
tY3TilP0NG7y7pFzAMp9jbf/cnTc0gmyX40NwWGuw+sIT7Ety8+YYZIDg3H4QV4vwVScebewcOkC
T16Pb1cGw2lqE80HB4unbMVdiRdRNsCzI7t59gWBHuRpi6SPJNo7r/hov5feDBFo3rZ81vYNUhaU
6V88IFlFmjXd/+35X9oHPbHgI8OytKUbJRuJD6vU0T0xS5YD1CANGDavA82kgPPDEtpE2k6PH+zz
3aFa2VfXfbPm/SjrGHg52cjyZ6Sacyt9epfop/LohFp2rlCPT81aHbZ9QPnfUH7gG4S2HMG4aMIG
K/rCccXCQJmyXv1MVo3OmS9nuTpknYkaS/XMEEO/TdMkaGBJfX7Muwd59oQYs7wUeRyMkPqzHGtI
DuAbHOFHWgu0CFWbNu38BUombudBieV7B2Hl6BXSRHXA8LvHJqq8k64ZQHQGlETA7JDBHehsvvbs
JcJ78BnTs+0Ld+uxDHDlNDpOSM4TV0bVyfYEG1x/T77N+a3wjtGi5DCfUHqT9KmWmj6zT2WyaVKl
dsoqKszVk2sz5N/J8CJtOyrf/gHl6/+I6jgyC9iTV3RbWupfUIv9Umk5mOyfw+ERj6WqMffk73hf
YHXbfgEWnTyciplh04il45MFuv/LBW+xZUsoEQAWbPtyJGVRW5WNeOzAhHzM5qnsIsBa575OqDtq
CrTlf9oitmD/gCVLGRSCf4G/vCc8rmRu2p93lkxKY+Ua8EVGcW+jvzM/Ap3woCxKud0XY958QUXo
yHhVYdf+A8oRold7y2hhntGW82HNgHlbYC8YgxzHe2SNc4WFO+A9BUgk8qffgXLxnR6vg6cf7+Kx
iF9hz/FstWQhs6ZldTpj1lL+6WOx3I9w5eP5ufBHTgSehf5sdrIEBrVFsag4hdyq5QBWjASzaoQk
GJA8oxh/NlqGO3Xb1WR+5aokJ7z6bMuLORgJUMAOfnoz9f74Wd1MaKKfIVFSx033qRe6FITY/BDQ
Cd8lnsJL78WM27VQy7Xt0phgG7i+nt7OC4bVCbcaBiR2t2bRRDZ4mrEzAAjlZi4VsKAm+Bsh+FiV
4lwz8rtwuUbp/7IaiTqY5zhyjNT6gh6/DOx1Ju1nqWa7tGCu4ufcZJG7cPDFk+sC1itQgO96qlNo
OYI8ETBNGwXbuFiFA5cRLzzAsSHeF3u3KYx9FxibkWukA9yoObp1Nm0i8PGYOX3lnOTOZa4Onu7c
dKG9k/paN7GGpMMGj/sU7nyAFemxIBydEfjTkwQZx+b14FlgtNsGyFCX/pTm2vBPpsOfXzJxqbPj
L2e87WAoA2fUaZhoyTvKdWNgu+iGbB6Uqk1PK6hNlbEEXmHOXCTtvVGg/EoExsU4U5P/7k59dJhV
Ys3ZXraR4Nnh6fR8RLsR8pnkyfactImxlK6an+e+bEgZglJNzE2A5B0uI8hORAQGJIMjN/Gy0af+
Z8ssK+9+7fMapZeeRrm7w/J/67s/HBlDS9cdQCExVss7+CGXaiNqHIuHcrQ6aM1B52xnpvlwgt2b
CfO8kNnXf097EBLg8LbQhF6g9eFMQBPQ7soR1Go9rkT8vV5C4WjJPA/+NForEHhqu7N0gaG6vXsO
PC9Qoj9N1O1bu2pfHhAm8h1kNBkA45BZHiSBFRh2uYzgn74VLZC8W6q9zN7z5UDgr3Fx3jbKGL9Q
I9F4e79TjIkO6Guz5b/LhHuqjjwx8UontDyfyQhCKIay9K4sHIA2NClG0S2A0K3nd2bZcRP56nFC
D05GcK/aH/iRoZP3fyoIcoz9Hqkp6ZZgNFzii8AHweoflE3fP+tMieqF1uMagOQpWLzMDwuV37xq
5mKS7w3NLErYyTbUdh7k2trnV3FeS0bgOjQjg2DwknFMiZKrgNIPUmq5zo8dFIzi7A+072Nve/+1
ZLpr+lA8j1YBFesVYshh9L2ChZ/1wMKh00mIx3u4kY0iTqzi7y8gtUjWB3UOqfQCd/puKyq2VM3v
5Z38eJVkegx5TwTmdSJ/Ffrg4zIGgcziPtLalmajmDs1LGVJxWd9yk5OOl0Gvx1AcUP3ecBhWNsS
uwH0jzjgur78LgWnWaa80iEO9Pq0Pxvx7kZGiorQzIziRkOCAB9ivT+Zi5/ptPaiI3DUVPpgUbEe
3+Ig6GytFHnJQrv2DD+ULX9vU+uK9Lq7ouDIzLZVZx6auMiQeegVtHX3fRYJSD+B1jMshVsPcgRI
Z/LwrGWG+oCpnv2RKx612zfs5OXkedSWAOheq+WSh7YfYPfErSUnLpVBNkjo9wAUIkj7uel4fZRJ
N/qCMCLTJB7xDgTDZ8q+Diwoh+W7c7V0dkViG5UvL/R8wVlMDU+V3VzFFWJiKNCsQJ63+bJHfeWZ
/Nz2NWp43kDALABvv+JcDY3DH4ebZPoIqiLPq5LsWXLVROOMgSTeic5Y4YDGsA6aOZOGHm8/UoF7
owLimwr2W5GtPF+SjL7wD8W3dYoH3a2ne6A79RPg9MxZK9BnU2ZD4HP0yVuahShrU38TtpSB4EFU
gz3DDQwu5HvDIzjOmmD7rCCflcU3yyLspbNzFRipmeHGB5xSvaooH+XEi0cjBh9/DqA3rhw+XTkS
ZnlUh1bU4zCi1D1eGEEz6+VE+/gYh6eqQr04E1+n8/RdyJUJQ+uYZBbSgcptYmUMvimGQGhSi+Un
Ywws0em8GW5kRpH5MmFG83wSaV7M6CrRaI3IiXEoLS9VxJdosjSnNZbowTwHOUMHr00HaF+rcVPJ
mkjDuiHSmtq6AzMHS0UXQ2k+x9aVRpuGpjep8KMbNnIhD0Eco31oohNibh0Gz3MbFX9KLyMwVCkP
dR3PAJaAOjCYJifnTAJPJO0NPm0lJugBd/C7BRZlDETQMNwQgGwyKnfjts7wettXH9SU4BSc7hNx
TWyDRFqn381lBCuYcZ7KWAFRCkgHtjgUQYd8pkodYKJzjOAk2JSanPRndBzGB6tEN0/PR+261EMY
gwbow399tZCx1cfRV3jlZIoumt/iFZFplwMnH8woJLirylIYWOBCniZ/Bifq95weI5zKK1Bjy9O5
D+2WuOrm09vZD2TWAjRM7BEK6ylfswdeG/2LM+s3S1yyohQvXOgt0vbe/qjOZUzao3tkdNDB+RIN
FdBcnt3EVbz9+jFNYaRWhanveCy06OOHIO7thZupuU87zWorylFsm+bwU3EE0eotLB2DkI7LBQv1
SFhtLhDa+P4Ge0FPCGbTMhKAGjmaV7sFLuhAbWzOCLDto9Z8XSzryUvadg6MgTjaW5t0igYFrYyr
nKExZRf1LDffToZr692ijS67oIkg7Zbfg4zzGkluRp941JtUmdZvowqoOT/Ft6Bb78P2O3EDvyB1
RIQMby3cswLrh/R4IPXODc/++HldjPneD50dUOI7VKidFSnUfP+e4NXHbQbSxW4ZQEJzm0uYC/Fy
hSQYo2FV9bfbta/GTLXxcN4l1dblcJHyi9cyCRLK5XgVdtT1AgvwtdN7YofT+5NiB3SEk/I+lPJe
0tT8pJxLHrikH9nKUwDoMZ8X06j0zlbW418ZoT8fbYRXr3Ys8sZLuhjXqq7Zt49OqNRlilj4Tf7B
Lb6TjWWGBjReS2RrLFHe+DJRoSRzwTaV+pfHFI2LvJNpPCfT6moDH2gMFrWDZav9pBqI3d2rbVjt
uKBzcSZt6r7bIJjMM5hSyWKn6rxYsnf71zRLZemTUEKbIv4BDN7iQFfau6Ln6mhFimiQHs4zD6oX
yvKHWWSh+GC9oEgcGF7A9Q/dNTriFx6s65goCnIRic1k6mysJEFaUmOVlKPWyOCVAamxERZHg9DG
wzXHCEDNKX8/1tZKzGXQVo2yOybZ9V0BM3ZCDpZ+j7Sywrx+oaJroMIA9PjdU5UY/PaX4wvixx5l
OcLZY0lDeQgKpcbmrhZliu0zuy76/lKz6Myo427cc7xy2g4XVP5OTEo7Km8YDanx+w6JMBkG0M+D
kavCiQEhyn7DiEpiAFX1uk0rLr5ECtM1ycdKZGGZyEYQMAn5LJ7ir6Bz/yFztjCBlZMafFcH85UH
xuaXpI/edu+rOuW6cOC1l0oI6enUFzCC6EytOMuDh6VzvVSloGEtnC6b+gOJn9nl3I+VzmK+7xoA
XquKQxJ+BsCxf0VOf/JgUKY0CRco1s/zQA1jGUg=
`pragma protect end_protected
