-- megafunction wizard: %Arria V Transceiver Native PHY v16.0%
-- GENERATION: XML
-- COLDATA_RX.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity COLDATA_RX is
	port (
		rx_analogreset          : in  std_logic_vector(3 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(3 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(3 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_is_lockedtoref       : out std_logic_vector(3 downto 0);                      --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_is_lockedtodata      : out std_logic_vector(3 downto 0);                      --      rx_is_lockedtodata.rx_is_lockedtodata
		rx_std_coreclkin        : in  std_logic_vector(3 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		rx_std_clkout           : out std_logic_vector(3 downto 0);                      --           rx_std_clkout.rx_std_clkout
		rx_cal_busy             : out std_logic_vector(3 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(279 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(183 downto 0);                    --      reconfig_from_xcvr.reconfig_from_xcvr
		rx_parallel_data        : out std_logic_vector(31 downto 0);                     --        rx_parallel_data.rx_parallel_data
		rx_datak                : out std_logic_vector(3 downto 0);                      --                rx_datak.rx_datak
		rx_errdetect            : out std_logic_vector(3 downto 0);                      --            rx_errdetect.rx_errdetect
		rx_disperr              : out std_logic_vector(3 downto 0);                      --              rx_disperr.rx_disperr
		rx_runningdisp          : out std_logic_vector(3 downto 0);                      --          rx_runningdisp.rx_runningdisp
		rx_patterndetect        : out std_logic_vector(3 downto 0);                      --        rx_patterndetect.rx_patterndetect
		rx_syncstatus           : out std_logic_vector(3 downto 0);                      --           rx_syncstatus.rx_syncstatus
		unused_rx_parallel_data : out std_logic_vector(199 downto 0)                     -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity COLDATA_RX;

architecture rtl of COLDATA_RX is
	component altera_xcvr_native_av is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 0;
			data_path_select                : string  := "pma_direct";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 80;
			tx_pma_clk_div                  : integer := 1;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pma_bonding_mode                : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0
		);
		port (
			rx_analogreset            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_is_lockedtoref         : out std_logic_vector(3 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(3 downto 0);                      -- rx_is_lockedtodata
			rx_std_coreclkin          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			rx_std_clkout             : out std_logic_vector(3 downto 0);                      -- rx_std_clkout
			rx_cal_busy               : out std_logic_vector(3 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(279 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(183 downto 0);                    -- reconfig_from_xcvr
			rx_parallel_data          : out std_logic_vector(255 downto 0);                    -- unused_rx_parallel_data
			pll_powerdown             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_pma_clkout             : out std_logic_vector(3 downto 0);                      -- tx_pma_clkout
			tx_serial_data            : out std_logic_vector(3 downto 0);                      -- tx_serial_data
			tx_pma_parallel_data      : in  std_logic_vector(319 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			pll_locked                : out std_logic_vector(3 downto 0);                      -- pll_locked
			ext_pll_clk               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_pma_clkout             : out std_logic_vector(3 downto 0);                      -- rx_pma_clkout
			rx_pma_parallel_data      : out std_logic_vector(319 downto 0);                    -- rx_pma_parallel_data
			rx_clkslip                : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_clklow                 : out std_logic_vector(3 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(3 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_seriallpbken           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_seriallpbken
			rx_signaldetect           : out std_logic_vector(3 downto 0);                      -- rx_signaldetect
			tx_parallel_data          : in  std_logic_vector(175 downto 0) := (others => 'X'); -- tx_parallel_data
			tx_std_coreclkin          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(3 downto 0);                      -- tx_std_clkout
			rx_std_prbs_done          : out std_logic_vector(3 downto 0);                      -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(3 downto 0);                      -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(3 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(3 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(3 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(3 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(3 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(3 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(3 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(19 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(19 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(3 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_polinv             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_std_elecidle           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(3 downto 0);                      -- rx_std_signaldetect
			tx_cal_busy               : out std_logic_vector(3 downto 0)                       -- tx_cal_busy
		);
	end component altera_xcvr_native_av;

	signal coldata_rx_inst_rx_parallel_data : std_logic_vector(255 downto 0); -- port fragment

begin

	coldata_rx_inst : component altera_xcvr_native_av
		generic map (
			tx_enable                       => 0,
			rx_enable                       => 1,
			enable_std                      => 1,
			data_path_select                => "standard",
			channels                        => 4,
			bonded_mode                     => "non_bonded",
			data_rate                       => "1280 Mbps",
			pma_width                       => 10,
			tx_pma_clk_div                  => 1,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 0,
			pll_data_rate                   => "1280 Mbps",
			pll_type                        => "CMU",
			pma_bonding_mode                => "x1",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "unused",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "128.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 0,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 10,
			std_low_latency_bypass_enable   => 0,
			std_tx_pcfifo_mode              => "low_latency",
			std_rx_pcfifo_mode              => "low_latency",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 9,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 0,
			std_rx_byte_deser_enable        => 0,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 1,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "27c",
			std_rx_rmfifo_pattern_n         => "27c",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "sync_sm",
			std_rx_word_aligner_pattern_len => 10,
			std_rx_word_aligner_pattern     => "27c",
			std_rx_word_aligner_rknumber    => 5,
			std_rx_word_aligner_renumber    => 5,
			std_rx_word_aligner_rgnumber    => 5,
			std_rx_run_length_val           => 10,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 0,
			std_rx_polinv_enable            => 0
		)
		port map (
			rx_analogreset            => rx_analogreset,                                                                                                                                                                                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset           => rx_digitalreset,                                                                                                                                                                                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk             => rx_cdr_refclk,                                                                                                                                                                                                                                                                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data            => rx_serial_data,                                                                                                                                                                                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_is_lockedtoref         => rx_is_lockedtoref,                                                                                                                                                                                                                                                                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata        => rx_is_lockedtodata,                                                                                                                                                                                                                                                                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			rx_std_coreclkin          => rx_std_coreclkin,                                                                                                                                                                                                                                                                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			rx_std_clkout             => rx_std_clkout,                                                                                                                                                                                                                                                                                                                      --      rx_std_clkout.rx_std_clkout
			rx_cal_busy               => rx_cal_busy,                                                                                                                                                                                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr          => reconfig_to_xcvr,                                                                                                                                                                                                                                                                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr        => reconfig_from_xcvr,                                                                                                                                                                                                                                                                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			rx_parallel_data(0)       => coldata_rx_inst_rx_parallel_data(0),                                                                                                                                                                                                                                                                                                --   rx_parallel_data.rx_parallel_data
			rx_parallel_data(1)       => coldata_rx_inst_rx_parallel_data(1),                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(2)       => coldata_rx_inst_rx_parallel_data(2),                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(3)       => coldata_rx_inst_rx_parallel_data(3),                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(4)       => coldata_rx_inst_rx_parallel_data(4),                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(5)       => coldata_rx_inst_rx_parallel_data(5),                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(6)       => coldata_rx_inst_rx_parallel_data(6),                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(7)       => coldata_rx_inst_rx_parallel_data(7),                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(8)       => coldata_rx_inst_rx_parallel_data(8),                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(9)       => coldata_rx_inst_rx_parallel_data(9),                                                                                                                                                                                                                                                                                                --                   .rx_parallel_data
			rx_parallel_data(10)      => coldata_rx_inst_rx_parallel_data(10),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(11)      => coldata_rx_inst_rx_parallel_data(11),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(12)      => coldata_rx_inst_rx_parallel_data(12),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(13)      => coldata_rx_inst_rx_parallel_data(13),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(14)      => coldata_rx_inst_rx_parallel_data(14),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(15)      => coldata_rx_inst_rx_parallel_data(15),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(16)      => coldata_rx_inst_rx_parallel_data(16),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(17)      => coldata_rx_inst_rx_parallel_data(17),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(18)      => coldata_rx_inst_rx_parallel_data(18),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(19)      => coldata_rx_inst_rx_parallel_data(19),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(20)      => coldata_rx_inst_rx_parallel_data(20),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(21)      => coldata_rx_inst_rx_parallel_data(21),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(22)      => coldata_rx_inst_rx_parallel_data(22),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(23)      => coldata_rx_inst_rx_parallel_data(23),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(24)      => coldata_rx_inst_rx_parallel_data(24),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(25)      => coldata_rx_inst_rx_parallel_data(25),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(26)      => coldata_rx_inst_rx_parallel_data(26),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(27)      => coldata_rx_inst_rx_parallel_data(27),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(28)      => coldata_rx_inst_rx_parallel_data(28),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(29)      => coldata_rx_inst_rx_parallel_data(29),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(30)      => coldata_rx_inst_rx_parallel_data(30),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(31)      => coldata_rx_inst_rx_parallel_data(31),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(32)      => coldata_rx_inst_rx_parallel_data(32),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(33)      => coldata_rx_inst_rx_parallel_data(33),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(34)      => coldata_rx_inst_rx_parallel_data(34),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(35)      => coldata_rx_inst_rx_parallel_data(35),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(36)      => coldata_rx_inst_rx_parallel_data(36),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(37)      => coldata_rx_inst_rx_parallel_data(37),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(38)      => coldata_rx_inst_rx_parallel_data(38),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(39)      => coldata_rx_inst_rx_parallel_data(39),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(40)      => coldata_rx_inst_rx_parallel_data(40),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(41)      => coldata_rx_inst_rx_parallel_data(41),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(42)      => coldata_rx_inst_rx_parallel_data(42),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(43)      => coldata_rx_inst_rx_parallel_data(43),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(44)      => coldata_rx_inst_rx_parallel_data(44),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(45)      => coldata_rx_inst_rx_parallel_data(45),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(46)      => coldata_rx_inst_rx_parallel_data(46),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(47)      => coldata_rx_inst_rx_parallel_data(47),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(48)      => coldata_rx_inst_rx_parallel_data(48),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(49)      => coldata_rx_inst_rx_parallel_data(49),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(50)      => coldata_rx_inst_rx_parallel_data(50),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(51)      => coldata_rx_inst_rx_parallel_data(51),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(52)      => coldata_rx_inst_rx_parallel_data(52),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(53)      => coldata_rx_inst_rx_parallel_data(53),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(54)      => coldata_rx_inst_rx_parallel_data(54),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(55)      => coldata_rx_inst_rx_parallel_data(55),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(56)      => coldata_rx_inst_rx_parallel_data(56),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(57)      => coldata_rx_inst_rx_parallel_data(57),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(58)      => coldata_rx_inst_rx_parallel_data(58),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(59)      => coldata_rx_inst_rx_parallel_data(59),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(60)      => coldata_rx_inst_rx_parallel_data(60),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(61)      => coldata_rx_inst_rx_parallel_data(61),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(62)      => coldata_rx_inst_rx_parallel_data(62),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(63)      => coldata_rx_inst_rx_parallel_data(63),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(64)      => coldata_rx_inst_rx_parallel_data(64),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(65)      => coldata_rx_inst_rx_parallel_data(65),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(66)      => coldata_rx_inst_rx_parallel_data(66),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(67)      => coldata_rx_inst_rx_parallel_data(67),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(68)      => coldata_rx_inst_rx_parallel_data(68),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(69)      => coldata_rx_inst_rx_parallel_data(69),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(70)      => coldata_rx_inst_rx_parallel_data(70),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(71)      => coldata_rx_inst_rx_parallel_data(71),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(72)      => coldata_rx_inst_rx_parallel_data(72),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(73)      => coldata_rx_inst_rx_parallel_data(73),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(74)      => coldata_rx_inst_rx_parallel_data(74),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(75)      => coldata_rx_inst_rx_parallel_data(75),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(76)      => coldata_rx_inst_rx_parallel_data(76),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(77)      => coldata_rx_inst_rx_parallel_data(77),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(78)      => coldata_rx_inst_rx_parallel_data(78),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(79)      => coldata_rx_inst_rx_parallel_data(79),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(80)      => coldata_rx_inst_rx_parallel_data(80),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(81)      => coldata_rx_inst_rx_parallel_data(81),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(82)      => coldata_rx_inst_rx_parallel_data(82),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(83)      => coldata_rx_inst_rx_parallel_data(83),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(84)      => coldata_rx_inst_rx_parallel_data(84),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(85)      => coldata_rx_inst_rx_parallel_data(85),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(86)      => coldata_rx_inst_rx_parallel_data(86),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(87)      => coldata_rx_inst_rx_parallel_data(87),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(88)      => coldata_rx_inst_rx_parallel_data(88),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(89)      => coldata_rx_inst_rx_parallel_data(89),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(90)      => coldata_rx_inst_rx_parallel_data(90),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(91)      => coldata_rx_inst_rx_parallel_data(91),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(92)      => coldata_rx_inst_rx_parallel_data(92),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(93)      => coldata_rx_inst_rx_parallel_data(93),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(94)      => coldata_rx_inst_rx_parallel_data(94),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(95)      => coldata_rx_inst_rx_parallel_data(95),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(96)      => coldata_rx_inst_rx_parallel_data(96),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(97)      => coldata_rx_inst_rx_parallel_data(97),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(98)      => coldata_rx_inst_rx_parallel_data(98),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(99)      => coldata_rx_inst_rx_parallel_data(99),                                                                                                                                                                                                                                                                                               --                   .rx_parallel_data
			rx_parallel_data(100)     => coldata_rx_inst_rx_parallel_data(100),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(101)     => coldata_rx_inst_rx_parallel_data(101),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(102)     => coldata_rx_inst_rx_parallel_data(102),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(103)     => coldata_rx_inst_rx_parallel_data(103),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(104)     => coldata_rx_inst_rx_parallel_data(104),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(105)     => coldata_rx_inst_rx_parallel_data(105),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(106)     => coldata_rx_inst_rx_parallel_data(106),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(107)     => coldata_rx_inst_rx_parallel_data(107),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(108)     => coldata_rx_inst_rx_parallel_data(108),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(109)     => coldata_rx_inst_rx_parallel_data(109),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(110)     => coldata_rx_inst_rx_parallel_data(110),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(111)     => coldata_rx_inst_rx_parallel_data(111),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(112)     => coldata_rx_inst_rx_parallel_data(112),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(113)     => coldata_rx_inst_rx_parallel_data(113),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(114)     => coldata_rx_inst_rx_parallel_data(114),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(115)     => coldata_rx_inst_rx_parallel_data(115),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(116)     => coldata_rx_inst_rx_parallel_data(116),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(117)     => coldata_rx_inst_rx_parallel_data(117),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(118)     => coldata_rx_inst_rx_parallel_data(118),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(119)     => coldata_rx_inst_rx_parallel_data(119),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(120)     => coldata_rx_inst_rx_parallel_data(120),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(121)     => coldata_rx_inst_rx_parallel_data(121),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(122)     => coldata_rx_inst_rx_parallel_data(122),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(123)     => coldata_rx_inst_rx_parallel_data(123),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(124)     => coldata_rx_inst_rx_parallel_data(124),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(125)     => coldata_rx_inst_rx_parallel_data(125),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(126)     => coldata_rx_inst_rx_parallel_data(126),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(127)     => coldata_rx_inst_rx_parallel_data(127),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(128)     => coldata_rx_inst_rx_parallel_data(128),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(129)     => coldata_rx_inst_rx_parallel_data(129),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(130)     => coldata_rx_inst_rx_parallel_data(130),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(131)     => coldata_rx_inst_rx_parallel_data(131),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(132)     => coldata_rx_inst_rx_parallel_data(132),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(133)     => coldata_rx_inst_rx_parallel_data(133),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(134)     => coldata_rx_inst_rx_parallel_data(134),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(135)     => coldata_rx_inst_rx_parallel_data(135),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(136)     => coldata_rx_inst_rx_parallel_data(136),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(137)     => coldata_rx_inst_rx_parallel_data(137),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(138)     => coldata_rx_inst_rx_parallel_data(138),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(139)     => coldata_rx_inst_rx_parallel_data(139),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(140)     => coldata_rx_inst_rx_parallel_data(140),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(141)     => coldata_rx_inst_rx_parallel_data(141),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(142)     => coldata_rx_inst_rx_parallel_data(142),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(143)     => coldata_rx_inst_rx_parallel_data(143),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(144)     => coldata_rx_inst_rx_parallel_data(144),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(145)     => coldata_rx_inst_rx_parallel_data(145),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(146)     => coldata_rx_inst_rx_parallel_data(146),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(147)     => coldata_rx_inst_rx_parallel_data(147),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(148)     => coldata_rx_inst_rx_parallel_data(148),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(149)     => coldata_rx_inst_rx_parallel_data(149),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(150)     => coldata_rx_inst_rx_parallel_data(150),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(151)     => coldata_rx_inst_rx_parallel_data(151),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(152)     => coldata_rx_inst_rx_parallel_data(152),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(153)     => coldata_rx_inst_rx_parallel_data(153),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(154)     => coldata_rx_inst_rx_parallel_data(154),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(155)     => coldata_rx_inst_rx_parallel_data(155),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(156)     => coldata_rx_inst_rx_parallel_data(156),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(157)     => coldata_rx_inst_rx_parallel_data(157),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(158)     => coldata_rx_inst_rx_parallel_data(158),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(159)     => coldata_rx_inst_rx_parallel_data(159),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(160)     => coldata_rx_inst_rx_parallel_data(160),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(161)     => coldata_rx_inst_rx_parallel_data(161),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(162)     => coldata_rx_inst_rx_parallel_data(162),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(163)     => coldata_rx_inst_rx_parallel_data(163),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(164)     => coldata_rx_inst_rx_parallel_data(164),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(165)     => coldata_rx_inst_rx_parallel_data(165),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(166)     => coldata_rx_inst_rx_parallel_data(166),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(167)     => coldata_rx_inst_rx_parallel_data(167),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(168)     => coldata_rx_inst_rx_parallel_data(168),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(169)     => coldata_rx_inst_rx_parallel_data(169),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(170)     => coldata_rx_inst_rx_parallel_data(170),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(171)     => coldata_rx_inst_rx_parallel_data(171),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(172)     => coldata_rx_inst_rx_parallel_data(172),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(173)     => coldata_rx_inst_rx_parallel_data(173),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(174)     => coldata_rx_inst_rx_parallel_data(174),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(175)     => coldata_rx_inst_rx_parallel_data(175),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(176)     => coldata_rx_inst_rx_parallel_data(176),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(177)     => coldata_rx_inst_rx_parallel_data(177),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(178)     => coldata_rx_inst_rx_parallel_data(178),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(179)     => coldata_rx_inst_rx_parallel_data(179),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(180)     => coldata_rx_inst_rx_parallel_data(180),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(181)     => coldata_rx_inst_rx_parallel_data(181),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(182)     => coldata_rx_inst_rx_parallel_data(182),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(183)     => coldata_rx_inst_rx_parallel_data(183),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(184)     => coldata_rx_inst_rx_parallel_data(184),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(185)     => coldata_rx_inst_rx_parallel_data(185),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(186)     => coldata_rx_inst_rx_parallel_data(186),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(187)     => coldata_rx_inst_rx_parallel_data(187),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(188)     => coldata_rx_inst_rx_parallel_data(188),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(189)     => coldata_rx_inst_rx_parallel_data(189),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(190)     => coldata_rx_inst_rx_parallel_data(190),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(191)     => coldata_rx_inst_rx_parallel_data(191),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(192)     => coldata_rx_inst_rx_parallel_data(192),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(193)     => coldata_rx_inst_rx_parallel_data(193),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(194)     => coldata_rx_inst_rx_parallel_data(194),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(195)     => coldata_rx_inst_rx_parallel_data(195),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(196)     => coldata_rx_inst_rx_parallel_data(196),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(197)     => coldata_rx_inst_rx_parallel_data(197),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(198)     => coldata_rx_inst_rx_parallel_data(198),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(199)     => coldata_rx_inst_rx_parallel_data(199),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(200)     => coldata_rx_inst_rx_parallel_data(200),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(201)     => coldata_rx_inst_rx_parallel_data(201),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(202)     => coldata_rx_inst_rx_parallel_data(202),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(203)     => coldata_rx_inst_rx_parallel_data(203),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(204)     => coldata_rx_inst_rx_parallel_data(204),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(205)     => coldata_rx_inst_rx_parallel_data(205),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(206)     => coldata_rx_inst_rx_parallel_data(206),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(207)     => coldata_rx_inst_rx_parallel_data(207),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(208)     => coldata_rx_inst_rx_parallel_data(208),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(209)     => coldata_rx_inst_rx_parallel_data(209),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(210)     => coldata_rx_inst_rx_parallel_data(210),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(211)     => coldata_rx_inst_rx_parallel_data(211),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(212)     => coldata_rx_inst_rx_parallel_data(212),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(213)     => coldata_rx_inst_rx_parallel_data(213),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(214)     => coldata_rx_inst_rx_parallel_data(214),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(215)     => coldata_rx_inst_rx_parallel_data(215),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(216)     => coldata_rx_inst_rx_parallel_data(216),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(217)     => coldata_rx_inst_rx_parallel_data(217),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(218)     => coldata_rx_inst_rx_parallel_data(218),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(219)     => coldata_rx_inst_rx_parallel_data(219),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(220)     => coldata_rx_inst_rx_parallel_data(220),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(221)     => coldata_rx_inst_rx_parallel_data(221),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(222)     => coldata_rx_inst_rx_parallel_data(222),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(223)     => coldata_rx_inst_rx_parallel_data(223),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(224)     => coldata_rx_inst_rx_parallel_data(224),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(225)     => coldata_rx_inst_rx_parallel_data(225),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(226)     => coldata_rx_inst_rx_parallel_data(226),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(227)     => coldata_rx_inst_rx_parallel_data(227),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(228)     => coldata_rx_inst_rx_parallel_data(228),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(229)     => coldata_rx_inst_rx_parallel_data(229),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(230)     => coldata_rx_inst_rx_parallel_data(230),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(231)     => coldata_rx_inst_rx_parallel_data(231),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(232)     => coldata_rx_inst_rx_parallel_data(232),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(233)     => coldata_rx_inst_rx_parallel_data(233),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(234)     => coldata_rx_inst_rx_parallel_data(234),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(235)     => coldata_rx_inst_rx_parallel_data(235),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(236)     => coldata_rx_inst_rx_parallel_data(236),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(237)     => coldata_rx_inst_rx_parallel_data(237),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(238)     => coldata_rx_inst_rx_parallel_data(238),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(239)     => coldata_rx_inst_rx_parallel_data(239),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(240)     => coldata_rx_inst_rx_parallel_data(240),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(241)     => coldata_rx_inst_rx_parallel_data(241),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(242)     => coldata_rx_inst_rx_parallel_data(242),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(243)     => coldata_rx_inst_rx_parallel_data(243),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(244)     => coldata_rx_inst_rx_parallel_data(244),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(245)     => coldata_rx_inst_rx_parallel_data(245),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(246)     => coldata_rx_inst_rx_parallel_data(246),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(247)     => coldata_rx_inst_rx_parallel_data(247),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(248)     => coldata_rx_inst_rx_parallel_data(248),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(249)     => coldata_rx_inst_rx_parallel_data(249),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(250)     => coldata_rx_inst_rx_parallel_data(250),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(251)     => coldata_rx_inst_rx_parallel_data(251),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(252)     => coldata_rx_inst_rx_parallel_data(252),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(253)     => coldata_rx_inst_rx_parallel_data(253),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(254)     => coldata_rx_inst_rx_parallel_data(254),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			rx_parallel_data(255)     => coldata_rx_inst_rx_parallel_data(255),                                                                                                                                                                                                                                                                                              --                   .rx_parallel_data
			pll_powerdown             => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_analogreset            => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_digitalreset           => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_pll_refclk             => "0",                                                                                                                                                                                                                                                                                                                                --        (terminated)
			tx_pma_clkout             => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_serial_data            => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_parallel_data      => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			pll_locked                => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			ext_pll_clk               => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_pma_clkout             => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_parallel_data      => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_clkslip                => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_clklow                 => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_fref                   => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_set_locktodata         => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_set_locktoref          => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_seriallpbken           => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_signaldetect           => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_parallel_data          => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",                                                                                                                                                 --        (terminated)
			tx_std_coreclkin          => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_std_clkout             => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_done          => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_err           => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_byteorder_ena      => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_byteorder_flag     => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_full        => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty       => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign    => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_wa_a1a2size        => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_std_bitslipboundarysel => "00000000000000000000",                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_bitslipboundarysel => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitslip            => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_runlength_err      => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena         => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_byterev_ena        => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_std_polinv             => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_polinv             => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_std_elecidle           => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_signaldetect       => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_cal_busy               => open                                                                                                                                                                                                                                                                                                                                --        (terminated)
		);

	rx_syncstatus <= COLDATA_RX_inst_rx_parallel_data(202) & COLDATA_RX_inst_rx_parallel_data(138) & COLDATA_RX_inst_rx_parallel_data(74) & COLDATA_RX_inst_rx_parallel_data(10);

	rx_runningdisp <= COLDATA_RX_inst_rx_parallel_data(207) & COLDATA_RX_inst_rx_parallel_data(143) & COLDATA_RX_inst_rx_parallel_data(79) & COLDATA_RX_inst_rx_parallel_data(15);

	rx_patterndetect <= COLDATA_RX_inst_rx_parallel_data(204) & COLDATA_RX_inst_rx_parallel_data(140) & COLDATA_RX_inst_rx_parallel_data(76) & COLDATA_RX_inst_rx_parallel_data(12);

	rx_disperr <= COLDATA_RX_inst_rx_parallel_data(203) & COLDATA_RX_inst_rx_parallel_data(139) & COLDATA_RX_inst_rx_parallel_data(75) & COLDATA_RX_inst_rx_parallel_data(11);

	rx_errdetect <= COLDATA_RX_inst_rx_parallel_data(201) & COLDATA_RX_inst_rx_parallel_data(137) & COLDATA_RX_inst_rx_parallel_data(73) & COLDATA_RX_inst_rx_parallel_data(9);

	unused_rx_parallel_data <= COLDATA_RX_inst_rx_parallel_data(255) & COLDATA_RX_inst_rx_parallel_data(254) & COLDATA_RX_inst_rx_parallel_data(253) & COLDATA_RX_inst_rx_parallel_data(252) & COLDATA_RX_inst_rx_parallel_data(251) & COLDATA_RX_inst_rx_parallel_data(250) & COLDATA_RX_inst_rx_parallel_data(249) & COLDATA_RX_inst_rx_parallel_data(248) & COLDATA_RX_inst_rx_parallel_data(247) & COLDATA_RX_inst_rx_parallel_data(246) & COLDATA_RX_inst_rx_parallel_data(245) & COLDATA_RX_inst_rx_parallel_data(244) & COLDATA_RX_inst_rx_parallel_data(243) & COLDATA_RX_inst_rx_parallel_data(242) & COLDATA_RX_inst_rx_parallel_data(241) & COLDATA_RX_inst_rx_parallel_data(240) & COLDATA_RX_inst_rx_parallel_data(239) & COLDATA_RX_inst_rx_parallel_data(238) & COLDATA_RX_inst_rx_parallel_data(237) & COLDATA_RX_inst_rx_parallel_data(236) & COLDATA_RX_inst_rx_parallel_data(235) & COLDATA_RX_inst_rx_parallel_data(234) & COLDATA_RX_inst_rx_parallel_data(233) & COLDATA_RX_inst_rx_parallel_data(232) & COLDATA_RX_inst_rx_parallel_data(231) & COLDATA_RX_inst_rx_parallel_data(230) & COLDATA_RX_inst_rx_parallel_data(229) & COLDATA_RX_inst_rx_parallel_data(228) & COLDATA_RX_inst_rx_parallel_data(227) & COLDATA_RX_inst_rx_parallel_data(226) & COLDATA_RX_inst_rx_parallel_data(225) & COLDATA_RX_inst_rx_parallel_data(224) & COLDATA_RX_inst_rx_parallel_data(223) & COLDATA_RX_inst_rx_parallel_data(222) & COLDATA_RX_inst_rx_parallel_data(221) & COLDATA_RX_inst_rx_parallel_data(220) & COLDATA_RX_inst_rx_parallel_data(219) & COLDATA_RX_inst_rx_parallel_data(218) & COLDATA_RX_inst_rx_parallel_data(217) & COLDATA_RX_inst_rx_parallel_data(216) & COLDATA_RX_inst_rx_parallel_data(215) & COLDATA_RX_inst_rx_parallel_data(214) & COLDATA_RX_inst_rx_parallel_data(213) & COLDATA_RX_inst_rx_parallel_data(212) & COLDATA_RX_inst_rx_parallel_data(211) & COLDATA_RX_inst_rx_parallel_data(210) & COLDATA_RX_inst_rx_parallel_data(209) & COLDATA_RX_inst_rx_parallel_data(208) & COLDATA_RX_inst_rx_parallel_data(206) & COLDATA_RX_inst_rx_parallel_data(205) & COLDATA_RX_inst_rx_parallel_data(191) & COLDATA_RX_inst_rx_parallel_data(190) & COLDATA_RX_inst_rx_parallel_data(189) & COLDATA_RX_inst_rx_parallel_data(188) & COLDATA_RX_inst_rx_parallel_data(187) & COLDATA_RX_inst_rx_parallel_data(186) & COLDATA_RX_inst_rx_parallel_data(185) & COLDATA_RX_inst_rx_parallel_data(184) & COLDATA_RX_inst_rx_parallel_data(183) & COLDATA_RX_inst_rx_parallel_data(182) & COLDATA_RX_inst_rx_parallel_data(181) & COLDATA_RX_inst_rx_parallel_data(180) & COLDATA_RX_inst_rx_parallel_data(179) & COLDATA_RX_inst_rx_parallel_data(178) & COLDATA_RX_inst_rx_parallel_data(177) & COLDATA_RX_inst_rx_parallel_data(176) & COLDATA_RX_inst_rx_parallel_data(175) & COLDATA_RX_inst_rx_parallel_data(174) & COLDATA_RX_inst_rx_parallel_data(173) & COLDATA_RX_inst_rx_parallel_data(172) & COLDATA_RX_inst_rx_parallel_data(171) & COLDATA_RX_inst_rx_parallel_data(170) & COLDATA_RX_inst_rx_parallel_data(169) & COLDATA_RX_inst_rx_parallel_data(168) & COLDATA_RX_inst_rx_parallel_data(167) & COLDATA_RX_inst_rx_parallel_data(166) & COLDATA_RX_inst_rx_parallel_data(165) & COLDATA_RX_inst_rx_parallel_data(164) & COLDATA_RX_inst_rx_parallel_data(163) & COLDATA_RX_inst_rx_parallel_data(162) & COLDATA_RX_inst_rx_parallel_data(161) & COLDATA_RX_inst_rx_parallel_data(160) & COLDATA_RX_inst_rx_parallel_data(159) & COLDATA_RX_inst_rx_parallel_data(158) & COLDATA_RX_inst_rx_parallel_data(157) & COLDATA_RX_inst_rx_parallel_data(156) & COLDATA_RX_inst_rx_parallel_data(155) & COLDATA_RX_inst_rx_parallel_data(154) & COLDATA_RX_inst_rx_parallel_data(153) & COLDATA_RX_inst_rx_parallel_data(152) & COLDATA_RX_inst_rx_parallel_data(151) & COLDATA_RX_inst_rx_parallel_data(150) & COLDATA_RX_inst_rx_parallel_data(149) & COLDATA_RX_inst_rx_parallel_data(148) & COLDATA_RX_inst_rx_parallel_data(147) & COLDATA_RX_inst_rx_parallel_data(146) & COLDATA_RX_inst_rx_parallel_data(145) & COLDATA_RX_inst_rx_parallel_data(144) & COLDATA_RX_inst_rx_parallel_data(142) & COLDATA_RX_inst_rx_parallel_data(141) & COLDATA_RX_inst_rx_parallel_data(127) & COLDATA_RX_inst_rx_parallel_data(126) & COLDATA_RX_inst_rx_parallel_data(125) & COLDATA_RX_inst_rx_parallel_data(124) & COLDATA_RX_inst_rx_parallel_data(123) & COLDATA_RX_inst_rx_parallel_data(122) & COLDATA_RX_inst_rx_parallel_data(121) & COLDATA_RX_inst_rx_parallel_data(120) & COLDATA_RX_inst_rx_parallel_data(119) & COLDATA_RX_inst_rx_parallel_data(118) & COLDATA_RX_inst_rx_parallel_data(117) & COLDATA_RX_inst_rx_parallel_data(116) & COLDATA_RX_inst_rx_parallel_data(115) & COLDATA_RX_inst_rx_parallel_data(114) & COLDATA_RX_inst_rx_parallel_data(113) & COLDATA_RX_inst_rx_parallel_data(112) & COLDATA_RX_inst_rx_parallel_data(111) & COLDATA_RX_inst_rx_parallel_data(110) & COLDATA_RX_inst_rx_parallel_data(109) & COLDATA_RX_inst_rx_parallel_data(108) & COLDATA_RX_inst_rx_parallel_data(107) & COLDATA_RX_inst_rx_parallel_data(106) & COLDATA_RX_inst_rx_parallel_data(105) & COLDATA_RX_inst_rx_parallel_data(104) & COLDATA_RX_inst_rx_parallel_data(103) & COLDATA_RX_inst_rx_parallel_data(102) & COLDATA_RX_inst_rx_parallel_data(101) & COLDATA_RX_inst_rx_parallel_data(100) & COLDATA_RX_inst_rx_parallel_data(99) & COLDATA_RX_inst_rx_parallel_data(98) & COLDATA_RX_inst_rx_parallel_data(97) & COLDATA_RX_inst_rx_parallel_data(96) & COLDATA_RX_inst_rx_parallel_data(95) & COLDATA_RX_inst_rx_parallel_data(94) & COLDATA_RX_inst_rx_parallel_data(93) & COLDATA_RX_inst_rx_parallel_data(92) & COLDATA_RX_inst_rx_parallel_data(91) & COLDATA_RX_inst_rx_parallel_data(90) & COLDATA_RX_inst_rx_parallel_data(89) & COLDATA_RX_inst_rx_parallel_data(88) & COLDATA_RX_inst_rx_parallel_data(87) & COLDATA_RX_inst_rx_parallel_data(86) & COLDATA_RX_inst_rx_parallel_data(85) & COLDATA_RX_inst_rx_parallel_data(84) & COLDATA_RX_inst_rx_parallel_data(83) & COLDATA_RX_inst_rx_parallel_data(82) & COLDATA_RX_inst_rx_parallel_data(81) & COLDATA_RX_inst_rx_parallel_data(80) & COLDATA_RX_inst_rx_parallel_data(78) & COLDATA_RX_inst_rx_parallel_data(77) & COLDATA_RX_inst_rx_parallel_data(63) & COLDATA_RX_inst_rx_parallel_data(62) & COLDATA_RX_inst_rx_parallel_data(61) & COLDATA_RX_inst_rx_parallel_data(60) & COLDATA_RX_inst_rx_parallel_data(59) & COLDATA_RX_inst_rx_parallel_data(58) & COLDATA_RX_inst_rx_parallel_data(57) & COLDATA_RX_inst_rx_parallel_data(56) & COLDATA_RX_inst_rx_parallel_data(55) & COLDATA_RX_inst_rx_parallel_data(54) & COLDATA_RX_inst_rx_parallel_data(53) & COLDATA_RX_inst_rx_parallel_data(52) & COLDATA_RX_inst_rx_parallel_data(51) & COLDATA_RX_inst_rx_parallel_data(50) & COLDATA_RX_inst_rx_parallel_data(49) & COLDATA_RX_inst_rx_parallel_data(48) & COLDATA_RX_inst_rx_parallel_data(47) & COLDATA_RX_inst_rx_parallel_data(46) & COLDATA_RX_inst_rx_parallel_data(45) & COLDATA_RX_inst_rx_parallel_data(44) & COLDATA_RX_inst_rx_parallel_data(43) & COLDATA_RX_inst_rx_parallel_data(42) & COLDATA_RX_inst_rx_parallel_data(41) & COLDATA_RX_inst_rx_parallel_data(40) & COLDATA_RX_inst_rx_parallel_data(39) & COLDATA_RX_inst_rx_parallel_data(38) & COLDATA_RX_inst_rx_parallel_data(37) & COLDATA_RX_inst_rx_parallel_data(36) & COLDATA_RX_inst_rx_parallel_data(35) & COLDATA_RX_inst_rx_parallel_data(34) & COLDATA_RX_inst_rx_parallel_data(33) & COLDATA_RX_inst_rx_parallel_data(32) & COLDATA_RX_inst_rx_parallel_data(31) & COLDATA_RX_inst_rx_parallel_data(30) & COLDATA_RX_inst_rx_parallel_data(29) & COLDATA_RX_inst_rx_parallel_data(28) & COLDATA_RX_inst_rx_parallel_data(27) & COLDATA_RX_inst_rx_parallel_data(26) & COLDATA_RX_inst_rx_parallel_data(25) & COLDATA_RX_inst_rx_parallel_data(24) & COLDATA_RX_inst_rx_parallel_data(23) & COLDATA_RX_inst_rx_parallel_data(22) & COLDATA_RX_inst_rx_parallel_data(21) & COLDATA_RX_inst_rx_parallel_data(20) & COLDATA_RX_inst_rx_parallel_data(19) & COLDATA_RX_inst_rx_parallel_data(18) & COLDATA_RX_inst_rx_parallel_data(17) & COLDATA_RX_inst_rx_parallel_data(16) & COLDATA_RX_inst_rx_parallel_data(14) & COLDATA_RX_inst_rx_parallel_data(13);

	rx_parallel_data <= COLDATA_RX_inst_rx_parallel_data(199) & COLDATA_RX_inst_rx_parallel_data(198) & COLDATA_RX_inst_rx_parallel_data(197) & COLDATA_RX_inst_rx_parallel_data(196) & COLDATA_RX_inst_rx_parallel_data(195) & COLDATA_RX_inst_rx_parallel_data(194) & COLDATA_RX_inst_rx_parallel_data(193) & COLDATA_RX_inst_rx_parallel_data(192) & COLDATA_RX_inst_rx_parallel_data(135) & COLDATA_RX_inst_rx_parallel_data(134) & COLDATA_RX_inst_rx_parallel_data(133) & COLDATA_RX_inst_rx_parallel_data(132) & COLDATA_RX_inst_rx_parallel_data(131) & COLDATA_RX_inst_rx_parallel_data(130) & COLDATA_RX_inst_rx_parallel_data(129) & COLDATA_RX_inst_rx_parallel_data(128) & COLDATA_RX_inst_rx_parallel_data(71) & COLDATA_RX_inst_rx_parallel_data(70) & COLDATA_RX_inst_rx_parallel_data(69) & COLDATA_RX_inst_rx_parallel_data(68) & COLDATA_RX_inst_rx_parallel_data(67) & COLDATA_RX_inst_rx_parallel_data(66) & COLDATA_RX_inst_rx_parallel_data(65) & COLDATA_RX_inst_rx_parallel_data(64) & COLDATA_RX_inst_rx_parallel_data(7) & COLDATA_RX_inst_rx_parallel_data(6) & COLDATA_RX_inst_rx_parallel_data(5) & COLDATA_RX_inst_rx_parallel_data(4) & COLDATA_RX_inst_rx_parallel_data(3) & COLDATA_RX_inst_rx_parallel_data(2) & COLDATA_RX_inst_rx_parallel_data(1) & COLDATA_RX_inst_rx_parallel_data(0);

	rx_datak <= COLDATA_RX_inst_rx_parallel_data(200) & COLDATA_RX_inst_rx_parallel_data(136) & COLDATA_RX_inst_rx_parallel_data(72) & COLDATA_RX_inst_rx_parallel_data(8);

end architecture rtl; -- of COLDATA_RX
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2017 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_xcvr_native_av" version="16.0" >
-- Retrieval info: 	<generic name="device_family" value="Arria V" />
-- Retrieval info: 	<generic name="show_advanced_features" value="0" />
-- Retrieval info: 	<generic name="device_speedgrade" value="fastest" />
-- Retrieval info: 	<generic name="message_level" value="error" />
-- Retrieval info: 	<generic name="tx_enable" value="0" />
-- Retrieval info: 	<generic name="rx_enable" value="1" />
-- Retrieval info: 	<generic name="enable_std" value="1" />
-- Retrieval info: 	<generic name="set_data_path_select" value="standard" />
-- Retrieval info: 	<generic name="channels" value="4" />
-- Retrieval info: 	<generic name="bonded_mode" value="non_bonded" />
-- Retrieval info: 	<generic name="enable_simple_interface" value="1" />
-- Retrieval info: 	<generic name="set_data_rate" value="1280" />
-- Retrieval info: 	<generic name="pma_direct_width" value="80" />
-- Retrieval info: 	<generic name="tx_pma_clk_div" value="1" />
-- Retrieval info: 	<generic name="pll_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="pll_external_enable" value="0" />
-- Retrieval info: 	<generic name="plls" value="1" />
-- Retrieval info: 	<generic name="pll_select" value="0" />
-- Retrieval info: 	<generic name="pll_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="cdr_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_refclk_select" value="0" />
-- Retrieval info: 	<generic name="set_cdr_refclk_freq" value="128.0 MHz" />
-- Retrieval info: 	<generic name="rx_ppm_detect_threshold" value="1000" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_clkout" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtodata" value="1" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtoref" value="1" />
-- Retrieval info: 	<generic name="enable_ports_rx_manual_cdr_mode" value="0" />
-- Retrieval info: 	<generic name="rx_clkslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_seriallpbken" value="0" />
-- Retrieval info: 	<generic name="std_protocol_hint" value="basic" />
-- Retrieval info: 	<generic name="std_pcs_pma_width" value="10" />
-- Retrieval info: 	<generic name="std_low_latency_bypass_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_pcfifo_mode" value="low_latency" />
-- Retrieval info: 	<generic name="std_rx_pcfifo_mode" value="low_latency" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_mode" value="manual" />
-- Retrieval info: 	<generic name="std_rx_byte_order_symbol_count" value="1" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pattern" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pad" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_flag" value="0" />
-- Retrieval info: 	<generic name="std_tx_byte_ser_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_deser_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_8b10b_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_8b10b_disp_ctrl_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_8b10b_enable" value="1" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_p" value="27c" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_n" value="27c" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_mode" value="sync_sm" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern_len" value="10" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern" value="27c" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rknumber" value="5" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_renumber" value="5" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rgnumber" value="5" />
-- Retrieval info: 	<generic name="std_rx_run_length_val" value="10" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_patternalign" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_a1a2size" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_runlength_err" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitrev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byterev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_polinv" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_polinv" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_elecidle" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_prbs_status" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_clk_network" value="x1" />
-- Retrieval info: </instance>
-- IPFS_FILES : COLDATA_RX.vho
-- RELATED_FILES: COLDATA_RX.vhd, altera_xcvr_functions.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_native_av_functions_h.sv, altera_xcvr_native_av.sv, altera_xcvr_data_adapter_av.sv
