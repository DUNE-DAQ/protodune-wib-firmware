// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IEWZFElpTRFKDtLY2a66xnyCuC9SJTb9kdxcoRyEk78W0dc5eSfx0on1IXHu3pmQ
u5e6rbB7q0KtQ83GY3m1WggePv6a4v+EQIltAIOEB4y9yrnx1j7aD4MUFMG6h17x
yVjg0cAesx1nukqM2tF+njkzIt4Mk1IggeqNpvx4110=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48608)
4GobaLel80iR6BSUZU3hcvg5eqkB+Zzu0PeXJQ/6pm2Mx914sVh7JKtdhXEtkvz/
7W9Q3PPYFldaZysVOEaSbIdV4O8lClMeRw3t0fgc8jwr/JTGUd8qiiaJH5TJzu/p
qpWvqvr29pJ0SdXE6NEeQkIKhMqSVx0GT71R7sI65sTPmiL+36GidMBykbxCP5nS
YmhDdkJlvEqMPcChTTzpBTbRTBTCfsYmERosDrBpwBonRO2YrMJzvgvr+mNT6zmS
9Iq5iL4H+1B+YkTQ4Uk22VsEdU+juThTTp1I1NUizZ67lGMXsJoD91fSDiMnU6lO
s5NgQOwee/XQp+RSlCSIo7lrPBCgjePPtREO05aG4sM7W0Q513PJ+Kbmd7pi5oHm
rJvpiDgtQ6YTEAz0b1uuirLZK/EOQTznRzRiVZ3oAxq95rexsAzB3JE6IH25PUOr
YfuZbNKrwS2wdDkdEt+2bTC3J/HHn7u0rCI4B3sg+q2s2i3V/9EuuiC/sOfktQss
bHU8P16ugNnJfVLB2jMtEfRV5zeK661SusGHor+c3fwdnDcJtUxZkZYnaabuWSlJ
FcVKPXtjfOLoW+7IlnwQHKmAigGPG0EvZBOmWrZz1kVx/aLTMTCUHkADYMCwhnvV
RF6LJtV6ghf2P6o/+v/WJLK6kaHUxQO9YTCEoGDEye4AyB/vh4xLUoGG/ChddzrB
KAbZAmUaxcbQp1cfWXSYNZQKSHCKdE879gr1gIkhylv4nsQkPFfzjz/ho22g+uBx
WkAHq6CKG1UDjYLiY2l+ekDNiX5OqdNAiPEhI8mF784odfHimCLfs0grKpDRY5sy
/4yF0aq9V086pl7RGVL8kssy9Q1iyQbStgV0CLJcF4fQVWp0IpHjbilFSq+h2jhh
Ua/xWtFxGQWsVRefmXMacuplbkak/xFUZODXcdS6+8ryhNgZHnUyY4vV3OEz0uiK
NJTxFgDnr1D/4E52mrkZLsdpg2bza3La47+iL5raLJmnWkqwYlXt0q4FK7P0lohk
EtS30PuS93P/TytHZajfDbeQSoJnNeJ3GKxAXs/T6aiHYhP20r0coHPcRZyb6hPy
8s+boLu/5E1gkJCfoFzKoCslJ+VFsaWDipyUW+Umy94NdZSDvkCzVPpdwYNusTZI
mZvUPkB7ashjVXH4fTQ1rwrQS/6bpg/hrt/hc9Brjc3bIepil0uR0jo9Kl/tSRHv
pwmJG6HFykQLrTf0UNRz+v9i1B26VkEKJzbWRiBfO2jmw2NZNX64fAyPDCZhHP4Q
rHyVBJrh5VnV/77iWtZskRLUGeTkb7LF/YudjoKxCZNA6RF8yVw89cyCySTcwYUE
jCW6Ht9jh4m1p26miFQ7I2c2kSfYjRSmJBcsM5/GhLikVs2ssQjdCd9XfU/tEMFl
IEm0C7WOgBvcPN+Ofc78Z6EIuT2j5nDw7uRW7aNsk3nnbjvINaAmHmF+EgdPfaRU
8ZQj24VudAZtf7FTzs1XacpP6i+P6Sqc1cqxruoy5pk5dSZEohelymkJuuyyYtjC
QCPttrBrAycdJjK+6w+iPBLJWPXFrc6zGUniYKJHt/HBFdLB5uh7kv2PWn658uCQ
H/5sQ4Oy5BZrS3j3A3TsLQJAbGJzdRZDRjOQ5dxLestcEj+5p8DCZqeDmoVE0MJW
TPYNpFNVvymlyBhYs+slTJSvgdNCHlkCCXO7YZU1jN+hDAFrEDzjINP2RdzBtZLI
97eByBNhXrdUXgugS1eQza++j5JCes3UOfH9RxLXjIm7IgyhAKhTTFYtgTJgVFLJ
1A5qFANg3sgheVpkMNCGqSLPdhM9CRKRt5GyCeRWoF1YUFz1+8WW0h9hKYt+c/wG
gZ2IFN9JeVkf+GZIAKuvsQluAkJGfbsbcuu7I8LZh1Cc/9I9f6lt7lQQ/Y46FsKE
nAaMOJCqGYGC7q4mLOcSt7FP1BOcokXGGqI0j602H4wPXS9s4gpX3xhISQwn9A45
oWqsFO/P8CmDBSeCxVYYfv8kJux7V3HUFtd5V3wL0TOPisHn885HtiJHrx1YtN5m
C5Zve9+EBSFqa5F31+eOaZzNVx2RKxLGwcw6vRmsgU/CEfIgpya2tvvBJCQ15w/w
IPxSyZdnAju29A4YdwNT4bTvjCjirTUdVxIrKud8CrVwm0x/QZRWoBG/m+QNx1BJ
j5LoNJwG4r1VkZNM479OaRhv2Rr7WH2ZkJrne7JRejIEi5oTKG/pVGXx7R6R+/W7
p4q9FBhh+DLIoprgI5p3bfaDWPRKTf24pdGXYxgr2uS14iNh4/JPGFGnkPMTCnhV
VWAIXhJhIotZWFmZUiKnlEHSZTp6MzVAPFe2uXQKuTz+UGRaX8F2K467Umqz5S1X
DVOSnPVhk7efmXLAqsnyMaCDhlr9vhQtRSasPXL4NcS/k87ksnHB2sKwCJy9qWrZ
YIXU1TdJJjIyj9fJwv4mh+0GsCt8wtWrx2kmP8n2KWDtcEzBYZS1Voj8ocN7SDZ9
Nhpwy3TJ9srS0ik/NsNlXUhHTyCymWdM6h1viC5K1WZg6Ypwfd/ysV4bF+uBYRcO
D1gPrhsF2G1NR0n3yhT1MCI2Bss+aIkB4DYO+41483Jd6+d/sYrGn5daaa3AcAE4
WO3uR0jt13VJJ0kwAwORzlQhqr8aekDHDfqcdrdE5+PzLWL4BLZxaJLeQGjGuuXv
3jbGbc5poTPAplCooq8NUknaMdCdC8u2HNY4JZTFtq5Jf4xwsuutOQdrfYy0xPNc
ykeMQyKF3muB/bfNG+yqwBfkcUV8QVJPgML7VwbWl1gPCvLWyRciBinSb5TRVjZu
29WkwmJC4iku4lx3kdC+BV3uo9YwHUKaigKRH0sJjLfxQ8nSLVTZwv9z85Rh5Tbj
IPN+S6DOMYqNNb6aiZAkOWraEW0yftEbtpoj/HhdLfm4lVfisznEkNzfqZC/pQt5
g7sUolCPtLIU73PNCURNAtFEPpEdqUN4kS5jWtFfJUq9z5q8+cvDb0FfhqpeqFk3
kXJ78dmAeiduOWVzqPvmbRyRxGcbTdp+Zk/HuDghvET4jwEDaT5lnN9JoRXnX5bc
Lne80OGZ++3WTR/vBnbIMMEqh48JfLQEJtnLZmtH5suEjRxvIMzVftdRkZi1akJV
rQvOdoO+xzGwef47hC3warWxRRojcN6OfQuRggwqXXarIpQsHGqFpRfwyuDdSH4Z
a9sbYYUMgTI9SLvvH2Vq6FdykgQzP4U44XY0n6jT5yESejjdnmwsfn6Qt1ydnlPd
55dRt6tJvQ7zbCywtEsidLwj4+x0bE7zjFORLLCR3N5/suMMwGaGQJxiEPD9hHY9
2lNewgLgspYalFTHjed8XnWQ7OP98Az/iy/+TfMbW8ymB96hKjQBzlO2Mpkz7EVQ
bARgWzIcln+fyNX9CftnV3x/deoW27+ArWzuQluFbbL4+GxTR3SVAp+WZsOU2Rf9
5lYmBGuQgSZ3g2NgM2IODxu1RCvT1tU1t9tX5shahUfCQ+vX1Dbeu27ws4Vam6u0
55yOLISXzd0YNQGWGDjyPcxl3yk4vj9dpxgr5z37C1Jnw5fYuYBd8zZEACKR1Bj9
ETC1p6UCAjJLzXaUhEV3U5uxeRJlC5Bdure87UvwFOSH3ih4O+L+guGJ/NRIBwLV
deQOgq6ZOMncv21s5qZKamwJWHmtCtWoXcb5lpDwzg4Ff/N6h4vrZDZaGlW0/GBp
eIHWc8ZbP30HnzXZ8vHNh3PbKQGsp86pWW3gtCnnU8xZ/IfvH6OsLaFN55bY62K9
1mcU8zLdm16jlo4u21iuYbrbmrk7v5tFycDIJz3LWyOjHtoAnS4MkbvQDatR6DBq
yY4cnoqYwcbr8tJuoifABGKqmbHDrKo/meePA9S/hkuDwi4B2lsMOH7SBhnNcK5w
zJjFo2HWiUXqlEnYQjAUoGxrI0tU2ovrC8Dm9pd2TgY/R6Gdg0Q1A3EhIv5MQu1i
0YLxZMVGtc7fRzVnNj0qdT2G6CXgihUCxi60IMvZYRgW5STBAq2FGKZrOu0PJv4I
l1a9XProZdlQBZAWppfYoCVlv6Jhdg/7ka6fGV6jicmKfSE5WHC0ncXAqWRXfd5Z
AeFfZjpZ3TkFvoiTVwfMuKST8qchq3jHefRwpn8p2x4aKt5U4OrDCc/TSB4nldQ4
pcUHcJ92SIOBQAE/Tjyjyd3DBlOsXx2hA6sdmhBfWj4Pkw0JCrVOHelBMWMbXryd
mkLlAvF3nJpM+ReK3eH5NcYmCEh3LhYqNT/P2EWNYoGNS5ISoxbXuEXL+e7glSGL
8mAoemL6YUxIXMbNOZluOq0UxkIwDW5WXTPDshWu9C/O14x8/gDoiID0nzO3MeA9
2+xDkQxDPvcs9Ui6dXm2tJL4j08iTjVcE1Bk7LFwQJaP7JeL906+o0hqUGcJ7N9X
8YRpO5nDOe3JUoMejhnMN47JURY/sZwfv5lpbIKip0A5mSfU5DFafuP8HDwtwLPu
RRWAOa4hqhc0jj+tJ8QuwpXxxaWa/fcIRX30QDknl4tQRfDcR1eT5Jq6mAZgsXoE
U9WoHydFJkIq9UOHsG3Yftsml71nthFpFLuX/o5ptN+4otv4eQx/JNYkSh4Pk8j/
mkjJuCQZMMykHIIptoqPuBSpNNFSRFZUl6gEPUylgjE463xuyX6JCoraSID9YAD4
z0SWC+49bGQ/p8tUS1Mo7UhFE3nIM3TuGNz9NLfWKBrmxEBfpFLaKE84U395dBHE
KdzHyDNrCRowXJYZzcoXq5ueVwq3212eOvopFRylHY7jg6pZ+AkBUkzHMe0LjYWl
TynCTVU3Bey/ECdWsCEQFW+EQMbgtc5BMBzc4jwgUcYiwxvQfjYMzX2NPA7jzkjA
I5ATafh6gziuo4uqGGd8XFhrbFB8zxY57iz6y7dfCNS/Am0HXPRDOEH1/u8Onzcx
illqcd7IOeN1Cn54bnfnJiBN7LgLJIdIPtebpzdFDkwYU2LirfqYF8sWmpKib0bA
wmR1ggeXKuXZKYzUBKTCG88JaCGdVCc/IT0+XVZNkwAPBMVpMSiC1n4T9FiHH5c6
GC5FesnAS1CJDUHfYhToXpzW9itwJvVhGEG/atLeQt6XRlHB7Ixe1MA7BO1hRI8L
44dB25gFq5ZCs3Tj+i4bz9lkSQXeP+bsATICAbtqQ/XEJwA5F4GbQoX0Yn5Gcrok
IF6vW2mrUFNFboHmpdcg6SVkXSR84d9QJWNiH5qdKR4xJZiS7X/pN0E0mC4CGG6g
F+AMfGsrNlEp4Suvz5w9g0MUlEkNnx6L6T8ZrCeHVDtkUsafqG5QZhPc9VJecDnt
l1yTknFQoTCctjznvVWEWYgKVt90QSeqDoNMh+QTKopYBCC4D/Z+D/lAAfPt9swx
5scK3QI2bopoeupH3u33SjmGtOoaiZzay+sBKS9DomorhMMjPV1KEe9ZUAkLWvRU
mRncTC9MqO32UV/PZzyE9VsXPFZVUTvrAl7fqN+TrTYXvmYCkUGSsWIsxJ3M18HS
0K1wAkNfP7LDum9khTvYQZxG+117ByYgi17Um+4gC1nvtMHWdCI6uNNoM/PD1sa6
AL7ALVgN0y0eBcH/hk6j0PIeg/msXlnb/4JHc7bft6zTipymnhWUofeOpz+uQdO0
JzhVYZUHGvYOWEfcO5+mCa59jmfsmyTEXLxOVCjwRjuYa5OmDLniytGVjwYVw2AO
HAcIBiFUVfs8SZMD8Qis/1TJwfe38T8TMeEiEFNiRG9U42neTnI2yqQZGEoi+FlX
rvR/IzfHTDk2vKjtFjT5cGVlV/FGyhcn0m+G5fg/TzJ3iEovXXwGLFFGm2iwgmN6
Nfl+dME2Jgo891vLRMIztutpo85C+nBxVtVzWW+bB7okCSOTiHSZ+oFOV1pOLsDw
6bD80GExF1QJK1iSPLSBXuZi1g29lslrev0hkL+r/LCuwBuEvDXp/6QZMSFx0fAJ
PoYsQ6L7cHUxbZrFddeRvkYzUmcYKrawe2gJlZFjejrf2PVndBag/EiOD8ckfWSz
ZWrNJOfEthIuw1KSfSuOlTt3lQrG+kVjU2kUU+SNmkqMOGeCCCZRPXKygjI0gRX6
vdnbFPyPqmcoVg2O/Vn1YUri1RKlLYSP5KiSf8jbickf2Xcej9W79koMGfU17UwB
2oK+U0SnxJxejcSv92isno3Dwl+PiCA2Mmf3xNpwhNeDhB0H4HSq9bir8Ttssurs
0S0D8apdbiK3dq7qBQjW4zn/UeGYdWK2oTVeChtuxc6YKPREBFEZTr32ozmOZlFK
zKSNUiuu0dZ1atuKz7mWNeHSWOuPKMXSMGnCgIqIFeLk0320+iXrDKlm8RW28NDB
sGFO9JKY/fNpE1WSt0UtGZZnylddrdaRDPvpnoZRMuNLc1Po+N4jMz/pIpO4o7Sg
1iiaIV1irqGVt+9j94m0pCdTmejC+LrGbZ9R4Y1tdMsOW6hTyZ25b87edfkcztRL
KELM2ewWUjujUXTGT75Mu2fY+GZMuCjWACXyNNfQNfo/5rRhf0KLzd8VpruTKRNe
461IoOt5IOnb40GJvVRvF55COcbeNcMA/RQp/1JTtbrMo8+2QLZ+T0csHRYddvm6
NytmvKtiI2KetrwgTxDByqR1wMYGkItYr+lOhHgbNXATvdU6IriifLEyG693Q5Om
1IlUo+qXJtrRkPA7aHPWAYx0YTqf6wyZRCjJ7X0ltZ+AeSEyR+w5FHOmMqSYDJ33
MtL/jtpxwog39AfSuncA8NobtKOKzowzOoZ1GDWIU+IwWSGq/AhQ9gDGW0lNcnAb
z/HzxJixiLO5458EkUjALX+hiK5MIeT+t8ZrNET87vrfzTdNiWxGOpGvChMZ/F3Z
lwDDQuR/mLenu/BtnXHiLrIuDWEsGOv1npUNu9Pk+lEjRYU8up653rFU7ByCH1Y4
eLAraqBvx7heKGpSkIPmeRfX+gryrhfrbDJVg/7vNUOwerldVGN34zDEkU0MQH/x
nNSu8ZI5ShMmEYo1bU/T9A9jvesdY8yewlAhuorSqf5tm8Z30wPA0T7sMbJzzpXF
TatwB2qWTFpKP637czIt1LlOxa8/Ua3wFTxgCGW31cpFp9p9XmUqQNQvoZKHBYaS
fiym/fgdzNPrZJyCSW+KbZVzcx+kpvIfiVjLsuJ8TqoCRokNyl2fGOtAlZgtbxFO
veU9LYdSBo4U/W/dztzcpgZutaU5TNgTuy38djDUVeAhfq9G3REZE74NOBZgJHsJ
oD/6hK3rEVuEMp3vCWf3ooo/X34M1jsbfidnIpFBtKHlEmzaa3Ebnla0usM59mCi
xYjUwv3RJnLEZb3Ou2zMg4e4qEpG5qzGBF5Pty3TZP8U0jwvLmWHICQ9DvWd2jrm
kZiB+MT2R2/aupuo8BT7ex51skMCkWlauEZGTgUmS2iWce0pXjSSfEott+Z+ILQ5
CGzvgsaiwzpWyejxGI2HIbnwssmerbqOtYsUSKDgU2EZTCkcMhE/2gAIVpWvOAL5
NbbquSlBMDPqRFpFn/778evteUQgAEPRnQmJu2N8yc9nRP1eNGBB3aLJGSx76vN/
3TYIHctDfFCWSV+lSF4ci+lGMAawV8MOFLQWI4RmgY8HQCFtmIiqfEow9c7TXFoi
ybX2ORBqcTZjBZGfyf8btFXnj+Vfnx/kbrQU4KxzVNAxI1AaXRChDjgMcG+WtVug
tJa8q1tk2ZzqzZeFTA1kDAAeI2g48vq67pajRvL2EnnMCFqsclJeXKpNCc6Ew1Yb
dGIXNoKqnxZo9JJ5WB/tQnqaNyrIu2H5JQ/3TbLk2zixzsH1SydmpUP0JGEYYwra
o8o4+MlrBz+dB30eKFLKflLEod6dOnkxsYaIctLKtI/LBE38KEY+BPD3RIu5CanT
40LG1t+Sc3/xuq0L17+5jUpPjAr60xqEo9s2Esguks1bYwPKQ3HW1gfDuieBAs9O
+ttsSR6sFgRl2gLDVBrO4ZlI2iHkDlQ/U6nutSi6Mt3U8hrvvdSJuT7U5ihBOr9N
46jqXK8TxWjHlpdqP5b1MLThmjQuIWB5AfG2x0oQkbuN7p3LADQmo3vqXNL998iQ
MMYsyL5dzNfr1QsAxp+2vPeQz8IBfudHmvtVTeA9hWX5VSO5Z49eTg1K3Y4WxEi0
7c6RE1xNsQAoOxeRw0EZW2ksp5PTqBcvcZYxvtl+F4ORmyU1yPo9zj0PcreraMxi
yXZZlSdLu33KAh8qNxmZq4hH9rTfKwNtzQ7EfhSSvN7QcYSyM04GKVc4UMzwm+Ky
wi1VvkhX1u+ZagnZPSvlKgyg/6p4iObvhXX6Nofh8KRV9Gc4//4o6BFpvpgVYC2D
o5nWDb2SFMPjdV7mI3EYCQVbCieNQ/+u0UQSP6v8iDO53nHtmpgtbvOrEFD+JhGt
2qmgxK1+wigBxrZvJP803k5BIY2qgz5b/N0P3W0RB2a57ZIpKETcDOk7on4nP1cI
y8VxjeBXQCz8wmzKhTmfyHXmnnxDYff2NE874Pm0HWb+WGDdFg7oiYhElFDpmm8O
K59SAVr4KffuWdkhG1bzHKpjNoZGHTQ2x7txbSYG8OeP30oNPZJ8+5r1ndn4nhnm
YJ8Ji/73ypHrczMGQbdzPpALLPqE7qKp6+mOVqDp59Qb/GdC2EVjLt4tZz63RSJ+
PCT4nEAUALtCWGE7t3F9a9pHUxkkONQ6U6fvfX9QDjPHb+OYZdC8aWLW45WNiRH1
Gd3Kecq0c5qXJUT6ETokriqF5nJ2CQG8nhPI8vCRo4wsmqzc2zzsAytb1EOLvGKB
BGyBkHnDtDJZoCYtYxYNe2zUu8480rbKdBQA5MDK4PaCdOgn2CNdkGneEhy9pOQe
/QlxA/f8n0HKyYSyJdEt0PmzJr1EqxSVSkYvY+p/k2JhI0k/mQYwV8dy1Z2KUF2Y
4rKmdeLEbqkx5rLdtNTGTlxJxH64rBbw12lAqEVbeebko1X7dgii49rxNs0A12uj
yTh9FVngYFaslJ76dJlfz0SeVXm3l+aHwbjxnLTUuW/7FFSX1pEm0MFLZRZro/DC
BO9uOQC0DAKLPGp1aqmD25M6bsyUL6FOA+66eBJjq4t9zTJLs1uuM3LQkvWTNDp8
6KqpOjkGFwdJBem4H8mamlqVt933DbMMZa22jnD6N0LSkXe4iUttn+i7pSeriuKy
LqF2UbNLXt/sJ0DrBbA6uyDc19KaORxx+WoXSuTUwlOy2qbJFIr+WSzsFLmC+g7/
uEgWpTpm28qL8RQlsyxY0MDa24bPO0H6y2mASBKDowI5+8z58bG7xxf/BNFOd8jC
stPtP8Y8tLtmVRrDNcwa7qwl4vl7PZZoVrWNo6a42FDAiNVMHSeUVBB0xRRqStiS
SkMspzhyYezyv3J5chIovI/uln0qFtlhho3Bw/iUeI2HtIqas218ggJLISh6GuDN
sjI1F8+nPh+R/A0iCMj0WgI5pphgD5hLBiBFOoz+/y74/Z0J1LvR3LJ+oU781mfR
Hg0faKF+ZQ7Oy8/5U8NGBJLwnXfFB/QOaOiSXv9UV66n26bfYNORtLN6KbwW6Cgg
2eZt+eWkBLze8HL9tICCoCN9yGSS+yw7jq1f1P3eDHDaw/F29mbk9i4S/epHe1C2
VnHTaxBO1Xk2xeeSesJimkH6gJKJz90sG4ZfvM2Hfs2HPpWfcz7ZzpKyNvbMoTvc
MAq4GuqXyRFHizwpPavZ2oMrC2AvZR94UHI+Mhdpqxx+O4ornxbKXDTr/G5CqfgP
xUyE+jcqfhkDxvzdQazlaO6avqR1jhI0AiUi9UGjtJ+YRSrMUjwfCkxO/wg4kQ9D
2cZcfSNuF8srThqX+OkP9O3QLeyqhRZJvcFdhYOLcX49XPhxVmk2z7JnNqTLalc3
1TchapN31g9ZJ60J3pHYwJ03s7Trgri0DgbLBUsuxQyXoB/vzETMkSwixQZ/ukhi
oJjaoXduXGjikn5DchlTSM74X2OPzG5ZgQHW5BbWGQlc3yyiKydXKMTWL528JvQ0
N76nttSIuNWAPyD9bwb6a3SFJE5ZVr0hqzdGTLn/Ouhx5A7Bu2SHQAs1ZLYEI9ek
JpW2+wznfPv9ztE3F/4e4JVbACEjasIa/cKd7Ljjyn4FVQ9SGIOQO+4wbwCgjBUy
tVCQs9CsgK7LMR/E3Njjvk0rAcg9zs2625dqnzcIw4igl2q/Lwt6AqLv53vMOW7F
QKPYYVDkla9HEbOhC2SU3jT8wud7PSLc4rGpwzLBx5Kd87X8jddUis9TbkzDvl2v
wvmI0Y22n34ln1tthUsll3BJEaCNKtteyLuANGpZOQMt7JNc5jRDA5yoBEodic1b
54uBesH2OzWDA1kKcSnB0VzGXAMp1JX0lOmoZaCAOu8YXDUclQCoQ2G3UQg85rn2
/FUZ2dwczGzuxR89BcJwh6viaPWSf6KUs32AR7Qozhognsw2TlH5DPmckKd0Uc+y
HFYNNU1ovgPrmmueoW4Y2t4GKdWUfut4Kw8nE66Lr1Hsvg0jejaQphMZjc6O3wHp
xG0c7tnDXQkz8lQ6aaNoOy3Ctk6hybDiTknpgroskLMoivkClxiWJS5teNuDXg5T
LhaRaL6X0BYNzpKpHN7QFWoHvGipN+ii6hKDNblbbEs+r4ovinXAt8le+ReetWVR
aXXksI64qCKNKb6RhnS2ryk/CWl0ilFeqap3hOSCMG04WDBmdQu4AGoGb4wUe927
o1LHEWCW65mHJ7SAYUcQ1hwdg7zyJn8A4Z5Ey01bpfEqw/KyyLwAcOlmEriUwiyR
u4hVtGfPvWxAg7IsHPbBsAUWhscn4YfKDaSl0Hccx7jkRo7hMG1t5B9fv4cNCYXs
1HH5QuJJ/waiI2LM9psFGXUkxFUFNW51OraXjy/rcOsxZg5l+pHxoTm6V/dViiVY
NPxq3nnjl/Hr8v8UEGFbISdZZBCSs7bCqo7vFa4KD0Aq9neGryGXoL0DOr/7kRrt
njYd0tPtFLIuBzoqON1TxsJVlz3VfrfwgB2v+5V8M2iN7E2ymyGIzPPS7hkzOtOP
FAUHqKLz1JseyLrqARTlvaslGAPuuxKdEaR8onysyQ7llaUYHOAVeikldoMgWUNY
4FAGlDD0u6PmMTGvacCIgrbp04Ekh1AYg5JcXr92eShyGyO+vOzkWQSb7b5Pf37J
UUf+edMCeUp4/wAv03ifZ5GsDNwBVFwbOGGqsscksbbmL7VLwPFM3PAB7HHljgvX
ewq5wuyAIl29WaS4imK9z6ZPcLtCirn/HsF747pG55NgEqRwNP2Szpu7idwaX2wh
ZZD1TOOEt1yj3peIPJo6hEk7GzzVp9jiTc1BRao2gjiArJ0yafcqp0IzZ/lXB3pI
qzPv9jKlN27WfzjQ24zul9T7Hp45/V/jI1fsLoG7SX75V5nxIhWnxsoglazCkYR1
jjdR3nqWUv1OVLeSpJZt9JBHLUZBnLvKl/5uvoTHUcXxlFJkleTqVadOX90vF6F+
NIFR+2FuDxNg0ml0+H1Gs951SPHRTljY/RPI+1RPkv2SQ2buTlqRkWaiis586O5v
A7SvZwKF3oIR/HijjF7to+H2YP+mtMaEGlNlWNP+tnrBPzHImp4oPqLBEmxRPDqc
qoM3dGFQwL1OGaTZj0tQWQGx6qSA6qfCsa3vNRo2kmONKGUO2CQLJSbhcwJKQ5jJ
qs/IufKGnDyEVD2f+xX1BS3ot5+d1qpLOuUReFZG8voC91WTLLyAh0fGYN7Xy8Tv
ZIzcfcLHsfzrlqiPIZR/DrbETz4gcpBk4bOgFkoXUghlSiUIIXKMvJHFfc+uxF1t
m36D+WVh/kSO6wL0sCwiPeTNVp9eOCXzQYzNEetGNk//+Flbvye2isgZ/TyXaBCx
vuNifQMm0jAr1f7MqHUSqvjgGaSrLwty8zJa47sJklYiqMONa/LS1cjnf1OcibBG
fEX7duwiWHiH0Wr6tWl803u/BB191RBu/7lMfxvV7Cu2H0AB826JpU7Gu7yg0BQX
yrSKts9JIB4HnkO47aeJvDNyOBcRDnIJnNDhM1r2Y3chA6J7v/vqC71CO3DtnSjG
JMP7z+JrvGXND8aBhlDvny9UcGIp0kiizcXfKf9lCv1EB0IJDO0hMeIZmXOe+vuU
d6YMM5FHBb6QSl/yZVaBL9PCNYUeB1DNAvKi9sgXYA6+qbeBSD+0LWd59tNybH0y
KmNOMnr1oflbw1QHwJooxN6kJGGf3AQh3U1Y2iDBBRLSFRgOy3UaWiOS4Jf+m7o1
Rdqy1v27msm5StH+qGj2BpgDUBzlyTHFC6+bwF2EdYY9fd0f8moAbEIyXglm/dUF
vJl852Y7cPHQydRwmO3XYI29v3g1sOXIFIaDq6QQH9nS5DaOlWaesHN+WpH3cbiM
CSf7XVrcaURokT7LAU5Qnv6564Hj8JDeszvIROhSYgI/PzxGjPiUaWslZNr5BrQN
39zej97DcUHZFxaotT9wruyLdG8WPlgbE/GwtP4Nt+7YLv284LTHEpKyvBehsdFF
HIYf3CBnislfrm3HmTkkgZ9SEkjlGghdFBNn7P7nnoc4HK0Jd4DCnwvHnqu07K+d
mozHiZtXx+cLTCnmZbBwhySWwVKGbStGzKg54X8mK61qtlYWGpQH3AkS0PKwwYIy
UWjO2W7qnOBxCz/k0ZUOtL7vInR7n3+4/tyD1U9LSsnOcEpEYqCv+9amZvCZ1rCn
vZgzn3K+Az6CMy/7hx0iVfHtU9YnN/ajKeYMXHDAwUYBun1BDWgto4LZY33+3s7D
3NLhSqBfM5psTrlM1YQMydOPn6A5Gm5jM98cg05duuLK0GEC530IW/2UbNsEWeU8
nbmvX9q3eY6FARY4Gjyhj+WFs3sbHU6a0un/oNX8/X2y4GCfQB1f+w3NuQvwTfK7
/qR6qQTYMsyqyzjn9OYpc9CpKVj7YIP4xXOrbyPhStIDIqxXZKbdfLVlLmV6Rniv
EhabL2fDy0wJnCW++zGfVN/nSuI7dg9LuFIhG1z5mLOtBLN34FLm4WcrE5wc5PzN
mPdEEKYOkYIQ3I2L/LPbIUK8h0B/sOkgVZmcUfCSe1rKs6JmEjrxc5ZDhu2bvsm4
Rd53Ggqy35R3q9X/qujoBlZcZ4uUe6ui26geaAKX74CWBy1xeushxwbuyP30dy0B
kwF4SgFgLfMeWgZ6P1dTN+r1lMOCy8guDdhVAcjaGihiMK/ibp2zuR4AHncUBM9z
KigRU0JAc5+/eIMRgBmos/GJSnmN1Jv2Rv0Gt7gwJqHAb9Alhy4PX40v5ASkBh+F
CMDXA3uT/t5VvRJRZB1uKTwLdd+aNcPMfdyZAWBjgpJGEkHKcpyefnOJWgxTQHJ6
4NVpstMgnX2malOclvpk+0XgcurU3BnEwntnk3fca4hwdD6naSirtyW+KbT0Fb/t
2q3hon4cEOGlRd3ZSeGx/gUZg4gzrLZ0gvP327hyNnON49Pz1jxaXGwjenCCehZY
U6frJAFynF039x1IKnJsotuwJi8BWdKN/ehDBsC6YQvbjZPHs1idMjAxKroqKMpU
Yc3TN+uHyqmc2oI1BAuA/+fNmdV4EFaXe6yHt6ko+cSF3Uwwv3fclaH8IKY1TMwb
LRmsA9Le/JN9GFoldklEnacuOiiwDWK53QU42tc7JufnSPkhCsauDHD0zbnX3oCQ
BWxaUGF+XakQryUrp5fo8yTONXVfitDey6MJobdXcQKWHKN4dU/63HUtiJEWEVI+
FmvAlttNL/gjUgafYIEz2bJqy7EFjS5aDiL3FvNiHSbjoPRgUxwPUvS2c6XgEoBj
ooN/HDP4jrrsMR/S4suwCvm952lbsS9S4dZKK/FsaGn1y+1PwUQ9etiL89RDz8Yw
P0Yq7ps9vhTWpAHk25VvmV9XyyfFzxHZYZtNRp4ja+dijI/VUSyUuT5bgzj5qyes
nzvSyMfLCkz5m25MAOypcNyPK5HcPC71pKFDNzIQOvgxZ1O3EbL4KigTMx3IIy/e
wJtXS0N0q4oEEGxkBn6WbHVadXtgJxSOeUxNsiLNRGlbj6rcNWqnh99fMg7WML14
6BivPtVFk3KKuqYDXMLBnB0aaExbAnA0zAfTRQzfWE/gIqBHMX66dRmNVQA9w5HE
DlcLAQJ/j2MowuAk9nDyRm1EUzlMTMUTFkaxmcR7dCzy+6yPFlZ5YN9Uwmc1461Q
pzhAsi3Uk4HnQyX2vbk0AS2nWuMTXOqppr5I4wEEqnsZS7UBv81gQCMH90h8NU2E
mhd6GFvzr1nfydhVDzotyaOEgV5fIii5pqkqnJgRjZUUcVsTUFxtH2duP1qyhSLw
HOIltp42Ut9jGM5xHRyJRp/9O92hLW7ivrVPqvyGUjC82Cgml4qtZysBsfcDRxYY
Kd5Mh+xMwIIcELkl7LzDYjRnb8ek9NWg7pmp9+aWlByWyGCSHngTz1pt4BnP5FIn
CtjQ/01a9Uw79Z6PMTC5uqUlQPumkcRxmn5qPIXAh6sdt0CKIIYHLR8TDRQjzqPO
qrUu7s38/g2ghCUmS+1vfXWRqqxQA46HyahjTWa8c5pwIeOSguyfu/fL+huAslkp
al4CJpLDQ2I47EmjH4KMcVNay5PkVI2MH20v44oMJv+HdGP5wM2MTZ+7uwEqJ82n
V7lAJq15RfO+CAq0azc+DUMlX9bLtf6L1i3Q2mocarAWkN91s2oVMMSCT0pwZ7w5
QaTYLEP47yCyF8J+cEPPghDQKEgFI2notcswaqn6RCaDmaFXX334GUo5mr/arnJr
PPeQxbQgZE7WhNpRW+T2sEPeV7JFIneeJ2TlATilQvLto6MElleQqjOl0qIGI4lj
3LP+zij7/5ifEDku488oYoQXRBr/61cYDJVoY31g2gqQzUaqiz6GpjGZ9yHWqDX/
KtdpGbtCsDcEQNAF33BaJQ51lsHYMAwhuz7Pb8YM3E4EyD29WCPkAuXVNXeCFE2W
pjv/sPlHdOgoffOz/eEp/JrSQodQ6NjYHIXViJU1e0+OQOyDT/dkIAyIaahyJ0Bq
OM3DpMcFC5NwdYBpbKMDTVIkptNKhR9p/nzDknObss5/Mu4+vfeIfzvD53mDcfeo
D6hOAjdCJg7he96Di5EOOvQjyOpls6zv1zDCpGvcgzMD//sb81gBGOk/skVa3Cox
DpSQLaeDxRErnbnLrVmy+3D5EyH9QOBvaIjzab77jQROW5Z9Wr0EKBQ7u41QDQHr
hi0FS4IcGkI35Ion+i8t8PduU9RE2gzZxoWKBxHD+mn2zkAbDwp0V6ao7kTjDDkw
Sb5dHNIw/ouWFQQ51oARq3QWDET4KxCnZm+1g5yC3FhhsQQK5V31z+OAr0P6q856
WB8L9r5woeh0XhcPxruvsYEY0L4CL/gR5LfI4Jg/Xn9OHWE5xlX+9EBMT/vh1blL
FlcoPnBfxl7WgH0Ay5o+QZZz6uiWnPxyeR8Z2ROIVza1PVsD64PEXRtFO/YmI1iR
2BWQkHT6tbF613ZdiySHRZfHY7ZsITqtG5J0910LvlnjHPffmC4mjWaB1leRKk3T
bxzn65BfA1U7H6SMVauNHEymnNq6o1MLs46dXzGtgWgO82gbu2uOCCG8R3tefHiM
7A0PcUIKEKf/t0wXxx3N7ybXLm3asD7K2wK+MfN0hf/a8+aaq4RCFGpoFA4YugBh
54GFbuS+CvRdAyF6HueiDo2tMnrlapuD3V4zuC9SFn22inwbojgXgwL0ixayhnN+
hOvakjQOmY6vfq8fdNVJBk/F8JZXHpbWX+oHfmiIB+py7pQ/iE63YM6BXb32IoLz
F4t4yy2oWXFGcmWbvipiNYA3X47j2phiyBegZHYdu9aGRWcS0QVEQoGF3ERdOkUC
PzsgJu1Rb1CnoEyW7OzJTok0K7OZjzWq98i+VDf6zrFFsmBbfvpVKnWmj2P75D+5
Fn//wEYe2cj9171UerjDGlJe4Pg+Or/suX8Ej0jxJVzmVAArTrtqjTYFgDJ5qlR7
qYnCl7lgfOiJew30B7Vqq+VUFJ7tmxvTH5/FaOtl7J9zmqnG1qfTgOkQe8P4cILU
4V51qEAJF8IViPB5Y83Ta7lOT+VfvoEcqasVzGYUxezwvOM/Zztqfq18ISialNj8
E8gmky7yQbvvVtj8rv6UNdh08FUpkgG9aMOdK90sxvSTgCzVzkVDrX5Glmbg+cb4
gvZHQlMv54uExYtFPDejegzN9XvbmwZyQVZGaVxOV59QbWPWQ4FfdtgFZTjsEi35
mYQPivtxXqloNp5eJdlTEHFnKIUIzZuPGBrbNjux1ZPgTBNrlJxpk2A4KHNKpgi2
VBBC804xi23H1FuqHmblIIErpNp73FHMMCTb44mGWDjiKH4CSW5BrJF9Vj+Af8O2
/CTcixIfexGUzui46vjP8axgdDwAyaAgkjheAbNEHtoUO3g1V8FDXq4q2RoEO77T
ioRvaIOZ4bnHuasMjV4Cg2ad4UC7F1N7thd4UlQxTGeUMfBsRCPnECmMgSaIj6uJ
62Pdv8fNU0aSLbYYY8xqX8LVGvj86ZNTFOdiFBPjWtp637NfKwFk9Ya/oVsI+ZSL
AJH469WTmgkRj4iH6s6HjeSgXN86W1cdKpU5n8hfFLJAfBpNPktbAMKQnuBgsrSX
hL0yy946RwmAFukDP3Z1IzrZv+TepjxdC3JQJ8vBG12K8MISCUyyMRSocUjErlq2
iCcYFhlHBZ4BBjWIKTr8bYvA5skqPamsLusWyMlesgHWLRpizwHwq+AdWvnqQq0M
Qs7VjPBpe0BMlMO/aZlJ+Gs70AeFMKKct9GaCYV5SafydNy4uBrcegXNW5dIjdV1
XO2TAhBvYDnFWPUZssttOZQ997oZiFCRkLkVVAlAO78BwbqsB3tesgtrQ32LHvXS
DV68tqeuuPbruby/GezGUIu1AkHs0w9Pyhll7WAgX/wOmdNrECTNSD9Eg6ExsHch
8AJoE+j5gJoMAh/Ep/9S4KHPQQnYW+3puCWd6biG10CLNj5n2hP5oY2bPhapBQkj
+HtNPGVLrmchLnlFwZP92X3WIC0lPl75RxDGk+cLa3f7JXkmK2yhlLkkmyfr+AAv
HpPg8lpm5VT4VtOPzU1fp8bT1UIGltlyDc/2A+i+ImfWNJqDyUunEK36gOkzqBN3
G+PEDL5eIKjlEoJTFHS+gvoa4BFFn4EcLFxeaX7273+BUWDRocrIIn7LEz+3SmNh
X9+luPELqnSaBE5Nbwlbf78SsdwDzY/x/A6+Xysuj4TBiFNesLqsuDg9SGL2srSO
O5tgJbEegBJgSoMRNElkUYknkElJKqutWL0rZtfgPfh8gRfT2veA7vAgaj1K7hbA
+IbHMAaz5pUv2S6IvoQ+FdXYi4SQImMZyzWf2jUr3M9CcUzQAOLP+4vdz5oiFIQp
xrlCZuq+61Gcas3U/OMDlVmlsP5snvt4u6CeplkzLYfj8RgYPc5jz3ucl7xLiDkz
gsBEq4rG5VU3LhZIvcQ3IXbA7D3y73gJs3qIfBeqsl8ucZMLeWiRU3HEZIKd7Jw7
/aLeV0N/xYjA/iFtrJqPhGEvdLR0stl02tsLRAcCt+LgW6J4+0GlFR5b/aCMuyM6
bTs+TeNkI/K8BX3pGR9EU/N1NhKM3PPr61Xll65brnqwgA0yyKsz9AHyCLeOdVNk
2c6CPZMKLxwAuCoZqiwPMre8kEzd5SkMFcQdPUwMUnQpB4AeDOzh47UvrNZzkeIu
O80FKpvjA7Hi47sUuIUUC8CrLGB1h0x0Tx2ujNfzqjyo8VeFtDdLt8XFXQxuvW4E
9Q8OajDvFga4MF2cE710gTUpLfoZBQ980c9+/KV4ZHrnBOmia0kU+F+IxfT/ncOv
2qprvR92rKMJcOGa5irMW9NyM1BoSRAagYOLTJPXfQjCJ86FruUl6hFwXuzpWgpy
XoiDoCsLev82lw9hmemnHjF4Q63b7uGtk8QFawb60TgXrDRjPTc1biBmaQsPL7Yh
xhoqtOtZ6C2DM/9oO9tphsBgRXb2MvPwAnxEkLuRWV6ikcJyRxdXXvYPRd73P/9U
qLtA/ZrVLEN7IMv1OMZwALu1U8dr7+MRksMmc5LR/3uPL1iV6kz5hTPLGfnbmWEN
RlhHNThaE+Rr/448SwIc3C3vKp5yBDnS4wGJFl65QgMpXFBws0UTmt5Nf1mpPkiW
DwH78V0LPwnvAKrQuZYd0cOKo/UMCk1b+UspqXEnvVERehW9P2s0QB//a1Zqx6Oq
ysJY9OgwaBGEAUjK9mxSm7o4MYh6GcipSP4S7b7GZyBT3Yvdssm+D11d2kHpjPqB
15QCVaD71Kyt6/TkAnh5pZ3tyE1PPVlkW5qbrXpX3FTpM0tZdFaMS0mC2WAWf6yQ
EgMKCJtX+cI8YrIfovwVavfUr2obJJgVIkA+k3PBzoQe9C9BMmhB5AzErGeDJl6R
bNj9Y+MLCjXBQlvSwHYyGZvhPH3zhV4jDH7Hgt8CMk5lYNNHK25BAgUNlBCFfWzu
gyELurPL1hFXSwDU3AUpj0ekyfMVv6r7GN5AntAABkhDF0wOboI9oh9fS3P2gUyv
QbNrXmhuVIPUHSMgRoQuDQH8uM/kQlOUWZ5b2k/X9i9prP7kD8YvS7KiMofD1JSq
3/timWAuxRu/A3x8QgZFmYSl1wpHtYGa6u7k0iDgF9/Qj9srqPPPW66FsO2qHIyW
VpzJaoYTOlflldfowsc1UJHZcMpuk+/NlerVuSY4jwJGrkq70SK/X+Sbn51PKRT4
0QdO2ktQr4f+wakB5PRjXy4HC4y99y3jjTxxumlCx1bGd6CzexrH7FXBJXPuzyAE
DxLyIxaKkWBuq009gqJw8Op7iOBLmKl+uTRa5HlbdCEh76WY8FLfhOh0/9YCri+0
iRuPvUzpCIfIfL/A1fIKp57GqlDvnTR3iAaWky/x22km47ufKp7xmmyCnSbpjUSe
ZnXKS4OuWrYsyHuKpEiB32ChDFJaVWnYxCd5XFQUttwWbWKm3in7SonHuuHqbboT
fYdqH9teK78m8reHnfF2csQk/HNP5qcnRiCHJWoHEJjgkCQqfy1JH4G7iMFZa6zm
FdaHffLCpPCm6eRT2oXuHuoT2gIpjooKB1n4m5vVSD3HRoFkDkaXGCxBRyn+rXmg
pTjdRQoLUkNtxRqtZTMerCUJ4LHzkv3/IjjpMIY7hrV2/tjhwNiOjw1gRGalPLVa
uWQX+Qg4SjVeUGzNER9FBb7r9y5BK9HoqMAkPBxEMxID4mXdJqKW3oG4EdDnk1Dy
wYukQg9csDye1OdMIeFot/B+y52Ef7GTeUrdoQh+rmj/9MnIksxJSPEzV5Bcbg4/
/Q1i4fhEhFloz35aGFyxXp62a+n2gv7MzfOPZLOPYk66Gwnmu9MMjMYvsURlvJyd
vAkXn652JopfFQ9XC2/fmO5WoTjx8i5EP4RZvyKZyUyvHZQMvse3bCaS+Ft8Qpce
z5ZDC4/nV62nCx6fje+GTeGsV+/wXz7yM3cOleQ6dfqUlfdXEJWEj1rjg2S20NHe
hDwZKjzla9dkGs0+tEgRi/mewijUojylWYjjExvLCrHzuOcOO4RHaW+QoKxXYkGz
VBu03ykKDO6nO5jBzYvHTUeAdY9OVb/WPftoliBMpvyrCtTXVub5b8xT7GYsoBIF
xbOKkcMfC7hsMpmzBVuxr92WONv6pA+RclJgobzysk0l53yktZijAOMNmBAN87cY
93uiFZCAmaBF0o/K2nIbd6pv7FcSRh3STc4uj+MiLcjkF9FFq6+pHWQhaopdf8i+
8Cwii+YxUIh2n0dSupnkIqYRNixrK7UWFSDeS23mNphzby8JN+iVuz7cnUZKAaDl
4d0ES2V0cxtEG9h91u92CU7Y681GPF+vAlITjPx/s8j3w43oeeHxcZhaskykg7LX
Hd/YxqsiocgeD3ZBIZBj+lYgue8sIiFS3SAhUnrm/29J+tC6w9/sR/dwMKl46ifT
nGz8nB3Y8gJgFqgYK6kXkjg/wz1wyGDdXNzSFPKf+1hp6VXVOFDBYJuVeFKGKoNE
Ioz558XmlZenzEiygeWYg/Ud0lRABnLAGtI8x+Xt515diLoScY6nSX0V4v0KjYcC
nyWrEeqQ3mAonoKC6tBedVW42fyvPcWLU3v77hfsRG2p6PDo5jMwcUozOZzTBron
Hqzg+LA6X7qe72E4AbtP3JdtY/KtmJWeC7gBNWlFDrp40pmXkMFXvSnhu4xVAIN/
ilAOGT2PT6sik4j7OjDSqykOC9Nt4KsMCG5qxKQAmZD38l7DIyVqtaCqkXzf/kHg
W2RnvV0Dju5zrQEnem1XsV8+k7x3/Dmkg/ffYv9K2OavQlAog9uyO7FlftkK9RbN
cU9D6K549BwvOBCV30yo+udCUR3U4BuVLRNMeWxuXs/VO0qAzlA5gHe6wAzaFtL/
PBKotDqssuIQ7NDzVc5NOcuGyXpgZuWk6akBaVfPTtHt1x5grLoUMU3X7I7hewR7
NYgwlLzf6+F7wEt6bydp3SHnzbl5JEWhU+2cmr4Vh16ZUS+aycsl4iYQobvqTKNC
pM6ktIz7aO/eN+E4YO+JMmeOer7HEEIDB/CcQir2fN44fAkW6llnnMY3MIOZFHIV
hTtrRGOA+FmVFT5/xTX3yl+EVgPBIPfTWdQ2oxzbTK1auj0lQDmg9XjptJH/twGv
wMQF8ghp1t+BKF8EJ3tZjKjyy26nEJwd1MwdpSnufNpIjOGR+C/S3nNMy5sCeBFw
p4NDXhpNmrYIvwyd313IfE7hGunaVUNqwk15wn5l7+fHfifStOJrdQzrdf+INl3v
EobikGm5iMuJxN75pf0a+ioSJxgYcIQPhzkzUzEasSVaV+RNfw2jHpD1y/7jHBDl
fi6S7sDZTMctAaaPlj+Egq+nZDr//PwYgANZu1XM8HJDZxI41gY+9Am2dQSGL2ns
dQ8GOGgZABg/79wajFoHegW5BNjIFronP5bTRXNFMtCV1Zo0ThwLSqY3znLf4SyF
zg7BRRR4bFNPWrrUC3+EU26LgIgrz9XYMFxKK2utzuTP0QS2EZWrf5wbxW+3htde
3D07CerVrQP4lxfEruleUCzjl4cQBeDBLH6c7XZEi3W8ur7oYC9lLYQNiFAXFfSb
nT4FymjqzEQYV55VFAOXozVxnTelB1xBeOC3rMhM/GqzOkFFisShWRuZ4EtMcijg
cQQxdzF2+ULNw5w+KRLqUt5E08R2Ulz3KeKepF2l9dV1YvcEQ5x4Rf3vrZVsCABQ
fncdYinP5LN+6+VmHjZOguggYx4DRplNOMdGSPurvJN2J4s0sUWKrUmy+V/ivGBJ
pY2JitSP6y20aE1QVj1NEwSBbbic84YvC6ixDAMbD1SILdRrLxjLOeeGTnvJ96sV
vwqMeP8frMJYQTkWxT6UgehK4Bki7CbiBFPQTz7/WHutMkPa5ZneD7OjxUyi6lF/
FqRUaU6P/C4ih+EirDAfXMdDA7uPC4STOSS4Rq4+Fnto6lKgdeQ9sOXLKSjiSpQk
LTg4q4iWApHfveOOaaiLQRj+FX8lLnrp/QmBgD41jbC6jryXBbLV+dpLdiKgY+Ft
icpeA7e8AI7MVbfhl0rrgH4G1disgs+ehyy1AcwUXTY5cdPf39iEuqiGmYxdPEvX
7KvdhAjb67zyY6o3GNA3C1KPOeepNE4yZYtyXDRe5X7pUU/BCCD2mFAvJBGTJjzR
eQkzrMczKsHB4d7vZ17Bzxh04SKROlosdhqcwA5KXto0z3WbhbYQM6HOCQ2jaJ5H
0udA04ERdW6UB9ZYtmxQHhqxQ379WNXiM8UPCVqOQSL0j71A+XW6tLasU/pU/bY6
D+fqfosf0rgQlZpkLtFP6hiQceTOH+4uylsz2WEYuICNw9f/ndwGe5LENRkPlTai
Le6Axzi7sAuZXJ3U38XQzaON3o19UmzTzVCylEEgeQL92xxk/fb179jfx4pNakuN
85shg3+RnOaQ8U4gB2HBCHP8sVaOOXOeWpVEzQDQ8mWnSE1vm1p3G1VWgaKaJtLW
4Z7yCcN/JM+A0uNYx//vj0wEEibc2PwTWeGY1Z8z7GvfoyLLLzYz++1/0yJP+WZs
DRuYLh0SMm1JlZ+qsnUUVyMm/WlZqfhmMFdq0Ew/rvZ4zjkWwkES3sXwnpeSpCdz
TsWgXP54BqHQpZFOGi8UQQOxNFUTyYh7837sZQy3ShPTrrVN2mSeIDdVzGYNDd6x
RVMs6xCBajIB65bRa4u6po8aQIbHKLW7HN8lejSpghehSjRdAaDLyxTKDMW9mfMa
j4kBfvDfxtI3xdNvThaK/vliMo3fRk0HZuy/dExyX9GJeELBO5MEB81kCwlMd7Zx
HEzde6Ro72wMV7j6io2PobfrCUKS2aRj4VuLvBdyqNnlb6XVa236gFKguubMtqzW
bj0HojShW4devrRxZE9FiCeX1el04ifJ+nYwzNwMTAmHIqY+sX8iS2MhHXu8Y5n/
mlhSosAv43p71tBdjkPn1/sphFzbTDBqOLi1Ggd1klbGQEkRHv3joslXB+sHLIfD
2xUsBByb4yI+bfIp2BxkAOPfHgUkkBR6SwITaipILYgnFUM3fQCX3fpcWzleCw/J
wLCtUSawrp6XH0h4+RMS8yQuYScTrAiXtjG39LOzQJKbHBYDagfMV9QjYrPlWOv3
/V70+N4rX4ElIa/m2384EyT85+Elg8X/eWJL0dfPpeBtW9jJBxQuLICbStlYuC6w
mw9UTtyYZWGPBKUQoePGQjlCmywnM6xFhF9FkUiIkCpLVeZDjFewLFAYcFMFbpnD
oXc8S8r5bit0u+GnnJGkQgfGtAtS7g+NHDRKrr+LNPrppObkidBv7iIP6qKIO8yj
ajUQ4hC75YRxUHJPzRAaCZycICqDNmvW+bqAh8/wLijjJ7rBk6QivPqhg/XJaNUl
J9RWWEgCA4FF20a3JLas15plnzIRVJyJ+A15QdsIyCC6bBSkddpIuYJmwa/FGAyI
g9Mxn0SiM5rUYUxBF84EC9nHuXGN6qvXZBP1albT9DjfmeGEe6F/k0/aDT0ATMsq
uup57Yt9o9sFY68DY9hf/Vi5jOTJSfJPO2KHdY6BPFvUaKM80xZDDkcbsWlYYyya
ssvxy4JBnaN3QtBM4UqxpfXxGKq5B1rAwhbfoL2btJixxy4+uuseBTRyjqtfZ5DW
dswoBL0SBicgTIens0DdACEGpnGdmNRchUzXCS+juNHqXp18FVypD7Sfh0Di+Ww3
imcK2DHVVaosjNERGAOPzeJVEEvmyVZ/G+F21CxSRXns/diU2o1Bunarg5/9m+ol
Qt6YrWQlOr2WjNVF0VoQoH1FX+W4kWlNKLoL5X9Ld1/qKMaC9BzS+8mVRIKe3S9s
P464dYUyKrgpft/FnXnu+5vasXha/TQA9ZZ78do4fPOae+WgLeFSsiO/+JJL472A
F6vy8hGZeBEOA8e7tU7DZUTCYgMej1mwgG8/thU7WAtiSH9CQQChh8Hr1C95T8U7
cUYGlbdx4O1KmJQaVMZnPCQ/jvkXTpX2CbFTPqcfQfHyDeFIunnexMAGol8m1p0o
EAtBcAAbn/CCtJoq/ynCh0FnEeRot2h6lsx0jfTynj5JzRiJDwD47Dw3sg7bVAHf
BgPlgH9GmnMJN2FiCz2lE4KhOC2EpuPEJAzfMYJaEuovj1tznr4tpkiEsS7Ejwo/
wnLczaJQl4sWoG0aINP0JJolAxIE8PIIvAb0qSFV2DUXIe6QlRDC2ms3o2y0oass
vjS+1EvOxZB/iQClmNm6acR/Um4fi/WQ+b5UMGOjLN1qHRDsJS0X6+KAsCjcWXxP
8/nA/Jqu2bBfqKewoMNUB99GRKWAoN6Ujpp/TQYU/7pBlcn7OhFh6khJgIZ5Ut+B
tYwp8qNmkminMhsesdD1ICoE1JpUnimNl4fSIkrUdsPk7IGvZW04q9og8CpauTzg
GEAlCRnCv5NgkVayQ7Lo39xRPQ5hg2RitbOmVw/gxWAeGEyDal84/icxPoO+g0LQ
Zovlx+5nAkYYWlz4qZU/8CS7H6yWh4YiKODMtzJmY0ko3LuLKzSZ7wO0DImSWQ4t
8A9t0cfFoKcyuf0jgVrIBIqjk0erLFjVBG0DSbamiyTZSftocBVSRY4CODzD0CCz
SU4s1Vya+cH6AitTDilLpL5/efhoRb7/nculEBQ6tJCrGxxpgYFtNY0za1UHlT85
PvFxX0W6U8/OnQb618vYe8TP+SR42mTmicVSk1esWUZwGYCr0JjvJMiWK09WwX4s
6GLEU4aHsrnSn5if2k/5TTGtMw8GnP+GqyMKYrYzfAz3CDLgCUtD61Km8Kjqgdqh
Ff7VPE1Z2YNgvlhTH+Cy+g/P0kDMiCN67sh9q6udgpkaVjqBqQbajdIepHNXpMs8
d7ghgLYekBDlHJlcKttcDAwFRjDFYT+yIeh1xjB3e+Vf3EPjJU0vE5gkwVquM478
JaJgtg5NmVN/YW5jW4DdYSBymXJ5atBZVWaDn+5s0RTrXPFIi3ePMbkA8bcCXjK6
wSnXWsuk9fgmAOGa8PEFK+5eAxiOcAkIhiEoq//3Pv7P8H7xxNbUuYM8PQqDoNL1
q27SOEM+o8/YeFHcdooog4t72MpywCh4qM0MKfHqHpP5fbK+FQ0519TTwnj1RZ0b
f7euKIHOa5DnFSM0vklFo3bb3CsgclUU2i1UTx3UyVMmq2t4OPOEQ83xTfJl0NZU
EVgObx+t0tEcEdCXVwjNa7W0T87MuwontYiB7NHniZYTH4myKHLZtxBn6bTTnarw
c4S0V27qSWn/yiWYpcrnxY1zkAchemyI6tMDnln9ySEY1TMoM4bppMTG+HAfRY+v
byEVVMulX+DF4XA5WJJQXLDFsOkl9NV+EM4MLy4V/B9Y+p8pcLAK9gigm9fZ8Bh8
Z6aG0Sy+SvlPdWwQBy+mvlu17/3UYvV7msfqOi9XWU1IIGpxP1cGfZ31pR7PAS2l
u/Ig2fBKqFpKeq1F0/iiFzgjIUmvSKTyKZ5BtmJFwEEpEoNX+hOR5DDqVS27qvj4
bDSu7hCUSORSM98qktojEvTNUvjj2Sw9ghkJXkUX7OL4qaBRqPdfCDRnEDH5EG3w
kQ8brNO2Mnyh28E+Fja/J2nRBFWUb4hY9nA4q1gki5o/ffRy71nzwFl22zV0qi8P
uDUlTwXf19l3iIR2XRnGcivRuixr3Nxs8InIfLtsoIQhYwy4HU9DyTVobpqi6iB1
ZBj3YPZ2NNSG28u72Hnojf/V4h/Bvm/77FMOGelnZ1eL0xyVSm3TM3yY9LIg+Hwb
Uv3Or7l5ywtEZ6/6Nc+Gv+CXCS92b+GJNMDclKGL9yzQdeHnKgMypRPNWRK91mtD
HkFIRLDu31zejYQYJTBXy9WANPXh6UtGeuQe9Y93jBrXj59iZfIViI0YBhoX5C/L
idsYwXvFfw5OJuGvlQXRBgf9rOdeIk5dNavsbA983f42Ooyw4TjkeDlqePqR6S1P
Tl7DkxXgeOf/7L9fCogz/Okl9faWNsMjjhXJ/X6RCeK0s81MiqsYVsuoX9dYF/PP
2qOMbKBZmKLoqc/mZNxIrxmWHQwN/ajpEK1ePw0firl5TfhN88KTI3XharKvRD6u
A8+GWIx9qC6fL9JSVgfe/uYM0AnSrMZp4yj6aRqnv9LfJbKGJmlwxL5ssfM7JriD
eAnrLp5QzrHAgmUanJRfZ/Jvc0/X9bYzfJHoI0S2z5y9BJrBa8DcIETYLxK59S52
GRRjo2d+Bt74mFFLMyjAkaAfEgRB50jloSguVGEGRli0GZZO9hyK6kQlKxE56+M/
/psAyxoHVKk2sJBiNy36CNlbPlaj/nSAzs+hinJhZfaLFq3JbIzTiLjvkmpwcGf4
cwUBgsLnPk8Ayk05BzdI8Zi+RyaS1KzYkx46J66bPossvIfWWJ2LtS3j+lpyd6Q+
xP6wrqE6dechpYyPt/D4ZB/s9atrQEVk1XWKn1Z+iTY2iGtRgici5U77vJ7zK63h
UUg7OySoHYp5xnjzKAPEcbeLEjDdBMdTEZTYshO+wFOYR5z1ONuE98kCRdWVNDyw
fAJWMxk7u46Kkf43wSsOAfdyOGSWE9OF9VJeTduPkvOVvVdVFJKTIjNmGGH+Hze1
yaq6/025IaA5vbdl86cqAndTYQSpTbwVCiAKMZrp+eVKC9XYWeaS0Gkmet7X5tlz
LD+0O0MAZFqM7vdzTrF/jpx3O7frGzln67FrAMW/5QtFnB11AVeIxHdDrizKBP34
9ZsVe3sUeS7fGNHuP2d0Y+Rd+WAsydXd8ql/MtaWCsM5+Hapk64mS2J+KPfh8/oi
HfQ2UWTHebRThB2SILur6fApbEe5jd5xrRYg/+hvCWHpOhSbzoJM8SEt/TC/wGO/
SkVJN0NAF/zfTcY2FXwRF0W7CC3Oa8CMikRu/EuhmkvH4iu3zDdoWc0hS/9glvZx
tzGP/b6+DaZhVIby3HeRS8T0/6faXOCwMwoERjzCJ25oHVlorgRAPWmgMg6wW6Ld
YFi202FBmPYaCa7x0ZSRD76eKfoyVwIQLVMXo7Bzh7n6LElKDx5RN8h7zl2hc+d+
uEdTeJ8LCdJ32AOqB/9hdv82KLeiKwyZTYWLUUZv4NX5i8NJSblG3S3wvdTrTLTu
0eiqIfPx0BCEBQAkkimlDgBMi/k0B5nWiWqgUI19v9Dq1GNeupkak+CBEPTQmgpB
AwIMaFDgrn1HNl9YjAAYYDT44MhASuQz2B8EFOX1e8csSwreWqQDgQiYdspIqk5W
0Yibnuq1hADVjoAAkX5FC7pBfpfVv2KDZo7RwnPaDXn9hlr/ayBzxDj/+DNsO0H7
QiqX0hiUSWebDZdk3fgHPfikVF5kEyrTRsaGAk0d9TGdHQizrZqpRuZIbqA6FO5V
GN2gGzYroybc5ydRI1M0wEBThz+aWAkEwXb0KVMG5lvwcAfjSLpAIRECIQa6zlW+
GMGMZRVOuGeN2cHqbo81GBIGli8U+Qa+vSKnyKuCgW+u+ObRgSW1REPEWY4iQmVa
6a3RrXZw5vFWfaID8azrAQUti55ytBbIWvKqgkqEDbve7t11j+rCGUyD7SZj7EVQ
FirCRQYx+ILAn+J5lqLke1bG9Psib1F2lhHBh065Epu3mwAKkWwiwoin57paiNQ5
iTqlExoMgy7qcmwW1NYeR4AtD7T9Wf01tzMhfTH5GqJR2tYMeZBo+Z9FHR1XvWwm
9ZhS4ivaG3h2OrlOajDkY6aPrL28dBns/VaCAGIL3A5rIpUD3OdgEOhj3IiOZwzm
Iv4zk4lotDDlJouTt+synurlozY/ujfT2kGF0379RghRl9fjXrzRdpaeIsZurZqb
X6wKH/4qv6qy+ywmN8XvlMzNzk9U6FIWFYklzyIwNPt+tPy8/559a9x+Hr85z2a5
D+ekAas+GGtfHEgij95KrfsypbaMQMEAuy4B+GTg6GdYnG8vD/Z6NXKvbG+J0724
EDSJOC7KcesNjk5Xk8me1nD5jdW7OMEjJqGziYev6Gy1roH1C13y8iLgAooRJqK/
8ZJwdSIw5+qrGo8ivaNhtN7kavLrcvdO3y9eOA76mW0kZwgTQBcyLbaEcBTsqRoN
QEcfe0SYW+MucHIfPtNWHv1yJN0FI+PhCYahBmLmQ3Wugc/3IIJWfGI97ycGXHEu
gT4ItJaOMmRVt5hxxS+n9pCPW9D/PgCXOFht/VC8OlzBC0YXvYOCp0hbO308jf5Y
KKHCK/5a4EZnEb2OxlTRnCuoY8DYa3JZsCUI7lcdhogUxnWHcWzR+MaN6waWEjJe
w+W0d7WMkyiHA/h3X+R+vyXoZW73APW+3EzYOsxbVm8Ps5SrO9OZ1zxe6Ld/h3gP
Fa+JLLvY1wzVqBVzEuGrEQybffc5B4Cb5khKUw4h4UK+QfdUURX5EC1ScfrGEkxW
RcV4WVgE1A5BhcBZZFNeQRm1xXs0Sv44qu36WfpaoqV+2X+wPMhagvqm9rnpoZwn
zqhGnVaLDqxHzoMEY7UownVFTDieuCxXTssOtEtfrUSys093ZiYriSKke1Re7NhD
qbG4Hg3dWe/fQdoo51xpsy+VMrubccrUzXze9s6+DxwU+/u4hHkN6LbNrhm9xgaK
T5T0jXgWqoZkAI8o5szenaF3FzWPMqP/esQwfds7qrkqpIjWGupSKD5ItxhvIAnO
CYBtXUltMzfdBzFh2v9MzUKLARY6XsVli6SeccMIrEhqAuFQUdL6MEr1XSarNPqI
uh4vkt7LEEao9qqhIof2pKmPsU1Z9RJkvVqWSr9XluoGtpni4RamYcnhwhobGTT5
BxdyRCqswYEgIxxXl1NSrUwFTHpaLt+DDEpC1cWY/X/PoPuB1y9cpLmC0NdaNHyq
hGYhwfJF03oq+LJY+L6swox59JXQtpRIjRIaOlGCkLHbfHYmQsLkf31gMHb4zKju
BKhMTLUWgwCv1BzNXfjjc+qk0bhIKnNEynq/qbEn0shB0AXWetsWdI7cpQyjHCoR
4FK1/R3BoBUwRCPnBgHlCEFXx30Vd1sWGvbv5WH4vEQsKIn9J1zUV3PnYDvkNoSO
9lvboKUhDg/o1/mxY69gHH1sK9IS/1kQNF6N3hOKM+HTuei7RUJDDApxQfIzC86l
PC+Y7+u7qUSdV2MCPEbHpYPuE9jPchPBrlL1MhZK1HVI9bujGcZ3XrlgyaDk48Ai
Chnu9LBBRJCZXi0dwCGUOm+nIFFG6Y01OCLoasQAOTqHE+orvbYB2aRD6f5IsjG9
ox2sIeNeZ0JstvdPZPPSfTqUe7EYkg9lrd+Dr5R1LvVwh2Q4Fh+fPKew/Ic43twv
6LCI+TSOy+pkNla6dY5N9WciVpAT7+sr5pn3U4loBfrLSpy+kmmPts+ojMnujPWX
ncaybF84i+apQwwyDG5uB/v7hoM/l89Kpo69AZfp1lx/FpzfZ1vpY35OEgeqyMNq
i9Q4v+t6+pu3OY2svKbUJZaXCuEdL+2Di9FlWAFKJChaet+C+2TdmjNnSJm3Az/6
+TlkOXx/JehSLSpVBCFyL+AurxFhi3nYODDd+xeagJJAIFooZIILZ0dZWpdkKkHC
ZI09ZQ0lrzjlRiXYJPi32wl2Fp4nqfn/3T+JN0Tusuw2KQ8bf3n6ubm3VfC5cCVV
hnCFfZVXLBgW9eh+i6STpDK/1rdv3kkV/CC1d2Gca8jmLNMT/mkbaw9lKZY9IiVN
eKyfFSygQ/7g7Y+3Hr8b9oFaQRWWXzUS7ec/rBsN3UbEppL87hUE98P65Z4zWpGk
JkftP1tJT60Grr/LuGehtsdew5msq2/jjDsByMNJIjyCFiP1iywitBdqA3dOIUk+
TRYvNdBou76/zy8G+36Mu+FmBeKHuObH9A2dbDitYkBoXbU2ChQS2VwDo8gUXHHs
ln5ZrUxmttIJ6YQ2iS9BzlnSEIewzT3m6YxUzEE/vGxWNoKYmQSqoqOkWp5iHHke
hI1us3a44Dbsj601Mo2vOsFxu2OAuyF5Nj6Zl3kjoCwHad0VUI+Huk0nyzQa+9bS
8Ynoic8kXWLC073Iqpdl5MPLl24eLUNVHIgwdqZOb5jJU31ocgvARf8GgBCqkxIt
G5GoskfHo6d5M3alSCvIWWHY30pG573M74EAATGkjurvjkLTsVnDL91nEJcBb8tQ
4WLEzjeZXuqNa5VJ1Mf+GrVTfBXzpXNYO/pVMmGl7tAC9DCh6eSCNaitvZ5clmZP
gsiQ/ZaVXMJtR8ppBKzZhhRx/1l4/AteF8CVB57OveLA/SWodzJ5dOXGBaIMjj27
Qhkfd/QkLsviAGMUuFI6wKOlYxOfKtyAKL3eEMrzB1VIHItfU9bdB+7ToId5bbEh
5/RgUlk4HQhh0Ts+9TGte3Dw79KhvhfWhaDEC3TmBVgrRpZWBTwhyBI55Y1MCsL5
Cwh29q+orP5s/yy9wOeUG3rJ8KcqNnp4bDJihcgjqLQCBbhxpdgMYD2Rit7dnc6l
6MXeKblRsrU1T92QFZ42/Jol5RtPEM8Ipc2vZDc8ohNvcyPoWrcHgTbovn4sBwZq
J8H/PIlxwqD9njWjaaNwtnajOJIlz1YCDEIAWtAfIAEOzroe+3InmMXdhv1Ricfy
5vjbD3XHcV0OCDyakY433BZREAdU+nME5kDGvIfKOJC0dqJ1P815ddfXo62C7V7F
GWsFqjLeErzWNhs0pMzM/WlDlU09qDi8GL8Pg3a68HJhNtAL2Enn9P0oy47b5pat
pNwUINUemTlRTGUCuoeZcSLBj/JFCzKyUV6tbTBVA2uLFfV77A6gc/b/2XUF2XEK
bvygGHw8hbC1brwxoAkq3lhZLnOd+mCZPIf+Es9BvthK0RI/GoNaVLmWLYXbjlZ+
1PmmjPtWLCx9GwoNJ4OOmp4OD9R6je2+Uy7GXoSByxZuW7aNcMx5S9M8pvxAxS/6
FBaVlk45suA4XIojai7v5ScHVf2b70bMjPC9qy3sTdu/jVrGXIcx9Ue+/bLb6nrM
GSNg5Jrlgrz9RnU0ufY0a8btdEGnxLhBx0kfrobHStIIz506Xi1EPA8SHBA3cz6D
APSSShgpH7jfoWDzSaLpXtSZ5+FiHrZ6rd0TMrv8FXUMDHpDMgfbKLXy0qhVEEH+
mAoIiEnEecssISm+2a8a0b7kLi5LNj4P6byDcZyTPuBTL/uzenyPrgbawWciV4U9
ek23Ty0CIROZTjp1VTFl6QRrmsaDAbxp5wzJMxPwIoUvOD2yYWXXxz6F74lvVRPT
cYBIqAD0KdtaoP/Pk6K4vRypWwUn8kJsg7irUTWWB1ZTzXU4XbKLkJsieKxcRQcA
bmqxHB2LH9Fzj1rzGCoV4z2JVeXxInMcuFVp1Jjb0BLZbK6PNNClpU4xHtzZNZwA
NcSotI+7QN4zmPCKTZv5kZpQ4B05kkvgrvAFZMoBW83PYKQ5J09v8wMZEXuGopt3
YUYbs23xuDl/3Nycv7xOBTowawXmSBDmhxNLMTmz6M3W87T+dp+XWUKwkMStTzDa
S3XajsZGqNFQEBGcYvf4A4x62WyCf2XPAYy4iGdDO4nlfbOIb2JwbfJBYoY21a60
tOITyXvHuO2hwKIGt/LLkRmsmdYkxWxjdprKpdI/4O+I6rrJauwIlHlgjfLwJl0U
1S2TBk1AooHbLUMh+8l7+Ej/78dhve7xebS2hgXZIQlcGIZZ7ss5Szua+kT/lxGQ
R2WBMC+L7HBuuYOCN1cAq1JELJ08UXDCML2GX0RrSbKNMCX5tPUSX9EHLpJ+wACi
9m9iL4HKbmucDdb+MLGsrTOXKiwMQJw/F/LAPxfGx1ImrNIQFLDZRQ3wLRzPy81j
LeuI8XoOVzNR1hWVopGVK9Akp8au1fl+1Nh3n4Kif4jpGozSvfy+G6V14oDicBnj
Sw8L47tZSfGBY2igbUc4snZR3Qe1i2kUApoLl0rdwYbR9/hwFXTv6WM/xN8tIs8m
2J6yT1AxJ0NwNdDUuMJGUck174C+hHphgifeiW0POox2Jq/r5nPVSNS7vx3x4X1N
DaLpdU/RsmmhQZ10n/voRlusj+XI2tQnALkGKUFGOBmJIYgSlAGciQJFHSANzWfB
tEU+zgpsdaZo2EdwScvE7QnQe2wvA/famLP9Pa5dPf/IetiISBzWOx3Oqk3j7nkv
MNXMSHTgFBjWWregzWrpPqfCZkdzvCJgau71YL72r7SHKKt+qdrdErk2fP6W5C5z
hnYTmSskEbqWMPp2jO2BYpIogY8BzNH2Uqt/6KETC9AXbveKVNlsQ8EXKciLrwdB
PU7MTL2n1l8sfRFC0jRyoG+GI6cz8B8FnQ/I9mMGOcj9JrKkTmLbK2+QefwpCze4
S2revRcDp+g68OOZKaDoR3QJ2FxGq0PBtr1r1sswLMI5+6Aom63v4NQ0DRDo12Cz
yzC84q4LGB0ULMHoFTdnZCCLdE3bKsxSQ7QFJve6bDhwuWE8hL+sTz7Z2yEqublw
peD2Saz8Cy36escw+tzeD7vGu0cjKqrzLWSgl4IlCX2JnGgsFME5gi+OV3YyEaNX
r54a/wwFi+AnFq5HgRqIby4wHeb7QfFjxBPdJz/mNZjEJhu1WZaztnYiatdrzxjM
83/1Wt1h3jsqUSRYCjLgX5wASpRBue/upmm7vFNhJoEfDKZb9zk+rnQ6Gv7YmBh6
ElXJyftHdILdNFoAjY1/bQ7NoV6u8W8NDIzMjLPybDIH/n9LlBzNLmW/PO8p+Dqk
oYCHON8YKnanfSiEWO+5Jfh+JV4Qln5Naxpd1KfAFxvpoiWwF2qb9qg5QVNxQkxO
K75V3o5PkXjg1TmKf2QjR76rZkcNaiEltrrcmSaL8BU+MCFNX+OpSKh8yLtfzTF3
WjwGZE+2uZ07icgmoZkmm4gOxUpDER7TlR5Bf09J4HOBbYfCQZ+ROkhYjnEZYAEM
SZ4G2mU95/1XdME2sol2/zsNb3S4NLesw4q6pwfbKmsdoqcjd1TjXaD4Kr1oAYLp
SeWlT2Rut4H9fPyNN+2JCqN2NsW579i3XpS3ahoxLm9hqGkVL5kJ2qqqgJZfXuJM
4Cf0iNYrIpRMU3t1JGUCVGWz7crNiDV/ny8N9CGE7mAcvLZ5H0inXh6Bij1nZ44n
uuXVCzulls2KJAT5WDQfPb1/QUipv3Z1cwTQuqhgaHLn08vXYFNx5xoLzH+7hnsM
ZjTKz+swX3ZfjbacSb8rZSpn7xjkq2ryT7oI3+CH6VrunzD/mD98gUHGnFh/iUcb
dw6x2u1b3sNl52xel9CniutrCQwAvwXsbCv8U0f6Pjdn97As/WRuD2VyCVS5yvVF
Sg77n/b0Rh19RSJppbsP8O6C2GVRdGMck5TGI3Ap4tQV5Yk6Ni6LfDOWmxfk2Rtr
VNtiLOXUQ5P3pBEhXKsmGs/R0oi5B9MhvMmSeOp8Ace9xnQrgBQxRnR0QRgXPwmG
+31omba8b7ySYQ1w1rpxvZEIbSx04+If1BiWmX5whrXrvdmUjnXRZUokJJ0Zjfi5
JI4hejIq0be4UQ5LhVHCaAxUhhnM4xjuI+palfGTIU4QViqL6oAz2eMsJBbAaOSg
oHN+EXPKApvxy9rrcfZAnUsNoILlcvKoU8sICwRh5T1SWIaDZbQBdcH8dHGYlk0e
08Ql0pvMUGsI4h0mgV+8nSkjVdSRZzHQ0Boecqtyy46KU4IK7uGKb0DSDSaLvFIG
YdBv1dQ6m7B/951ltadkJeFHvxVQXLr+pEshAA26CdxSnpDp2qfUGqSBj1nfAjbf
z1t3ZSqnLosS/0v83v1fCVSOY6RDplONlBmH1B0+QTwKYmxEKrKEvVs6LvXIWxso
/4Fon06JzJzbJa6MgZE9ZyopJW9tMEk5pMlpjaCCnE9kVeVWBMtF3/8HKU36YyyP
J6GsMk46Cjsu770gLz2lBLND/c32CdX1M68rmp/X3+ohX7hMlUdywe2ZSWynJ1Sh
0pghuYgSHlivJ9AYG1MjG0XPTg0m2aDSrpXtY9R1N+y6+PcUB/jv4OcXHAM8uFNx
Y4opVRYhu2ztMMcGS+aHcJ6vvluBhu7QjA9OI1pDJ4zxxawfsZLTehl5WG45OETe
FIkbYXJdfLysdUAJAUpDrsgJ1FfIb/fIc3LqurTHAlamqPqaXaQIYDMAbvETgRs1
fT3W38VNoT4PUycB6oOO2UEUPvO+OqT0OyHhlvts/XnQZIJWAxksDt/4lTJ4MeQd
xCLy/5OKZRvAaUZCRNtIEEZkVH3xLU6Mrfu1cYRgrb9oEm35YxAagTXL4rQEWVlY
4RnwF1cMUkuFUYfD0at7hko0nbUHluK0EGr+LNMc64Vy2fY+4lfX33XOvO5xDgcF
ZbRpYmu96iUUbNOytfxEzLFuC+idHkO9r06DCKhAk7yKnppkGzy83nbnsZypj3dL
9rqtOXOEPdEePDYJCyLxerA87xj++iY26L2D8vBeg0y5KX1fBuQ6sNo99OSToHFb
V2FGDDGo33b1Z4bhDNPYk0//bYxeo7t/RsA523a7Hp5OrBLEHvrTAmRUzV7s9Dku
o0e9c8ty3zzi/FKEj/bBJYcVgpcKtN+f418biO0rnxgv6i2hLoyIBk7BSWL1c0Oj
3VbdP5YiSJjMp7AQwxuGr1zXfdHroEQzvwfNLhN+kbRwYd/lHFcTkL/qp8AEhAVc
nuOw5CltnDAJs4VeB7FSUNNFhD0p6rWZ3z9eK74LN5VO4f8a8Eg3DqjHirOXbO1a
2jpt21Cfsqs6Qaf6AVH5UpZ5nyP7CW4D/nyuSHaTuj2ODNosJIMscgvIb9xvxR8j
Z4jsVkfSHt4vH+FHgHDNuwcfiBKSX0LMe6MmIMe/7elmuY1qj+mE9M16h0cifnnZ
+Shm8lf3cEsErQGdURq/vN+lRSNoEfoc+lQRSx7ux4r9FpyInhpqgizBtBIeaUPo
M51t6in1Wod2pKToGzn9PgNE0iFRsaTc2mTAUxi3iGJmpw7JOphEmzeyKczolRP1
F7exoFVE7b4P0zBYfgG33KlouPAGJxBwWCMNLQfHWTPV9W+7RJIWyHa7PtqyoMT4
4urXW4yE7/Da7oBmMDC5y4W5ZTx+9dL1LBefaJUxa6707r+n9yrprx3e/H3Krj0n
B1GA9hexOedj1MRXinh3doAzxyaXMzV+FbmKONKUHIk+Cji6HVdXj+YPI2TQFlIR
O9ij0OQltZ2kkIN1hYn3VWihrInAvUArg/dITU7lxs0GrTzfuAjHTAhZ1aCeaPJB
Gwi2QjgMvgCDM83ehBdnosrsyGbIB/jpI4vJkEkVflBWQ5XCU4ghPcJyXF6PhT1f
nu6jsp6mxE3r5XMJ7saSvpwHqubGKWAEPhaieYPfYxx9v5doBTcz9DDG83+/CHGU
hn5s2YzxgGn1T/TRnPrf95ciYuOWvekUr6V8BV1RXUd+5OFYhBK68S2iwal6ISwc
2Zv9thcuYnDsqRPvltPHUFRm6nL8Xo80EtZ4t1u2YNYI4/2tJ/UZhMzfGlRwomhm
DQU1FbxeyZrena0WYofJFfYJ9nHyCLAIbMi8nlkd8v8jliPiv6t+4r8xeFKM1tQ8
xgZI3c7siUwie09yM9sxtEgJTaCT1JgVceCWG2DLTSEWtd/IxzFZcv8XmY7x0L3a
NPzMVcr5SJxhqkDodflINLTx8TcAqjFFN1Y8fKv6Qiw2BcpGwswp/6tgytndGWUQ
8/Vr+lKCWUPaTF3hnPL4dIJAdXmm7NBFAUkcl09riSv/HGWWYsJNMRUEnzfDBqNg
BDGrlE1hlmCHj24Xy1GYsDrM+HBIJaNyeNuEVo1WZcSV1mCpwnoYD90xXrRz5kNv
j7nyQ0LAyJoDEesirp5sJOKrH+O/jCJK3g+hwe24krpJqJe60XGNilxHJii5SDRf
Ct83N9LBOEGcXlf125BAc6IqW6OP9lCljN6rNXmEEOa2GOjop3p28sDsKjUePt4M
4UT7VLc+YG8W1WbDHX2T7rPG8/zQOoH0jCSSgGs6qtrPPHNVTNj046y6yLKjU/8q
DUiC7nIfPLrVxvyydX8cBBihFh25Dol0FOtfW6sn0yKRhx89fJmxjl/wXghbzrM9
wrW2CgTwA3PF4k53C9tMafp3I05oXiXGmlvL0ztggW0q4IZvWwunC596FIjqWcHr
4EYeTUAOFfeOEMcQZcqUSScwcpsmNNhJb2ehc9M0Ji2+nHTCXbVTcOavWOuo+aRG
37//LqpyC8/A/CvgT/35sQHveWO6DIrVA7iG8VlYcwryvsXjeN/JTNGPnTIOPHvT
Pfl0N/arEgXKobOhKe35jRrn4ssjd4W18soB7VQ6l3xuRY/tzS17hSSpHWpVPMv3
GURrUGuRBSAry4EmTy2pAYoc68rf69/OofkZA3NcvcuUxwUlm/OyUb0Ek4G37rwF
olSgBjrotWsDk4JnRxGVVit9Z1CpcFvm50s1+msKCgvVe9nuNowEkbrzaaUxzKJQ
dXZMY0Z9r9OHSYESgNS0XjeA9rQ0Ig2Az7DaNEF0xWAf6+LZqz3HIzXH4ZL2cd/l
aLbiUyy7/GmRSEp8b7dh+dpJpLKPNC5hVWHgkzDOyj8HRmhRpvLxurjnbN6+PzJu
k3YwiQJMXJZDy3o4vku721Umk97ujvozfea2V3M6h4XoecXBR0iWLCWbVLgVdyHH
e1cFPmjuqaAqARoA7nREtCb64x0WeaJVVISAreAwORjKXaBHdUbc4CAuyjHH6zXN
KhLwu2Z+ZIiXvqCS1Wa5aSMbaMHWr/6T0QAJgcpcIq2jjkyedpq2tdQZUwHF6uHJ
H2XjNP8YPMVGYeKK8AoE8UJwyUYxDo8T0sATYtwaWENFmlVxIjyZZ5HuM7CkZtaS
pjO/f+SFvdBlIJvs4Vsx/fJbugGmAl6ax4yyvrHTCJjIa8OcB5s0ZvolXZcgmmC7
C0TwynddjwjOmKGBbMLrbmUa7L47DA3Vx5fm34tiHYAUOeif/zANjzfBZCw5qauf
tCmpnh3DPOtHvU7kb35rYMzMR1iOPAOd3aJcSrlzOYZJh2cexfgeO579q5povWa5
sSoOcBx0YIyNfrTKnSG6Ykh3sqw4j5uqVMDTmZQgOHWR63wVw2QJ8/fiTtW4YwtZ
Wg+xnwrKN6q3W9h187KO+DHL540Kky8GHbQywj1TWLXJqvSRGzCwFro1v2wr4FD1
pR/y3NCWSseDgIaX5Pi27Mw6bxsYrx8HJyO/JghdAhIg9wJXecVK3XL/nPOZposL
FnXiEQZ6QCPWtk5RHlgPUr4UVVnTTDVcdk6rzwab8TM8cjs0EjefFl6pQ/x64T8w
MVQXEJHsxVDSi50Ns4TYNVqb/n08LsZqkG9sx1b9wArNy2CJfsHcJxffu1u35WXC
1vc4kegJkAqHxpcX2SzDkJrxQNAMpTODbv02N5F5JKclASFxMPhNVFNU9iI87xOY
JS1p+ze/pJmIFj5PAFWJClAL6ziHPZ1n5u24cEA+QrVvHsieZBVIzjpRyUnITtku
cijRdeSBRAdQs7EtbIinp84eMAJrdTSuWkQUM0ieGPES3HmoDLLcBo23ePSwssmh
EumImWacX9RFD8fMSQRaOZ9Hz9nTCZISCiqfj5skaBlh0aF0haW4ehQxYPEnI1dV
a/lEb4PlY2dBCFbUVrZn2qtaJwOobKgQDZ7FqsBPH75M6O9jlqkI97a++lkzveHs
zhGeahWEbV670zbZSEPFgwThj+gyZxomCxZdqGUmpsUpoYcOZlkF7hftP4f4v4Oe
BXDrzb2a4glhSkiabE7gOuGCQWsw0lCB6kkLggGrAvbi2IxGrq4stZcahMzuW6vR
7f7hL5rOfC6h8hZt4D1jXQWsjMFpb12o5x1c7PsRDPF6aQK/7mWX4DhwCEoUK6fg
gL4JIRv1LnCaw+WiCj9BjR/22HcVYSC7CTo3hiHm0evm25R7TtjbWPOrk7qN13uN
sCv64/W7JNE7lzmzcVjENpFtEgiaHYbN9xljWfHz5/1mie5WN/HyzbHm+sn8UboB
fehIHn+lCdkb3fBoWs3SvAIdKylJWWZLOkcndGDylTOkwCYr8Kefeu92gmRGkgVy
rVmoeiiOvc2rWOp+2fXSZx26Y3yvgMMTT8I2Bl2I9dvGpr4IwRd0lbwPTlNEiIao
8D6K0rxudjKBTETOUa9kky7q8OLdM0qNcOYHHWIPiduELDUMcEjXdGJ5H+aVNnAr
E0O+bgkRrGbptf5zQ3mWWaRXTgvHjm26VezuLIWyGanjbESNHucVZbluTCiyH/x8
Cl2LiiGm+MzMp1neq1E6lKlYiIMWA9IWB7i0dqFXpocu42WMa0C0ZrAqZ1ZRjybx
ge/ST3lHLA2cusTQOmBlUwuOQ9iaVGnBXgO7JLtjDia3mfrv0Jf4epRSy3RhP5RY
nTkHRz0Nfa022jrZKt5nzVlAHuxFUCbU9i6NiNLXhvtIkwp2icxLshCvzTFInOuV
w+TgcIYMquW0uR0Bq+mgnKEFkQhprJRbqQXR5tQPoffQHdhZG099hWhANMl59RyA
BKUZi1qrdUpIXpTsa4zTbL3QN86NrN9H1Vy9MDErZass1/E7jlHl53lhllOrd7ap
/Oatpq8sTJ2fiyw6dqvay9VdJwGYaKg2DBX4B00yhaSKbF4EyuS1Jfcjh8F4+uhv
gWJ7yow+dS6DqN0JrnbKcwdh5Fj6V03zGa+bgPbWIbo51WWrcUBhRAJnjJEUQmI8
EbeuBKvBZjX6sxTNaMrMiYygGev423BWi2t356Okx+jQyDPzW1qZxVLFCkot0il+
FUw1CR2CVzLLjBhooJb1eIfsFOMOF2Nl2iHfxLF9xg83+OqUtyHK74ui3g75Cadn
+Gew0Uo1X4NTAGwwMBI6xPrEj/67v3oRoM5jEPGpjSxEYE8re7KDh0ks0ZwEazUV
lQvLEcnznBb5H/huIjMghWXFKKl8D7VjUMqkicwijL+pQRbRdYkjdEchnWhQWESc
D25So7AqCrJUawpbUK8q5/Xw3/mAIXldhXY7QXG0Wy/suqvXtpDYa/EngLGLcQ4L
8GwJHQ8uCPj3UbVPQzrwIy63rvsEvpRYTPnUyh9/c3ac0Efq5E/MPkziu9/6UtX+
7DBa6KiFSIyAv0W1pZTw5YU4fm0medBKDV2MlB+M9XjUIRdERWyT5ZFRsW2BPXcZ
BHO8S2AM4+BESwlv2aWqHJTJP3JuMiDOb1qXYJI/MRPRBROQzj4krpwUVL2Ypx1u
FLa65PSODC+ggIPhfS3Q9D+GprPTuHsWk3/on4kybB0wngORM8cGdQHJegKIAjZx
Y3vNPCoCxHI/6U6uakZCOR+Jq9iitB6YHUwhTVhzIHivQSrP4yJrzDSdyNlwOjqQ
+KnduXAh6VuqsvhHgVRMZVIThra9QE524Ev9cvlphQJ5fqzPwE3ItB3pWtJpjyg/
afwLtMe6wO6jXd8C+mgSDHkX1LViUFTDbj1ShrlOT8XRT6jypLO/56oLqE26Qyk0
dLlzdVsIPBc+bksgPaLwGPrjApCGtQhOq1PY9HI0LF9FpTINmak3KE4Da1K5omBX
8TGuxa9MOY3O/xJPaBBunPoat2H/E/2spAEo1yQK4EiEomXXHsMC1eC83Mh9KNxF
Sb33qULEUIYgvTPEh+V4p3kTs8hrRfK6OFrIuU25OwSGhYQrp+bquYNoZ9vEZw92
yemEJiAPK2klA7FwpAJOJXGdA/sG6vPTYXpfpVC7AhJJ3/o+m+xze9j+VvvkjOt1
/KXU96DFGH1UlQFCGTh7ugY5ekPlsZ9+yq5T4MuMKcuRnE6bkhLtp+gfDFRtIk5e
RqCFsSJ+a59aoVpQB0GEtA7tDko6H/lom9isweBTGCNhgoC73RJu3DaLykNEaQDX
g7webLAxm3Uzpl/xM3TJNEr45Pm9b8BCgwi4PEzPDchOne0B6JwYVAFwWlMMFJIY
Kp2FFcYxvBPoGgy8RDpbUAwqLv6SDO2/b1pXd5LGoLpqY9ApWaf6aNpO5zOIJN7Z
ZlzKu1n2XrERk+qtBFljy7QSqd4xD3SKiVyeO7h0UZaej2S4eswAiuVZQDM1Nbqj
BlfgS/GODdSWPFPkH1T8OUX+BU+ufS2QvM38+v2hlUDJ/sn1ZKb+xWQV4vZOdJXX
/DneuLV8ClUAukDQ9Cp08xBqDVUzbq9MAoqk7+6ivBeTGq9lky4tEu5KhOeU01KU
/tmEFm3C08kjyyhgorW3a7n+cA/xejI9RbMsMrO2PnMMyHofcAwbt4fJMXL356sz
9SLlhOlYFSRhvwY08D1CAu8FWJU7KpsR+BdrLRThi22gSMxX6m07rrb9n1HBt6jQ
DzuFkrpZ3OFQwPwJ0fSspKuUxny1edrjA9GxFZNc7idh0NAuBURS0XEuyA7cHIef
K6oZrkb8o9QwcU8Rj9Q+5ePGUai/JkLRZAqWS+qep3+oPcmQrs1AfARNIsJ3GSLr
j5RdnlG7uNVALYcGIg4U79bLGB8Azm0/Gxn7T4n/ibr5qwSG3zhJM4wrcJ/Ureci
Ohqvt03fV4EnwDgj9eUNCah7hA9spb+eTqtHbdS6P+k9emRL0tcE00rwhoZRomEM
nusLeKqsc4aaUUd53cxVhubI99ufgT2Jr+eXl5YlIyb+7rw2LjihvjjfkYYa9hW3
U+PKeKfieOUMUVJVHDGjL9EiGxU7jqBuHJrodNhnS0pdXK9z66lJVUNoX5k3fQrn
jinoGe5n6NMCIIGNIQUqd3r8NAsM0V68GRm583Gwg34pEG1BPLsyxuozVDReAbrx
FN2skE6leowWnzYq5jcfhAVGA24Vkw0XAIj6Soj2Y0tM9l0Wo0dDxDVSCEpFvsxs
fTjanxZVrUuhyCqJctOHw5Xelnq3uUIwrhn6+nDPTn3g4D0RCIpw0acMMTLkczNx
om6KY+q4azz+O+Mn3hFQH682uyE/ihiCIh67krZxTndVFiYoqM0I8gYhNXduuXKn
y3uowmgW21FmKUdPOwLy7plKtSGT1ZXAQ731dCxIhj44x5uLZ3gBo9owjPBvRwS9
ZRrVUkN9E1Ik6XMNSP+SuWV0z/TrJA/54zpDptJZhtbYtVpDbR5HU6NTzYYKmwe1
8Zm6dMZ2Fvtsdy1d588iU+BHzMYj68Hr2s0s65ViCBl+yXdQR3wBjI9Go/Rrt9BP
kK6uJYtUwhs9+YXi3TQSykuNNRoQpCb/u3fZNYYWQI8Feh40VmMfpZJ8YnG8tCBD
B1ALu/OAiqRAlzlA+9OcUIeqQm7Ay6+NSFDoBPIq2E68Ab6NlLcvkrRDw2ZZTRmK
klYKSjNHYU5n8l/7v1w5e0N+08rnBvH/TITtq8ctV20VijPXFlhz7nrNH7R2mj4O
wBVH0+3AKHBJesSAGAC4is9GPPjQVKt8okXRXng9RpmIkKSdAu1sI6/YplacFir6
F0nL6YDkg28iZtwWvsc8W0k4L3T4JHOulXFQIb9/bYydJQMTSia0xQ1M4Zuji2X9
r42xUK2dXDYF0wIrHVc4PRuE0RYnUDyq1w65TaQkxtRxXaSYT+86QH9ko+HURVrl
YvmMMJpUoebDK2LLdXBRwkVw7eCVGW8bFcihzV4LthEB/sbRGBpnTRIBRk6l1dPy
AH2S16OIJzGBHt/we/4tuzRk9UnjxPG11NdYGSHalmhJ0iTfewpW2nZGj/4STePG
dZcF15ANOAk6qLf2odm/4lSj92DZih8HL+dCtTdt//CRdX7NDg2VAADg/guUfTeC
/H56E7u1I6hTRFRs2wx5Q56cvlNu509TWI+CjNJz7tlhSYpCM1cgl/U6cHOxTZDP
wc2JsCwWvmgp324I3KcsB9JbjVfd8aJ4wCsV2g+mLJCto4APCtklBUER2HhkpZ90
Lche012GMI4owR7uQrL02T1r8LL1ynaT/3vBnfaSY2qgslSfCmR6faLu5Jtsj92N
HIxrcxDGHEW3XlugPnJTFtP4P2SniL2mZs/AjNkPT2SJCIdfGXqsrXuoxqR5ICbG
rLcWGEMG64fq/XsBcCTearF9O2MTsUwCGy3yDjysjQuuuGGsfZPoQ2Q4Zkq26wZV
yqOR8a0m/OoQh+ZgRB4I1tB1xjMdWKvoXlpXrVuJCFPQWBIkNgbTy1p7D/c1fqXu
5CxsnGAkTFFuvWhBTmXY4NKajMKvqvd7u9CtJCe1KX/jEEuC3kU4a2ZDuHNBMkbM
LOlNz8SqP7iXLkxC0JsJyHTYOJ4kYQ1aomY/511NReuKi+CgY8/fW4efUXjHhHGs
essndmd5/3id/Swm0sufiDA+8qX+or5YPCvb9SG0A7D3z2Sdp4Pw4rxBwWaEWg0S
ssRzPsvQs9EZxsX/t/hdlH/72gt0G+GYJYRgm383Gmlygjd5iiRdYb91cZS64fj0
Uo+3GoYlFbNznoz/V1prCMPGoLzLQ6ulcX4DoFWpJYc8xBiNUG/WdfDXyWaHDBcT
3B6kvv6xjTzCzoD+0CjWOAkP8xxaJhCanWUXNZfnab9Qi4CYTlHaFe9hCD5IuwIo
wOPKWG69qJ5ri51Wl/Ock4pNvoZm8APn8038JpgWD/4LXP5ZaKTpP68mrKHuo5fy
GNFKSx5aiWS6Dl8squ3pABL1yUvVsBFr7H2Y3laNtXerpmaKAPv5yISNyOo4zxNv
I0Bl2ljsNnc3qQAaY5Qv7WRqOPkfyGjrw/MAcZLRQuCnd7fDAqvIFMxCy6V+gZM4
xXEiVRCCJqDiT5KkHdENiugwUIf7muAQ4s4Ozod0QPVZFFhOy2eCvztCilVwTiWZ
jeAbZXeDZ//ZqM6tUlPgMWBoke4rqEY2AVqyH8f3OlsaTvR7zDtyDJjiG8nuoylr
B5prMbwC+0KygJ3ymR4h4RdaKv5vPTagd1lX93HdG4bPVBwVR6rpzQRmOViNR69l
9QB3wnIeLpRv3/TEi2NuZZBbcgHxhBmnpKSJUleuufdQVkCnTrWbRSA36WPmpC+d
nBbvflDbslb+2FU1pjnl/Gj96MC9Lg5uRN65eZexTToazFgK5SfgcE4gz/kKfkX7
cFBecb0HsX5F5uNcJAcRakdzpC24lCnz3YHzLCvjKs3lxNHGkXCqYNzmNknkmvZT
StJnJ3BFeBP6sQM+HtKIFIyOioVN9Jj0kTuUIz9dFPkuB0We8OWAG2YWhS0Ub1zL
dCHRmu1Z0ihC8K2udv7SzMK6AwwjIzAgxHghq9NEk+ZaFo6Q5x4KpoquRpZlHqfC
E3fDjs26xBF+zrIxjBKpmwgY8YekL7/+sXHYwiED4pfWjc0FP4LvWLlkDiHzip/9
wSnZQgu22F4DnmLAAKz3rwQHPwKeaYkugZl4ze6DIkNqXA2z+4zYYebtQ+xFuxP6
rGoi7d/hATkFUpvEPPYCvozlFZ8NXXcKqM3y7XHJBM4pKOx/0YoyCSJbdtY8egz5
T3nV2pq6NPqu5FClom3EYD06EmdxeYTwIogb9miZlpZpUPFBrd8ItmzJM+yk5p2k
HkCsFxOIJJ4mGnXUs2+1y3GqYOW/1SsCBjONokapiYB5Ta0K8D1yYtS8F4LNKjq+
jsBOxeJvhTIuI62r0/Qp1ZSPVNjFOUUraZ763uI0OtmPKqVoWNxBKNmu+eS5DPka
eozwwSPujp7B2rLBBPoD7Bi6Rw0Gfr7isPucYh7qDxzoXCb4LZM7ln9CBB624lXv
lYvE/nAx+Vks2wgwHXTro85NdPg4gEk/7DUHa05lp9pfxIjZodK12avWKTLRcT1a
ftf9g+zvpO7k8RCRVinXc3JTAAU6nmhZ8u1+iHf+E1WEupmMal01aRfJfZxsyw9n
jgRbJTHd9AgS77x2tpWuUNflIeSudMe2U+JH7OU1VOixlNQSrfCrfcW3BsieO2bO
UUSQAUAiykxPfyKb7zOR7m2hk5Kx2Ipsbs4pGmEHSWtDhn6PqQ7HeEq+Kz5K5hOr
k+jkOHFsWOfayMpxMk6d9Pw9zzCV9/2OnDf3zRYT0U03aWB1nJkuQUM9sjbBXZV+
JQPKBUq27xIoV2q6ZJkRQE5cVDa46NuzXDYM+u8sszuOSS/rvf6LPVNsvsnxHqd/
ar+Poql/Y6fmwg6jX++BjcKOZf55QpxW0VSRgEVdjqJCz1OAQvEnRMNK19/2DT8d
iGDdX+8wpZFRUcLGKmJGW9X3cn1DePTrH77t63qP55PmHC6f0uFfRhj+8RJwZX5F
P1XizNoP8XBE1RHUQWxiJN7NV3MXhWQZYdHvmgTOZErQk1RRwyBJyVp/q/9aavs2
Lso4/LRVeWWjhseu4x3IoV6g4gP5LY5gGLxMCqJr6HOaZcKi+ZFRs+0L3Mp16h63
glbvFLFS2yYU0SROH/esyWULBsyxxEH96Lhgh8AaY7R+AFwXotg6HCH6rTBBNac2
ktNrHu7ehrYgBeCmkMOnFohkJAN2n5LH0Bf56kDKUSouTn0oDnplSlSwAtt5RtHW
2lU9EfPjVojwMOtY6TJHPEoyUicc64z9pBqsPF3uE/LbS5zieOZ1IULFxxu4Z/Cf
+9UbulZhccGO567UODAh1GaZnOTVJ+pZln5SlGJWroguoAsGI5qLWdbGPraJ2TLx
QnaqSIPna4Fg6b/JeSsukAuYnNlZP+KzYIHuFX/A2uU1UAcb9szs87j5L7Lo6s3u
0xoNcIVCdvZhHktNULInnol7K2tNFUpGnevmQ5Sf26OJBsdp0ZCgjGyzW9OTdzxG
Pj76ifsidO+q82aEjwlSJ7r4NEGjfsoKvy/4gwq6EXpiMCASJAhHqKXOhm6ubUQL
PqCEcGRF7tF9VjvCI1WnIEg6Kq7z41QR6IqSFo2sDnMm76djT1L0BgT9W74LV2ru
wO3vv3nbVjQkPOvPdDq26Ts7OeU7FgUcymmxEwoOxzDvICtI0FS/gEMpWGG/Qbxd
1h5jSR1wACRSSEaiv3AY8ojDtkwlg6SPn7ftvX6AmwvXu9DujKAp5ne7qFFisXHU
88uHSAlI/4qM1uhxIXy1VaCD/t0OrjFWyvjzmgUqzkJO8Swg/95y5ZHTciy0sDez
o7xDV6zC8n7DBQDiBtZ4TM7rLLmUIxfcsVaa+y4A/cv78G7hI0eNA4pYlHPzVsCD
wyg4Afpd6+3l0s6PrVHvACjRL7RfOW5UqurD5Mx8eDVezf5IbGsCC4OyqTcb6UNJ
IrES4cEiQSkpjwTa8p5ER1muj9WgmZVSvlJX65503E7Tn8xPucy21Ajx0PknyOXm
kCXlHQ+vP54wRZTkjN74O/hC+S2KbxQRVLhDski72wnXmO1u6ixLqJRoSz8t1PPx
tcKidtQZlcMpFVjIzTReJb/t9xzo6E6qlBCUxs0tFZTgQqWJ3fI9z+yQ09d/3gZg
uRzTh5gvVm3nAyRVYA7ukCjFtIsHV/MR2XJ5LU/1p76SwjLzg0y87N3v9kZ57g/T
FxhbaJW/od1yi7f/Mn1OwDO8FrQeJkLy1GVcw09tCIutJ97EAsGIBz85CWViKN+d
C2O+IHdr7Y6ALU7XPP7io+RmhukkObJAT5ECiukgV5pms47q+ssvZhQabGMMBqea
1Cb6bMCkGGJU/tq8WUVUqO34XqngfG7Jpa77KWI66+eICTtVTu8fPzML+N5Mz4Xl
uswmNMepjpd1FgVwkjT4Enqx1ZDz/0tp+lU+uKLQorc95xyzUH2axMU14MxM1Hky
fM2GCGJPEjIybuuAfWy6tUAxrbMRgSU4CpiNy+iBSaqAWOzs2Lvg92olBwEmUVwf
AtOo4M9w/ZvIYvHDscWoG/u3L1/9vfJQMfcBY9yBAz7JiFXN1AU9itCjIusRl6GY
+iSNX8AvuRcIJ6VzDdwrE4SDLih/32TTZxfQoppImTGfgLgOKJUdBIKyz1Mbw0fA
xAtXemdiz4Q8bBuAOsRLTv//lEJ35kU0/UgIMV+GCILT/ixzbCA9ktPDvM+4P2YK
/+r3qvB1S+qB5zFq4l/OUG9SOK+Nym1zNE0n9a8/0ic/4CUUr4deWM6UNyFoz71D
r0O/DfTFKHQ4E0oiwi+UiK4nyTHQkmEm3btbgRGLehnF/irK74s1SwvY5hG7GP2Y
4N69OKdSyOgK8wyRKJl8vxFF5j2lRNxYm1e05kvt25uf4/egwvMJuw86Wzl+kneu
lxRkWhfBpywlRk7yLSGJkOe2/qCuZXdSZLfdeDo49u55waXutG1/CyVLT14X5Ent
D/fUq6Com29Rsj7XKVDBZqcaf8f1pMYneC2KFmeMBLj2QXa+9Y7JOW3Kws55JLiv
9kxV+Euq0aeG6e59kHRsfRuOONSs6Jx9E6PGUTN6JXEVO//ofFpjVmBcd8/+Z+ql
4LhQDbjKhCnwEV79XyVXQeGtuGAMtEKL88m/hoLzrQeNIt6JNfbLXtdX5O79iw8P
mvAaOnGrhKGCuyYKCeNDjGSfUSdY1Pe/pkbA4p8+4vtwpw2hIPEApQJkn9l150vs
f5Kv+4G8DtLsM35jAoiOc3mYMI10e810Aw2xwM6TCvd5540zo2UltGGrmyJv/Ruf
jHLVNpUVZDf1PuibEEa0X9gH4LexyMPHR98Lyg80PMop1XCm1jOEvrnAXJZRGRYT
0dTBagN1RgV+Sq4HSuBNF0mNgQoqVqQPcPpFz1wJH/OOhCDWDnPA7vIXHQI3IfNh
vloEjt1Tejf42QHPOH1P4T5EnE3h+lIN1wfXuvUGtnqg9EbNz/udyvLdKGPbjBFN
EQPtWD+Nw2mQSlBQz9puUNvaXrdA8CnfFfQ8skbgYOJ6XqQ9pJRBz+NUvV8CtSd5
kB4FHnBljbD87hjkioeIIwAY5Hr8kg3vfFU/eZ0DIY50AlzoowQ2VSjCYuc7bc2m
PuBnPN4ff0t4e2iqifm5YzysbeYhoM8YYSlP4MQPc6+tDb7LtzL7Iyao+YlWyj5I
WYGD/SQ8lrStQGgy8IBujSIARosKp/VUNrFYEP8L+CXVsUQ+Tza1oCn6mVM09UXL
u9aJN83RtMo2ez0T7gYicYAJaxzELvveEtw7Ei4Y73wcCYmpuG1UGzCnsVFmrx5+
wRtnv/4+AIFs5tDuFAY7Nuwvl4WRw9tunB/cflpb3Z2NmIvjbnx9aqrmphXtVSnv
7ZQ4pt/T4zZIgRaJvV1Pv6qwgbY+5R1DDMDPTsxR9SiNdsM6DhwTMqz5tjtreN5J
7dyZ49GUUXp4ynAJugGZ6mTVi7HDZLC7+d5p5kJPHhTBUyk3DV6MQWZSCwWO2vc1
jDvzYmLY9yXmfHezCU84o6jYtrVWPPWMMyU9LVASx+S9/BM7vWjznN3utsJiDeyC
kor8Thj7vJmg+0fCKi/L526aPn+6Qpo4csqlYyyMguHU7JbtGUUuryYKvwl5xutK
MDNfB06gO/vQayxBKzk2+OYFgfT2rOF1kevufx/jUjQ2QLX3hEJlxfwNxQbpnDD0
q9A0s7zPHwK59WOF94W369ed7wFgpHiJVQ6HV0PPMVxh3JzO4/cnG2mbgSlZRGSu
bSO1VZgAZNQDVGmWrAhK/fHWR2d2AUyP6Ew5PQknFQ4Dn57X5kFA67/TPBbMEf0q
O1AFnGdjTggHpHnnXFyRXdnQepUroeQrF2QPtmCK7ZfsuYRonwFSPBrmTcmtrU7F
i6eIZIlp6FJFvh4ay+tb/02bE+PCZmQdbpTxYN//E7oSD3ZBqe7bmLwvdoYsUFU9
gCRuCjqgYQsmbotTkgIgbx1YEtur2YFOoHqNUal4NY9Fjq4vGgNBPUj80kx0TeZc
zLeqvxW7QEph8Hy8NjTUPlL40w+uPnU0K4mO1AauOrKE10qRR4zo0hcFZQ8BZNUh
ZQ/zProMEugDeORs+yd4SNGZPyKp1IU2bqW5ytA2gGCyUC80BZrvX7corTbW16DW
zoyYLmGMcvWXjeqw84uVKmvK33/psNPbmYP+cJk2zRHj7293e2UujTg8nCOaZtOM
pHkjahLMNH8Xui6BN4o4RHhuAsGF+DXd2KdsuWMcAqBDLStgEjdYGQnrdiNcsHb7
igRGs7hxUR65oE7RAyVzXtHEqTGVyFYeBb/JXyHFxIKp2wqvlIy9qiB6tZ0eJPX2
uEpyKFhBwfyIMCvTFVp2yAEG/YLpHNspLEvrls2pFtP+RIs3tesiDA9Lqnb3Xf8T
N8wNAjhkRux9oQn5gDVl7A7NQFcNDlqtuZrEXcD3kUdXOplRYw3fSp+S94Ay8JRz
Hyo+9LdqihQC/kmAefyFlxWwM357I78t4wIdUfan0SBOyllbWcdckWL2rRbM+1TW
1viGNffjBsqvv3V9UrabfB54mxTIVebEaJhln5YAQas1CGRxpK7Xu+QH8ICBTdim
kVKG3m0sk77K40N08LzZqRYQ5Dco84+C9c9pPppku5FickXd4AooBbllRjk5PFYh
SzFpjIkEFTUNNJD/c3HayCCaHHf7hjphIW6DJmLrc1M9q/EihJonBS1SRgc859/t
t169YOhXTgXG1ODAywHSu7TtkiKXKr3SDbOdJ1nTUSQ52yzDErsG3573weKA+b+G
3F6oRR4I85ISx9vFnoOqgUY2kntTFdjVbsC5Sg/HGc35kYiEWawrHBa/fhWKGLe4
M5EKEsTrp7IvNQL8BEKvcOohhkO0s5bx0xUSVKVYTiDYur5yfMqwqPcWgeOBbiq6
hqX916C20Q/zU4+kXZ5Zj7xUt9pitgN/G5fZd1BHS2QVUMybXrRpG1lEvebeFaM3
9B0lnOVzWwUKCyvjBwPEyYleYt9346OLWws8yG79FaQ+nvwPXsmlcOTe4HHbBG/z
U4DBBA/OmpnTvi1n3DPAXVemxog8dWzAIYp/KUhUvlYD0M9M7fN9w574/XidaNmR
FL4yqyLmhvYLUrJVgZ3FHXnLlZAMwGWTLJ4362R/Xbxdp2DfQ9D2XbERnzW2GvEs
ZYVcr2Pv3BD1r1tXt757Forr4sF6/z6GWEmHD/1UmiZfVQfO8utkSnZ+ZhZHUHGk
ytntK8S4Rhy63xy1xbXk147CihJf8I74T7bN5nTouY+vkyXgLsLfx7CqIiv7YjjN
wCQTExoER9zCTuFKMbXA5uZ0rbvUQ+2ukAMnsWj8yvWRr1WSW2ktrLv592IQb2tx
M+r845NmJdXwqglZZki++lxkcxWrciLU6w7Ov4L8mqCzx4wZ9AUQrYtt6c51soha
y/MxKLhX+OhQqgwed+nIEpBBzlDO6yPeLDl2ET+cxionTUyR3MI0+s1MdudNHItR
7ySjAJWds07fqdq74hPTyYEKUGu+k5Z6Hc7Deh5a2/W45xe7oLQ7jjyAQHcveUgH
ol0aK1pj7nmS/7qOv99yDb4dvqgThnQ2wxk+IaqL09vxoAxAr49atiFRBcrhgtan
BAu8EFXFhvcwc9gzXewYQXc47Z4KVoQx8zGYS+Jump+BTZEq+3kqAjjD2ZEandBH
4eo6ZVTNoEta/9bBtXGosGZXPJ4Sq9KRr0C5CXhnUKF2vqmkHhYEpZFYg6OkqfIn
dB+DbTIVD6fkpV3LGJTbv5/mkB3TSzF2+6G8iYz71JaCOvHpU0OLDuG256yhHttl
Cq/z2t2qyFfsfJ6Jx+bPw07X+axvIV+RlQm4CH+61geE18BSBxxnZ3G3aaODy+jK
QZuD4Tj/Lzpcbc4bYcpWJaREKPXONTde6lrCmgP0QuCqmfvcAjOm46jk1rlos8If
eS/SwnDZqj+PNoquxvSloYmklPBewigdAcJxbgd7AvGClHEw/mjiep5slnJBqWzQ
aZxFfrV5kRbQT/fVTokRujcAYvsh/4zMV31OEGuKMmoFCRtDBzJxKz3lkMSRSlS4
E4CbTwBBmSbiGL09XOOlzR2BFDvtzCSDq0nJKkqiHN/4qpMEeeVFQeqHg7N3HuMP
unPeR3+OqTUVNyh0pPp9ArIK8NLxbiimdoOZIw1xWfL+9EwJoP9YgziZWpi2/Uu7
mwB+bETuDpnwv2uDZQgJ/fJMb5ZpzqSjZNGzzzfFtihOPXQVG9RUgLx08giKomDi
26KZ8eC07HG4dii1NubmlcMwZl5MvC8sZqMH+1zl7yqRMTs4TNv7qfEVoq/ZV4g8
j5HHoONpYVeRR25zSA33saOEgfwiQ0TxzU7xRwqEpw7l6dPjLLJwCANJfekckI6f
MKQ6gtrDVxBMZrv2ae1Fvpj/m+5zfTtT0eD8RWJDvMJ9JqRPTLWvZ43KTDEIcvbT
xUabg0/6xmEfcUxkBkHkbdFfayCpz9CVXO4kOMV9r3duTruQw5x6a6n04D9Z3dgr
GUrufXkbU+sPqA29CWUEAf5f7L4PDy4Uaca+DRnmUDFo0GNb1UzoQkWqHOxjfTZw
0ycGEASnnWsflKN21igwhgreDOKxOBEs3nZq8W3S/TIVaUEtqaMzy14xY/ZaW5DG
gEAilDxaDNSVetAx1A5DM0Gpeq9ICdlC1Rb4SKArOYAVmyx0Q4nFB6pg2EuWlEPP
J9VlUiOBvXOH2Ze45oquzSM2UvWqwGYR8Df4700vHYfDHljKwS9FaqoBjUgj7Mkx
8m3cFvhjjwFeslSvlcpYmQsW8wy/lIYwB0jPFiIy6v8sk+gpWvfqVd6hiPuqbsTt
RvYmbfQBekNrKaSKbGnhNBBOr/WsI7ari9IlIhqX9pg/gww5582w/rT7ClwSu7XN
43z7+1QR6CgGHetZDjEinTJp2VQKWXPQP2T5+RVYOd+TyQa08m3ljXpMwf/jv2mr
LhuW9yFWP86ngToescbE94ENV8b2jGNkI/dADCdj+19WHlMY7ygWeVbMJUur78ex
dNlYwYV/m3oSJyfLv4MFLIeorw32xCZ5afe0vS+8Hg70Cfrqv01RwBF8RCKe9xP3
miDjx4QhjhQQ0bAx0fXT40YV3gJ/9Aq9d2u6wKSGu7/l/aB+02hYR/100UNrUngI
Xqm9LXmfRzl8QjpxuhGF62yVl+iLPBxTXH2/6MkT4wSDcSUs97ah6mepB6L390jL
I8etNQb6PeNlhar3S620DOzvgVrWyqsYN9nkWXFRIDzl3Xf3tuqKu3GQ0Hbxgeg6
bNLojsHCT2FLBl4bc3a66x1LTrn1cK52ZXi1K8iQEIED9yuR2nSTl8WUJE2ebs68
B+kg4dNNLAd1E70sOc/MOWGdnUg/fHe+2wbjN1Y09rAIiJ1iiOhHZu8EMcwqe0kc
C8qGSkhdawZPeDNVn+IXK+RGu5h3y2R03myN4qk1OyuCDgMTk8HkAhMaCz/6HEC8
nTe+6T9L0/P6hda2MZ3oSvH8kN44lRmN4fR15RFuU7bkofPJBkvUZZqSYxqgqc2F
wLoBQWaNAfdIvzsRpvnUQcYo5Uw3y/GnxsW8x0xaYLZGQvIEYsifBNGg/6XWAriL
NijuWg0Nxd0eorBShB67prRVaIlN3ClYfujraHI/1tRkjlOQXdnGFFJsLdBhyAJQ
OBqTEUn4w0efUQNNW3Q0meV3UJhfYsDQFk7E3BXvDkPJSoqc2ce5d7O9iBzV80Oq
ZbAt3cPAT+0XO8SbxFDFoHiicezDQvAMvHA8zNf/4u82qpwcFhQ4oMbUfqSjwRYY
vownpUgfebb+d2KvslFNpxbCJsocvY10uRnxqVBAj+lFyugdlvyFUwgJ9OdueVIy
8gJ11cUoul1sdduyivJBnIUrVwQmpcbb2+uGSE0y2n4hl9C4expCuxbYM2DGAGey
NmEDeeG5T6bA6rqzGPUF2yA8Gp7/N4JupRDKwTfMIwZ+VUpZ5b9jngjbqYoGXNS8
MOA6BC5IPafILYnox+2MwVNTbrUhwc/8KG4SVTck+GMi4URWuHFC9NAp21B7vAiT
CQqYOtk0L/fDWo3bMDSMPkEvDaRiJ//mD0e+OCW9FseDOAl7cCPCgv4fjMJNnutG
37134R94POPKJUXi1jjfxhc1EzK+iAefr6IcvwOmQ3w1EhDyKRWGf4MElMrcFu2g
rlCyUzn+ttswwpNF3Blg9ythvAPh/jHoO3yoHsjRhN2BbX97NI6K3QsUVmem7ZCy
CwALzg/nNAgcYS+vZbdoWH+V7oC8V5hSxqGQuzM1eVjaBu+ghQ9JNJgGyEH7mIRw
QV6Xx2lNKAlOf6JtI2yQaniVsNRVf7UwV3nh1/HxlIT6q2XXRvswWl5kQuSiSxXO
eG1Zppz+X7hXSGkaqErq94tTgPNBWQqHRcL807UeUvjKPrqxompPgy7GFB/rBzku
a5Dq4Od5TjvatXl7H2dEehqNEFug/3OVALcNWc515Noo1r7JCHfjfPIkfk6vYEgF
OouHFXstd8sv2J9qQwGqTVdEFAT82T7noynP48qoh2jODkHzXas0d72yN/6Q9sqD
pDGnqcM11UwK7868li8zsV6KE1iG8wSTIoNP7Wea0LQRgeXlyfXRxr5BxxttuDW8
rGT2v8NYFmyxJTZ9ugQGq7xr3zQUg5/u+o+jGlElDBmTV/XooGFl/66WM5m14/lH
hbjMne1X4iqB/3stEUg9Ts3XFaHcdlD/QIVjccTeUGDiCmPKYxkUBQw6we3Hi5Q+
yeQkdmSCmWxLegcCq20j/A5Nxt81ZkKBFufb9H4Rb8EsBlbAQa0HcN1UDqfSxlYI
0Hop+xTueBjIT1TJjOoTTU+fzA8WFA97YPWUx5ZckJgHLjYfKKwxp+Dd8qEnvi9f
zebNNU3uYO9C7cRKhfRObXxCivu16LOECmhiXo9ruG6kB6110K/u/frroCPK0EWV
wdMSGzFWANiBzVvVapu8pnnEcgkFObWY0tTonrIVM4JsdW4S3bbXztkD+rGJkDeJ
5WSh56Z+YYfmJfUKeq3LKcJESpjKwCZ8fy97JZB2YTic8+w76VQK/3VEdgMyGvc5
KlRP7uAOOyon3b0HdZyqhfIKHc48s+7S4Tww/5z0ehuRrrdwKcc5pvGR9K9hffTP
8iMcul3mifvj3wFRqLckuTBl4zIv7vuaG5c9+zLfY4AlVTtVOzoTCm18aJW/u1Ka
drp8eCrJTn1qjQpTSXgLnzt7TOUxu4/953SVCwi5XIAZ3ruozpX2HpHFgL5dSLaG
JkepD5FvEi+Ayn/AnoM5LTjK7Y4o9AQq/X1ybk/92kzfMBiw2bcSJUZ0QkA6A0cA
CF0Kmb05xv381Ap386rxVMITPP9o8DCNOeCO3SJEM83NIb1j9JRaBFZ4r9q+AfzF
U0Fezjwes50sgV3FNbjUcLAOxiFw8VptiJxNwwAMN9ACTW5O56fa2jh/8RHICFgE
gQFX/KRNib7fQq/9Gbwv2A7Hh1Y/WGsuO2tYrio39Yx7u0bUElVtetZPVLBjB35O
FCPFeOi+4J6bqHhvle7eR/9ICVDVdSIAHJzeLgX5h5odcQEHA1bbRrnrmTZ5p9Nx
oez1SJYDGBvNjpKxU0uZv0v1ZsXNH57A3q3AaO61yU9d/YDHHudjLgtInONrUMbX
I4I8xQEqFPDwebISHzh+V42U6W809KIliK+Kaq97tfoCfo/FRj6UjE2r43vex60A
0VVJ4lun3mmLGuuyMyqgk5xXcx86KCDNuk/+nhOEc6J6gDk3S3t1X1GXJNuRAl8P
fq/DKSyM12sluhJWZ6eF4WiVC6EM85JlA30V2vhXzJpmmv1foSPM54gSv03035oC
FBllERr0w/xnXL/qnCzLpSyIjdutxE4MuOYKGx9eb6ePaWB5StS/qYELHogKDpXa
/z9jTLK0TIiAdNrPoJ0t7aPnrgxiNxxwc1ZJh6+PbzlUHniemMLAgkdB93M5xsIl
1i4BPVZ/gu5d/GTNFUiwQK+fHDOBNCbluIsUfh6R/D5ts3MuezClqkINDs26UbXx
ulB4L45zGi5VTnf/0m1zGwN2U4SN6VpgZlzwAUSxXRoSA0IL/9p+VEGBQ/fQp1jU
nl7yFD13P1erslCAtH1j6yvUb9JAcp/pzDdGOswGZlhY/HOM7L8ZHcBrc91DOePE
VTEZElQPxReqYTPJC+tYU7nQoDcW/gZub6Ojt4sHPENHcgE3FuF+KUpvrughVBmQ
vHUW3kpzBwAVGghowUyFHqWGY/ZCjUsek2aKWwJ9yg22Q0ScO3rOBHNLtavnGPzL
WE4wPBB9sReYED/CH1wGEH7Mq9AKLBlTEucBZ3u83vdxl5wuYVyphIZeAyTfQOLf
gX9iodr9hfgWGMiws//ihviAD4Kqj9aH8+urawxT+2C75QeFKJU/9NYlD6qhkmHs
UVcWQ73rKqZC5yw54H1G1xnKXbNlxr+eurZYtM7crRcGl15BKAjz83L9elo2fiWo
KzfGc0j9dDrIwEbdPtac2U3EWMquoulHCR9davYzZPeseCt0Io3Pxnos1310ZY0G
bXEI40nf6cac9NvMeQecJAAJMi/yOOTdBreON8bj5yJ8ruAS05SBiXdfG9NXSy82
zPjng+/hdSZQu8lkLDLvPlgh6iUVV/EHYIjs2Yk4yMilcMk+qiZINOCWQo+prdFl
eqDZ6dCbv3HEYaHSOMHTLgvE7Ak9mzBHTyMDaNDmJUgKqDGnrIu1ebDqWISz6T8E
AfX6eao2q+zG/F++68bJxtejUZj/0sMW4Mln1CvlnEqJn9+HJmEChzmQuucWbBSi
eHpEBqrOIiHMRFe2HiD05MnkPYvzfVIzNUtl3ex3VgP+GUcHd4Ht1WN2r/8aNnsO
71GV+ydB02lOWTGpwX7NmXQKbw5Ahe6pvoxyg4norG4Xk4HeMpBWG324YMqdZuQC
NH4LaxON1NEI0rG84xxwuzBUrxLV1aT2880xpWdhBNgnUesDQoFTlhOySunYWNVF
nmQVNuyp/BTRD2egGazkxHMAyNgljjfKJL6uJKOg0kzpa3Mgz2kY4++8ABjGk5Iu
HE/qXbkIRFRcynf1w+u8LzYi1d1oDOZwcW/pXHavkGvTBPs7PPzoGYim4Ueedikz
W17ZQla691rMdQJqAM1PlOU11YdCDY8omGOOELQanXBePz96bNN1oYobHGq1+aL6
U1GIeK1CKnWSo7G/4XkiEdEVVxJ0Mp42qUynCSm2P640laX3lkA3v8J74L1fJRVh
goSm0WITvp7hXquyM2fY3qKyMlCU9IU3alzgtMhpMwJiogaGfEvegX8KrkSwx6Fn
haledkb97aBsbnhtnNJlOOI0JXjR5dp+BLakbAuxKBn583BALN0UhuSF6uGEKjU9
u/BjkL/eICf3UtqNZeFYFhPezxVgrfqy9BGRcScUeHiMWe7wX9TQ4ZrpJSrfOCWy
geBcNKd1fLVBTVXCFd/DNYpmeIBUmV8sH9LikgxPSqcD5YDouJ+SQIcs37I8GsfO
wiMGzwIybgVbI+3PZgL6zFXdv2SX4x4NC5M47JBHcSNWePZitaPHveXtV2p7CDqB
F5JSu5QdlEbkokBSzeuu1olgmU+5+SWNBYS6KUV3WgpzX5WhYGqsxd6spUsVE1se
8tzRMTyIOzB5WZFubr7gr+c4OZR+J5nNPDvspV7L6P63NSD8k71UJJQfJYZ7gXDm
/fmRLxxVn3oAtoBZ9H71jeJZfauwiZeZ6xvHWiK3LYTOQLll8cv4REWdexRuGGrJ
QsUHWgiORajweqM90pKnAUJzxOwlpWWcd7hXjm0SEC2BC3YL3Xu35H22ake0x2Kd
Q4/0hmTUja6THIj8NA1LMrPBiWcRCqmL9tNny0OmSbLvd8sW0LjsMH6i3d8gGbYf
qyhEneeRT4XsRSBxEvqNn+fJkPaeO+Qis7eY5BeTeTscwtTrDXmOzC17zSTEABV5
wkn9DgU1xZnIhntadf7ftNyjzxRH3wFyJlJX64JaBLbuHE1YJ0BNlyUVvtJhRHB7
ao1DCKno+/SUP9Ycpa8XXjcupox5aGdcdFKMdYj7YPcQHOO2wtxukW2euFeU/KlK
ToD92j03+akyXwqPjft+xotd34lgDE25cmCbVVAus0Dj/DHv+9//hbHpV+va0WkX
3dBszSm2XVyKDG4vYe3l/rvW4QI7ibElMpGLI9AFIPbo6GjbSmPzVQnCfL883Ukx
BMtuN9TMOrsu8IpmVxvu/wagVTm7PnRjQEinHnOhRWO8NRpVUA+zlMcqK7wb69rg
CtRIYm1sDfA83wGAfLUxESOalvLUCwWF2MJn2PmwR1zjUPOGubEXCZLNTM7HYl7e
h7bS8Q1Efm+oHXb0oGhQeu3KH6awxvtb/gsZkhPCqBr845uPh+KOsZU+inhrGF+U
U8+pvw5MpyHdzbujyAreYATf2MuruCX6xaeOrZ5S/0NEBwQwTouW8PkhL1KyVAYX
rvsD9H8WvwrpFAM4LrUgxrfGrb9O+m972OsjsJE5C7QfzBsRyw+FkwrqjYPjRzBb
MX2PEFyRfJqKWOJyra6BrB/eFrOckJfe8QU431qV2s/C1gTOpYUROyb6bJu3bHOu
L2sxFqK49kpDcgbgbLaul82kl0Dw8HDHxWZG6ukKivfLxY7IzHEIVONtsAW/ix6k
XqFiG+PkwpN+ErriR93I976hSjVh19tav0puh+NiH36rcGpbF9pzz05dRPC1KYTc
TtNGQixBTsqWtNfa3lJWLrtJLkY68l3klc8+k9Now1jTqgjewBiarNrtNmP667ry
/FHtnEeaWmJdO+FT2HCDmp1D6RjMCHE0VppRUHitLNe+sTXEAu2vBLH+JkwuEFxV
S3CDUSv78ISdUEBhkgtBUy4SQqij/v3fNaEqelBCqvC1XBOwnjpYaOs5WSgn8Kss
qgk2fhLketCAgxrCHh/7wVAnSFYUBPznrni+YiTymMugpWb7Z/Xo0PhQwND7A6id
aBlru1lO3vldnOR6AOOP/FMd175vFYnxe/Yt3v1cyENCGHWqmKCBnz17Tm2Vllv6
RwpDzXFdTztb5SVsWC9nuL09FCCq+y66eVbSUIK7AEkC1vK0ObutkwvG7/YDdya2
4WWbsIQz4UE2ICRWmBaJTr2eEYXPHY3Z6k/zcEljoMIpZ7HgqMJhcVcX18eyHDh2
Jy7UVJqSke1TdGWtLT6gteLcPh23TcGVEa+2ruEiHEqoW+l9UGw3yMuWNAe8tXir
Dkzfdy0AAcVXzkeNWPbEQOj4GhBG9GIZSXvRRIDJibjOj4AcCflBqKfPYiuTXYaM
L02PS1s+pirtbdiRQrzoi0h40YNBSlkvFteUgxQ41qGnVewXxX8Lh3WylgPaU5xB
SQK6EOt3QCgqtcv/xN4tRdbtERrKi8YiHkqLHvtW/KBgrIwYOiWJuK+kryR6xwTk
l8pb8SR97e156gpyYexZ4oDTMFoj5fLPFVWoIB5Wa3heAV9osf462YWJjwJ8oJNF
8bWzkCrHAg6f+mBEC12OvsJibfZQh36Qa+jwFJMTvIS+JwgbzEJgO6FUsCk0HrqJ
BXTvI95PjX3arPotrzectzKsjFxzlAF7K6Dsq3yPkcB3kFUZkfiPQqsVtGfgpPe5
WMJ+7rrgk6pcn76c7KypRdlYWeDf8C2yElaTzTixiTWx9Qio3/EF6+SckG27I+cY
zPkCu5AlbBWYAJO4dODvQisJh0/nOcT+0MT21JH9qN2yjySQq90taSqGlrKtGBvl
/B1+NvtcjL4dCLQ6yCPEqMVNC+6QHZdVXWHgjw9ZN8NSZ8mD+dT4CSiH2lHB8SNO
hfYuLXsn2hlL2eYv51d2eZp/A3y6BL6RpWKgLNP0dkklXym6mDAkBM6JGqsDD2R8
uuBgRFj8NhD6MyGPVILsWXSKyf97hlt7jBi7qUUkAcRSprdNXsx4tQYbr7+xy0Fm
HmgqAFYL3U7Qh0xSKIZ3JsphmGG1Ubcf3rbiSZSyGAKPmXXqkxDFf5CWDQdrvxJb
U4FTPfzg0kBKTqVwWxU6qbWs0rZgNPO543y5rJBo1ovXXhTqw2Hunzz93oD3QgJ+
Fc6IHdIfHqiYWnCKYKaURr6fi/FWSt9KUO0E+b/cTX2ulESayV3i+4zprYDJ3+XS
W53aaUAnRO7ap+i91vl5jOcD7WJq1qjMDOc0qRFKc1/NysVcMjSHyzza6d3NTfVd
TfHEYaKhsRp20m5rzlMIzEU7mdzX0j085NCKVGQHxPvM/2TE8yip0+bvaO2APgrg
EZ51Ri/Q8TFDtVpKP8zPy++3FPFzRLgy+qVdKjocqGE6o9bFtuqnegp9aXAgcNAJ
XSho6rXIinTENNAi1SnGhME9rMAr85Lv4GBNi5R4S8B+MNRZdBU0S1wNkYcXYqdt
DW2Gk0g9nYjQ7/rRUL/wVa1fSujKLKDh1WZ8ZhBSA52+zsc8bVGDanlWi+wy7WiY
fVeRIH0x4IqeDIcwHUrHXssX1NnjXuFAr+1WNjQp2V//Oe5GgLMIeCJVOsiUVblD
ezEUweg4oFHvoWmhjDG8uGqjEiUZm44PY7CD7y2CNIovT/HgKzpGDyUYDftrLW85
hPXsYI6Wd+YDzR5RPjDTAxBP2moos6T2srFtDMHRLjRQXDCWDnMcs12Wg7Pc+Bom
N1tq2dkNLnYCd/3adNNpyG49O4FhvKa5WidBTK4CqlGzKj1R7b/pNXFEb72kEIxU
NbaZ7+ZCnPpQdDejQ6dNqhLY6nbOksXBWS7YQoHFe+aBNgdxe8IdxEKYmiTfhSlE
4T92Nwc9FkNjMTqczO6w1Oc/Ru5wALu/VT1pd/d2K8X0Mjd52mojvsfozKMEtvEp
N+NTzh5QKewIsTNQupy2ChB8xu+UVohXrVQ5fwIhemvywrLesH0MblTK00bC3KCI
k3AmbLC/kkmT5nOkE0vuZm0U0PMU1miTv8tpj5Q7BDffAwGYYHnw4ARlXmlpkj7x
cXCWqFyHTmGjkNxxFgI+xKzu69YL2nMdiOwrD8zj5CK4C5A9s4Fes323whEtsHJg
Fm18+aaLKGP4tByt5fD2QJwmdeOPwMMPq+FS7bFmqjtcmn/B0DpjCQlMS4NAuGqp
j99LeZNpg2lNJqy13OE93Ko0Ud/QL/GGpzaqo+K8uNbVcwDfOcojGUS9T8lajJmT
uNfdE2Qqziyy3M9gl2utCoHwXljqOgweriVvJnIOJD6rdEkZWVoSyFPb2DO+tWYR
HHd0H/zeBTHd1KR63kb3MGnklkFNp9iNGacdemOoZ3+BJPZikg5EP5iDdywloEd1
71aMVH2THH9Vd2pMT6ogkvt7qRLS9z5Chq9LQUkE9JbAAjtIgd83TtF9N/jgzOMh
X4kfG37oV7U+GLjIX3VLCWPp66bX1EMgqM3iVQLh53G2VoCjNNYF1iJt4vwqp8qe
id/bDlYzPDXh6lRnXKJXhxmhS36Lgg9eZcM1IEJwPzP5Dea+w498lYGFMMVphpz7
d3eGn9vkyee7S5XiIaxnY2/bdWLLJWixqEzk/FMv+5mEUFlq9JUyq6UgYPjgQy+0
Xtn+qY1odaKIwFDEHbJzUdqukFgSMKs4fxvuMkkncTaHGDnC/uQQrYhZ4chq/lPT
kYg4S7ieHSUQXUzspI0vwAqC1tjcx4IIFMB+H7Xw1P9x0cJD3u6N+gylfYxnoPNB
xdbxeCOui5kq7euj8wdQlO35bX9WqNpWPcqsHaDfimoMeo1o4OhxQUTcyJ/k7BJ1
VWPgM59QQV98rZcyxviWo/yFvzxk5I+8XQya+jmdNwvijGrKH7Vn/1fTr4l41sqn
f2ocO6sQ3d020iNnRA9z95A6O1rMlK12XlTrhZHqbsKNE4Di2rAlJhwprXjlxkPB
rgMJ4E4+ja87g0ckakGrRTF1j8cVEhKfPDUigZM3S8NhqcNA9+q1/Iba8v84GsKN
O6anUkRcxYDeQfaiG8+JiOF9D9s9lUiEaeogWyRMX/b7mc3nozEy2XACeavLE2Z0
KH3NivKuLGiweBWz7ROyadcd7wfiRNKEGGevWrLnyTogEG4oZEMZsjRwc/I9kkeS
e7SsZoLqlGd3W6MVCQfZQDxqnv6AFX0gxD252GRx1IRmxqE8qOEJAoipn95jPsmk
3QGvmXYmOGnp9hN527Eh9cNhC7EonSZ66BSvDhM/foLlNuV8sktOiVoIyjWm5oWo
VfGfskowLClLpTtWQBvVCkD8a8PdpdOWTYrIlS4HrahXFlP8WVW9J10SL2bWl4UQ
viuz2CmaJU+7mH/p15PqT51iarPq2Y4xSIenqJk7AsBC0Z9mZkDtXK6k+lgt6w2E
4h1BUV8PpjKkxmw63yBXFkp0U5tqhNH7hYR8LzczJn74JNkqwLaClVPYi0W6FTSD
71q6MElfBaVrmKIIBOEODRaE4UbBAHdug25s9RMAk9b2bNYV29XXklr6gAuZrv3C
yDQQ6Trn3ohRiGiY/0EOO+0Z6ckBCOh9Q6rmAtU7tG075arbY/GtPyjQVDMeAr8W
5N35iAHs+Ieh0TncAWhv+0RdCYoFE+miqUGVFCrOt0Esqvam8y+G6pr1bD3SyzlQ
1ddjtlgxtjzY4Sf+9rB69sHaDhywN/U/QZ7RyRH3ov2WMuE1FzCBE9+qPn3JA73X
5EihnMA6jQo/+fLWQ7bVm6nBYkOYsJT7pWl5zMA4cfl5V+I8+E9sG/NEIzcUD2FV
sy2+hly8zxPxVYHD99utnqOeYZLtFkgcURplNrggCjwws8zh68UC2F9jqVXcMMU/
W+a/1I6U/Eu7Re8aj5OEXMu5Mf6/vfeBoNEfvG27189bS5Qof/ZeZzx18OiHHUFA
xk1lN6SnIJxOp3gjpbTiG6FaXHVFqpYOa1nN70VzihH3rwdlELUGmtir8JqEw6sH
A6PD8oX01/DzVQGwmNFG76QL7U1Q/9RNRF4U6trrwUm4HckbNskmPRShRcEQF28u
7jZkloVjG3kLaW7DGcsipU5fMVlyLnuqGaglN5Iq9RQtJBWJGWOc6jKmdslvec0u
BwWzxi7NQ790Dq9wm3mYYS+kBtXupFAk3LvQyBMJaESvMI57Pk4p5aw6+smTNBYX
TP9Bdd6x45tHFh6j7dqtQ3UhjiGFW7QlVfuqV6G7y3ngI7tJDgI4itaTJjc0fzAm
8GL+18c3e0MjhgUWElYlXpUQ54kJmLJdt5of/1QtUQac8FmUsIzIOPdbCkf8jznh
3j8OYEVNGUqxoIzSvnqu6CJ6iH1NP3IMiTwmyHrm2lGNgiw672T+4Vc3QRdjbpE5
4DCuGG+IbRALFgDT3bnULUtQpdBdrDefeICi8JLD/VmdyYEwZSBSUCuMZhtLH3Qf
ZFx6JvosXD9BlVBt7/VYSzfxKkV6DwMDCW1xb9ouwjQL5R1P/4OnUvo9w+/Y6u9D
8U7GKvq+oeFWfRNMWnVkWPkxwxlwjbzRxcQcp3BffgGy3FRWVK2p1hIlXSkcXG5q
yTIdmzSF/5yTkYdzl81X0G0nL50Zx/RNg7ki0/WBiwfItPvkez6bkwfbgk+s+CIb
20GTX5euv1QIt1uhLDH/pavuZWVQLxfogzTmvWAYo5IjL2P6yS+LCgv/T6Toc+jM
6J8v7ZfWr8EM2q8OLD6AOX643JgG52zYfthqNRLPQ7TNXBj9YgzFlRulSGMtwnVZ
L4bK76sr6nTbbqJyINLgZ6PvbGDCYaQxcbwRVpi4cqKVyUZ44obCJwpqG1IH6fqn
ITBpyjnRrBT80Wmu++OGn7I4L7K6AcTTi3nyXq0CfPjR97S2MRYE+kzxbN1uTAzx
4xllh8QOl9x1ZfdxAlcGvOA2Et6W2WN+8IlFK8N8DlZWUBmJ8VKgAYpjn49I+jnv
rX9uGO2HUlJqnOZSg5b/HS+87ifVDCWJ77Tq2jjPw12ZRBncPm7g+Y7x4p9rXT6+
2eVFQJtn67yFzGLLwTkqd6jBbJRmutFlwWbDDi90kvB/nhN9pm4Fe7ao92jY+p0/
vASbiPp3TFo0l+Vq1EzPZf/HKlTy2Qj4tysx3r1AVbrZKvTjT352r2vaT+uYbtZq
RFKcpSBFgjFxMMDhWz85ZnwTHkBvON7aWBzuNvgDJvGD/N9d1ZR8DnxiklsMEM4r
PxP8epsKDUtQ7IKGiX1gaK0jv3jAJU28XBL8J9neZyrHbhv3ri8IEGjGSOhWJslx
oaZ8ULyia8eOYvIYmvwY9iAJmQKJxDsb2GXr5tmo3I/qbWo38mf/UHY2eFeWuM6W
qCV3uo5nnTNUNTrmNa1qjcSjIf0I3sjZwpraklDGmC8dJbavuBuNIi1bccweBml/
oZLH6Bu0Uomh1sWowz2vxklQVfFWfs75Td+/jbHnvXO6jh0S5Vkp/mW2j/lBK/CK
mpI+FvnhGfl6h3fxo+JMt7PNmmBAw7M/Rv/R3Xh4pVvXy7tBCDxDsszxWtmH3R0e
QWIXKxp0rGDVOpEfHJ/acESVJHeEP8DMGxwQV2ncs11VoNPOJuRquCoISnUgE4UM
b8pI7ZlQ7cVJzTn1FDh6bd9Qnrj9vRe0qEigmza7XDAh8ZuhVqAEvjo7T2g9J8H1
pm4lRbQ2c+v1eINVtuy13Mijy7m+dLAvx6xdKDrXr7fU/P8MU7FdzcT0rFuwYyvl
SlL9oPR2uFH9ElbZfVTMKtPZQBygNJQeuz95cwKNnj2McRRGu9MhEBE6gi5jLLVi
HHX4lZf4jg1/irbthDjMZhKDQavovyOyr3rJb4xM+R1WrZoQTULhdbmvWmB2ftVk
ZQlRjQ+8C1VfwPPtzlaM/wpo2LDNfyf3oOHISdEiXBT1J4AgndBbiC9rqgVt2e9e
Lmz/fVBg2G2cgI4SCMEGQcbhRXHEUZ2IZbx7EWzkKKz67fXsjDEgkw5sJKmdrwwF
kvckOOBK6/AdjRr/Owwe1fyCccaMCZUeKvG9T18j7dfKFGMWzZdB1ct6O7GWzXU/
YkiphQwJns5GN7QmOcZyEGuFwFzVLhCEWEwSkm8ZuAT3KXAoeZ+mkOMc8F32ZDVQ
6Wvf17mgEOEXISKykuw/Epn2Pv+JiWJWvo8KfYFBwwymwqy3Wc4f4TyI2ZMht43w
bqVX5RRdiTRfDCHoyt9TPWIJGBxXuj/V9PmwrziMWTwBFd00GJB8m/20cnHTR47J
ZOVBsGiMB9/fV6abcgGYrYEPxM+5aThR4HW2OhWiSSinIDSs2TlF7Yzf4P/U7yWI
DKnLYLL0giVBNnXjbyBEyVxfg6TMkB+Z5CuAAtCGvBLoqf1Kr+lUpvmK9bfO4w6+
cqLU06AidVJMLZ/Qznscwt6nFIZsP/9yR5OOozQgXmjY+uE4oeL7SubY7bSX0Jx9
ybqsDPRODRv9mCYmEB+2pg7Usj4ByMuG6tftHX0GMfqNEbjDQwYLWx44d8NVAnHR
mIPTK0H9j4uQA77Q75ImcfqobelgOk4URxll6guXOmcx+POCwDsAdaF4Dmi0eeLZ
9gw4jO+E5rekvzVOgMHD+KTDwVVs7BUArMsRq2F5S0IWzWATDG0+sl0WEofM/w0G
ZLjsRmTmPfnI+Tc+XC9nUeQybvmsq4fqRVrD8Tk19rc8ma9jK3KrIEQ7TbDMVDxy
qaKFMy/geIOjOOGN9fPBWE2SQ/VEhXourc+7MpgvuRpbyi+mcPJH3R6OXRdgG3bT
o2OUq+3oIBB08lVXQuokZGEN57EheLgj+08ht6N//0u9Y3j3eTxg1Mjid86NbvLG
y5M9ni0tGyIPK8phpaIYtJC5cnhMAt/85tkEXf6V+zkr9Q8t5Vw67BQ21vpHimXX
g55Ar0EXUSnSjWnlkwZWTdsuBZpaYN1Lf1RfVSktGlrT3jOOmbVMAWOndVEZ10zv
nFOI63Gj8PJ/pEEx1hPFvybCnjoPaDf+QviNNgPFs4NjWppiC2BuprOkV6wP7qpz
un3QpWVndK2+OQhGc96LwapobiECoa3uhpbBTNqM1DexW7S7hUS0BlbQXAnsLT+D
0FPfT9TAWXmKIwRgK4e8ojU2bLlqhqXmzbCylALYghUEVeLkernrpdPtpBPv/Glc
AE3gOoEgQm6O8wpqNQkwkafPTeGzzGgp5qnQQ4CDhi94yl9jYfKQ3KUPZ+kq8f51
VQHGwPa5NfbXt6AwoCMcXK0PS1ru+tk16tdsvlfsQfrbExBRlEZYFcYjPLcP/Rbk
DBmThE0X/H/uCy7b4TSLYGEQIRTAx74m1c7zygHj2fTVpm6jdx3qaFoRBNH22S6y
Nrjg9kpSvCXENPGD1n3bsRQXF64LJ1sOhqdpufE6Av30R2i1GEabbO/LAya6TueL
88xYw2vrk98QIpA5LEeTenL2HDF4pO4DLsxnNULchMbTUWsbmuW2gP6sRUGW1Qzu
f75v73BSdrcZWSk1Qqo2Pq1NXVJ3h2++f4/zQaokPnNKLp18BBzsGuIusdDfKB3q
sgniulm9kUYxmnFmqX9vG7nDN7aoX0OhZYCIe615thO77yPQDMjy/PHYewwgJk9+
thlrmsT+8DV4WFkROv8LtdjkzN28lBKgFdXTruFAn8YviG3L/ZQxs67BaWbEJm+4
ICoGWNpIBPVpS+ze3rTYdnAgLPzE3kw3RgvCz/aXZ6X9w2hVCu1wN6SMV2bFlQL5
6B8fZlApQJHPx6eMJj2kbTkpbV71CHF4ImgoSYi2t9rTYwi2YvKpRWJMJR/osckw
ujBuPAocpsIhuTfI+rFVx3UXDhS5oPEusV0Wu9w/YhpYvYN1aOs9f8lxp6jnLS49
aVqulrayzsJsbB9p6KJPLg/Y7tPrgdJO/5whOYfmaJAtylfzSyEHA1DHA13hwHh6
Zgw5mIMCvQGofNH6SFN/U8hW9uyJgioM6FeeuafUDtL2zsRbCc9B67QZkCEwOw2Z
iC96tcWabBQ8RssBZ8rKKFq2wcRSaQbmxmnHds3vJ7dTF0kThhRkXgeB12TiB/DC
8HNc3z2rGoBswuWTZcANZrYu+yPK5SfCyIXmJfNi5l323506xnJSrwxkCU6/Ji1F
UWvRMnjFP8Z4LwBkWD1TcRUrHpNRkMfQuLBjlSJAQrNXZa/XKpskl7k8pZ2DgM/W
sxsEad2nOCFGl6PLNw6z5fYOx5p/YzJzwBZHma2x17+qLo7IS/PuxhaXWgWxx6ya
iJB/SUw0TkgVmFfF3iyHP4u9BXocC9UCandq0rA0Z8GndEDhuDydJZ/UDlUF8K9g
AtkKjb/1NO3LTfq4aG8fJky0Ljk5s6lGEKnss9rZgno5HFH9egmONhKVXvcdL7bD
OHuB9LZYrOu9aU4Mee9ctLsn9rHtfQVbhcMxT30qQAPAedWY9sE3DrlU2O7FI0ZQ
crl1jHS5b1JNp6nrnS+K/2LtiWuFjYuJZpcyK6DZ6Gh8q/m8GS/oP0cndG0hs2xD
EUmPDHH6Qwomr44DAjsrEtR3QF4ytve5CUv2HWbB2Laa7ckfhE02WKF8ERMijZFU
eqJ4KQydH3S7D4W80n4/YVPJNUEMoyAoUmveM0w0ICAJxeup/PBvzxp2y7KMdxF0
JxvFYpYsKNxjEUD85jORHIWM5riU9hOWSecr3OjJgL74PCTwDFiEOMZIRlsMkNSs
ylCOpnBxRWKpvDTXitcRJ+ptRwS60HVQpFReTQGz7Skh8GCNr1pwIbDVeG8e+L7N
Q2ud+KJMY2LeUHtLTbH7CihUy8hNcJo5DCsECT3fS9iMNu6xZZDY4+3kiEuAba4e
3RZ5Nlayb00zzOhozvGvMugIvKP/OyZnEyL5YfeiBIDf26R4IEMj6sz7npEMn+sY
NtxkwOwT3t4s6Q9sJ4PoF996MpVtjIFHlGVHaBStzhM=
`pragma protect end_protected
