// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qwR96p+c2x1djFfLohmI0osFmkMq09RGqdbJGIRHfGl+8/AnPiaNHeYkPPoZWA0lTPQOHb4dCiuG
iXZYm+VTcw9emYaBDxNhmw5oicIhZ7PNzp1hFxcLcWGdDNR6xx0WQApbEi36dB9h4zafbyzehSjv
WKKsN+vBUV3b/hnIPDe8pzl71dTMl0qV7eDNLTDMOZDFXu5tQLQyihMq3C2L6cUl8hx0bSeS5VJC
WUM5N8sadtSac2fWhGUoQ3yeuroi+T49B3fNxQTVvrp4lPi57EQF3vUndtzDNRJNEpeIIPupfcNr
eoD03fjUNg/zT/eMgCgObEN0A3qcsQ0Ex2G3SQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9264)
8kiI2t6KW8DdZxNEmAecLd5OSV2iBm21jHz+sKzGEG0mjuJrF6ikOLkrQ0C6xH+n4Jq+M/1Dh6KD
p1XYaPU5O/njOkVEWVpzlKXTVrjlUyXgJED3+nP+rfFmrtRsU1badm89hMyUXJ4LHARfU+3X3x3W
7jkCvjaoLIAtWVh4HhAOfpfmxJ7efk66b71z5Ug9CHnh8xaW8SoJDbCNEobgpP/8/YftbxjfXw1t
cwurFQKkwBZJkQRp2jCIk87sS9qmUT4DkjZhC6ELPK2uvJd/vQur8uKzivRDIDWFbCCckampFvC0
9yEmZwFTTolYTLSME/szx+40mGzmDsJpvGuLzbAZQ0OM/1Zr+Vs7XPj4LqANbVz20EGswj8dokkg
2nh+DmXdDzuUcjjYoNhsewJXPre8FEo9PLC70xydWe998Xl9AbK4wKPQtSqo+ggfAi9eukiyte4q
lT6WFMx4EaTYbp6xR2r/bv65jlLBjtUXgh70wqURXl8h57wpfhQXwQ8bcG0PhNFFkSpJ2TNH4/eq
M8rIO4/oyHam0c0QM9yRZ4DjvY/wCZk9hNc3JSTljs1Ru2VVUItVRBfvxAbF9Bp164WVc+e+JrC5
GunCKIbdbHJGn9GoyUHWPQc5C+KVWwYozEfJFwX8L36Nky2IIX3+sCQzRBJ1rwH7c7QSBItINJ38
+mdSq2FuJwPnuA4RmcF3bMqtq+w+JnBCPnM1WGXx+s9XgFs7uHwywmxrtrVltjQdrKP0UyWKFrwL
YkRRBgLLjff1Am3zPL1JWKANX6PTRj6VAYiU4XKDUFi5E7b8O4zPB7hRITfq7jumeS23JO4MLuMq
Gy4WZD4ELY/0CQu8z15o+tNXbwMMwiq4wZvTK/7hlXh10h7nFL32l6O7YauLYR8t1aenPzfqIDQ8
N8bMvozBH75THev5/fs/L7jQXGz++ciCi3hG2IAMDIaIgih2xdrJ3MCCzPa9gOgQ5PzvpJ4gTae0
5MRRjn47dFZ5ASpYnJb7eFq3LFpO6CYMyeH93gJqQ7S7LcqKFPn3bqX19fqIDRIctZrxqVGwl3lg
c4FFaFUlwaj+wSmP9QgEYabBj64Y5ezNdeQldG6uciORI75I9WADvzdVrWIHGr8wDOsqGUJJE+Uy
hnK04M8V9UVcGEnO3rsomLpghrSPAB30MQE3G1PHvVfrB5U+QcIYyYDyX3Q91QQv0Xvs4mdyEzOs
fxiexp9pf2YknlIOlvOU4dQu8v8yJnYf6TAcV87oUJCkd2PgqSknDRbAwstQSoDLduLK6icUJKhw
ISQlpeqZvjk8NVTUJ+JO9aNarCE0DFpVD8zuNRX7o6XKe1sI5ufTmlQyxDIqFfxXmvEG7reiIRC2
2M/soiWNMlgCJviQXH1nwstY2nYg6FxmHB97hahW4Da8OtUNx2BgPC9Q+Ya5JMgzd1wdCdZYXAXP
DM3+VUf53RNC0kYEMk82KZfZsX5aUSOTlLGCJjrLhHnhdFHz9WjMcjBpAM9VJvEcGZsAytBrapNY
LyYAQ1wSHp/UBj0MacUoqss6cn8phbdxvJsujZSw+XZp2b2zBe5kLU/0Ps5AVzImA5kLwUi+nEcT
aoPBe7SKpzeTNFZLq8DaaP6sT+w/tEhX5KVicY6DnuyIWoEx2+mA21Uvj83XmWoopnAWDaidYjvj
4RJPvu87dEaf/r3oq5CzMGji14feUnbJVkI80dZX8rxB29jC3j9wZSaPD4hrSKLccjp756EE06QR
Dm4bMERzF7yk9SLLrAl7iss0WAseEkW2aIiMXhZm2e6j+XYQjYbnvwG4abTIF4fLZNtW0fe208Ef
p9h5oCjzUnN5fKAwnL1Ghwh4vykNz7ZgSBuCUGA4QdwX46CL9NBE6Hy9GnwgBvfWD26pRYxJ7zT5
XaYSLYnAwb+WftbE1baDloCwqh4YBeVUzwnGmZaBhUeK6ZHTsi2Ub4SLbah1iS47ebcbm5rtWgpG
+h09qcMhg6fMeoz3YN3NjcQ/bhLLSmidEXgYjQvo1M1tMX8IXgUCbFTSYzY5hPTvy51poKvjlrVV
I7ij33A6H4Rp37m5MKDvAT181GKOzjA6gRKhrhNyRUio39w8bSsbdZFvg9fphyyEb2KYdzMXH8ky
1wn2mJtgyJVxqZvNcjqa1gyn3rK0wVABda1vKPtHITcoPbwJek0MigtBC2AJmN44dzsxJZsjiMUN
eS7GdGayBe8T5Gg7cHt1f0GvHax8KVCMM/oGoCtklbeX434WYCT58364GbEQwLcUY9haBP581rw2
tu4eX1rQ6xlNiJ5SWgICDa6rjOwSmBm+cfU9uek+YB+aWIk9KBzoJJI6cJC57nI1YkAzsGlY0ytC
Bw4gQU9Rs6afWuJwzk5IF62zNXm8ukBYmT2S8FQKsUBy0gKPnWjRU9qTe1TgRPp1anc/Yv8FIgSJ
Rf1Ks21FiD/lKKfmpdjE94ZdSiN29IAZXAeqI1M12oiPL173VwtqbQxpyfDYlv5IY5/k68gLR5aX
w84QcfpJ3xJhJbzlQc0Lja2V9Kp4SfOn5wb5x8/vbMU0PDz9BtJBqViyMl20oVaChzhZPMzyjjjQ
zr4OUFawAy+PK60Y19Jh6DwcpfL4257xZ7Q7gIqz+BLxPZREDk2sAHOyAPYSvK9enAECzLb4cH2i
1PJ/VRk0ekBm7AJ3XE8doDzqhIJ6GOD+HWDWt8V5acJOx//wa8x9RcFns92M4ZtHQydx8PXW5YkC
qDjl3hH24CGBxTvkmrar40A4/ZoHo+hJpiE9gzTeNSAtCEJ+WBXKR0cc+24xg8tnrscBKk/AmEQu
CAsrGiVUuUSTgupsu9OwgyTlg1y/JiQUCQDWz3ct76Xn/x4QkjWj2xBuADo47L4j1pJOVkRCIFmf
H3/jV+3GXQEmn0tMRzKr+9LVgA2APcpRHfb7GGdb8drfhzqqK9LUi9J9bIp9Qn9TJWB6J/BbGNIH
C0EnbFyxVYFn3cjrLWpA9zaezBQuUvPov/4EsJI5HTA5jj1R2BYv+Nwuj5qn7OdEl8b6M9IX1WNu
gWJpBUfzh8Blzd6igCKaQfi1QZUx0qJUXzzrhn7P9WFmNwuu+COpPZ0UPbMp9XpX/9lVfL80WMSV
V3079tTl1kRqSE1PVxKzAz63CdhUPganc5bS27s0uCuqverMvDb1YRmgpEMlxsewzAVC0RKeDOh0
pFPpf8GhMLCx+Eah85sW0SymqgWiWXjZdbVZwHPP9LZ5lr/jidg+19z+1z1+DsQppjRoy2TbZ8Pl
1Ws7BAW5xTZ5kQ8dgV3R4hy5i3OAWvuc+tikht/DtSU8zAgnWW5gsfzQ7FzCC3MZsPuINF6p9qMt
PaYRDC4QcElxtAmbwZSzmzpb3V6homH587SmIzi0+TbHRR0x09fwPtEZx/c5I0gJMgxlBil9bica
2VhIFMvL0+2IXLewKnRmMrWDsPr1KcRV9Hyln83DmOtcnfJ+evo0bW5lkOY8F15LV5BUJvaAWxhL
mHzNM6NWHRsoyXP3BueFjA93dtWiebRRWi7afqca34Kxqho5FjJomcNlAvsfGa8GkVFeYt71jcIR
tNMzWgBu6u6v/AFzqBFQWZjlHlGphV9O569dLBqIOoRWOncqVDfBuGzrTdtfJihKbTksfc0jATgt
zfpYGJwJ5yazIxuzkTYXmHlHS/jRSggK+zTo9qIPj0krOmmxXGF4kGCEHw88OoXs80VnXQLdaHkx
AvMUo1kOqlcCMtyHXoKbV7gHPpVnzESoxFO7/p+nalyLzZW7IXSl6MOxlIc27bo6P7aqmQMPt+f2
28GOAvRMy2Yf5ldIQg351LL4WbaGnvmX9D6V+N5d+MI+jCDzTJdfHdzJReyemIfn2nkOzBpDuCGS
I7DLYlW0BAVguvRHQ/JKj5v0drkL0p5fyEm9fXUAd3UHDbrW1cbTGU8rY7edx6834YDdsZqQuERi
Trqmv9LfZ1K77GuPFvAbUuMf9qrXCw/BrCgoOb7EtXSHxXlk0FoP2HZnCPeCbdPelF+/Nso2L+pI
WtxWZxRAy3mUmen4tAD1JRokak1YPYNBUGSDsq/C1QRvl6OnDKjzzrJwr5JnYApHj6EzL1oZNpsi
13XvY20bQoX8edSu5vXJq8/hDbaonEVB8/RftEwKtfsYbVLwSC8/+lgHo5QuUAEZWLNU3Zl4Z4Ut
gIOSe2G9Wz1GXvC1eA/i3HjerMPrYn66LOO+4zqLqvMmzHpXkKfc8FUxDDDT1AH/y+8VngudA5ei
jGXYuyAOa0CVNqoNKd3vVFk5X/wILUZrhhKfHNilHTz19KuVEZTOgt9qnpf7f8gb2KyO/uQxOX40
nqORx48fdurasNzfPgtEVGT0zJ/BT829odGcLKaWl8RKafiNKyE1f9t74M6xhskqsVodishnz71m
rhNTNBj0Ga9C8fy2VJ6TMLpbZFJHKon6bQPRGV3Snxd1enREXHDtgrGy6ZkVp3zI5NXZf1nbG+QF
m3fY9nVZ2mk8NRSNsML2GGlgdEuaVcHuOyV/pFrd8NsMH5gTN5VcozILaw9F2TyyM6n5pXFz6uX9
o0KpRRRTnfVEk0zRlPdm2S9lUI0zvXiWr3iHeqauFEAueyRzxwzIMzw4Kl7Ba8jBExlZ+ecQlszp
TLYwFVqVD+Ss8AG9npnfB0vrwT/7n3BD2+4627dij9bEDpFq/yzGxelapA2UvH4IpoqNQLL+nlvC
EAMl5AqMnT8GCgE8AWyoyzUMrUeWEMzS5iyL/QtsvUbvH/yBbFV4l7dN2dXSalEADHZxQ84q+I3/
HEj4tKs6prNphcg0w9fVkLKtplEHDXALA9Thqkead73xPoO5sxr0M+6c++pa1V+mq0GFyGNykBHC
3yIGYfiZj34mxZqTdTbCx7e0eouKOyn/HnCipZWAEmYDnHaTCB0cREcKwRRduAIDbU3fkKognFNU
+hOnUMc6IMDsGj4ZcSbHNk5YRAV2OgQrtf0rYeXi+Jx5PSlvg2Hqp9a7x+ccHTfGhtYiRWUBGw8t
1FQKZpLPYVP3zsLFKoHIk2hGWTGXdvuqW5AwWKzcBtAX6i9KSm5Dm7z4Y7QAQaQSkP1+Q9tyHhwt
eT9eFZkIFhPDIGLshXXeQPh/QCOVOA71WEjfgU1TrLNH3jrBpjp58OwUY5AZo9nfNH+CNBe1zUVL
3QGef3+a4WaAP8QPJL98XpO7GY4jgAA1aCyFIiBiufB5slWtGNkQR1t53DWg67fT5EnHUMO4U0G1
SAX9nIw4c2e1NC1T+inZaA6HGY37yU2UKESDaU5WipONYgCXjlfZfXafVi8kn9EmV8tChkdYoCmq
w4NEKDT9is302yQpZFBwjrc9wyB4T97LQIqP3HCuCCp8KZfAySJHXYIHbtyBjOZhkoAUr/jo6RnQ
Bd0+Wdmnso7HO1Ymh7YcULp1n9n2fzbo9u9AogMXcBBlTN47YonaC5JnrhoIKh/VoDUqR7A3BoRD
oyWnvPofBTSg6YH4Ff1sYhAxpZ9PFY5N1tmJ7tIXIqft99I418UxLtkC5eeFgQuseHIonYZMaLII
IhFYcwNmq6oZmwFqwm8GJGyOL6Wl9uPrjb7V/pFHZfuhB9+BL6WC7ksgsY/TFVNR2PqfM+HbrIlK
ULmtZSrTcqsNeuTNJmOT13OxICWqP+V1ZcbvhmrdUiu5Nh5A7SnywjLG0GWLidWY66LosTXepvJA
EKFx+yYnLlFflJQTYTfIVtwZOZ0xs/yECuc9m74Z3j/PhtP7IhupDCNkAeqcWsZnmglpjNdE4NEZ
w4OcSbskhI29quU61BtAcxqNOBvmLjjaW3VqlA2jpQgmzNWjxy+bMooJOrM2XL94WDMjH9QR5mO+
jeLM2s0aXsv7oLWANBZesVV1vy0fupQFUc72lAD1WKpydWrsq7zkHrfruLUkLwbdRlydtLaoqhRc
z+SzFKAEuJXI3u/sjBVcak060w/JNmesEd3h+wPVJq4C60iqr+y57PwQytj0VQ5trBojNyYa2GUa
Zx7zQcSB1+dE3lZ9yUNdve78Ncq/2Y4dFjgag2RszFPX9QbinYnSQnn6vVXHNWEEUlqXwzsiIuhS
0z6krM35To0Rfw6EGzeVsylbyA5BbXgZoq6t2/a9gPn6KlcNVf7xlQy8QlumYOZ1RZqOz5vomlge
AiJ+XvJMLXxVfsNyEsVqzZd9RnShbKL+zJt333LRp2wrTwpj2IUEFH2VFqBDuf8tLlLoyurzw2IV
9H6PGL4olJdUTko+mJ8gKExDXCaM1umPMyTFnlV/WHXIP+Mglt/XkMYFLyc0vtEvArx7urjbUror
/EkGNJX7sLVLwOZvSmNANbv5qf6+ZaGPXjKVytEUUowtRfdze5W8ZSCg7jJORrUCDBrDJnfIBz7h
fAAyaguL1OKzMw283F3NtexkaXHdCjWd+6eab+48EC8oMqW778ojbU25gpBmfbE0BllAdfIEsThU
efO48qQiGOYrSZK0aukcjK3PMNjz1LyCKDnvTod454VJ3hfUYbaUL+iSD9uDN+BCFPnKa0zDh529
SnmgpEwyGSL81v2kWuzJI2C7G4EMQCnUOLVsbKKtJX20iFYWnwlDc0RCzpyw/8n4tJzYEXbGhc6z
DAZsx8N5jcW8bk95CAvAf2WkEWXmd0p939xIh7CoRrZnp4pUqmNRNOr7Nx6bnntsh7OLtmcf8WUf
8IVyQfPufvWN+E1YPO1c7BJaqzcn6URvXCv9FXS2fEvC6aE4AGWHYgRBAw17y+5hZvB+ehm58/ps
SQHEoiwrLfkoqnPoX8SJyRQTi9ralcyRC/yZPbQqlaKQ2muNEAf3o0OIqnRm0qum9Yz4nrs3D408
bsPR0hXxgi6Q6qilYixQ+RuEEUJqan9r2wQN5VNitoDMBKW+RkxrFB0nZLG+iwvHAJRriJ8GqcnC
puyNBE2HrXOxznEVz+B2/i3gxr9wKDhwXMHmTm5RN783k/EGxrH3d4O7eSYhPr+l4qTBSno3Odgi
zdQJWVVCFVHuJ9vxRG1xhgNtX3lFEjI2I5lDOonMRtfwuev0Xni4O+ILbsS2tlQa6P/hqhUvjyed
JFUuMO0PNrwoL97WFWAWQu0IGh3w2wPMbvj0WLkOJ9Cjh0E4+J0ABl34j3PdsAK1IZB6Ja7MliMl
kEsRnrMgWimaxebjWPOCUwSgF9iIaWnUAo622SyWWpesQ8h4znrzIPWnB59/StoOAppL3V95Qlii
qqZe63oRnHPWH1zoRvloLYcCnwi3wN16NASGz80GH38iR28olnrP8ia0eFrcrh63N9Vp54SzNbMu
LDn+AULOXEZKoJMDyaSJ18Nehk623T7EVwhLyD1vNsxQPYZ9bxNmm80naDLgS2b0hO74FNBG/kp8
Jmugl/M1qXHrwBxjcUH788/iVG6RItzD3+jiuxcnal7bL0uu8LCVLAzMRHwQdFPSgIeh/02Xh9xM
aX0+g4uj4g4ngRJwKgZfxeDha4M+5zGhHQ1JRJH7pRyRpXiaSonjaJF48VTlzHNvyNNPWzEEja7S
xiBlUiPyJcfCUfPtgdf0iYx4grZYZmGHTM6uS3hbzCpC7meDJfoTQO/bggYll1gM1NSPt4gSb1k5
WddI1cj3iKK/AwHk7Y+X2FBGedKCHvq/5J69ntHAUojLXpLvL11w6vqPWt5In665l/2oDoScEvrq
6XZWWrphNyUNTqytGLUzoyFdz9UhYcb1xrWAcwrs6t1g/moEjf4/wflJDq7S6sY2f9Q52+smOeWn
chATnAsEsu2xxQfJoZrHVaD85lSoC1m18VrUnUp0D6E7uIQeLze/nGObVP85fyh4ALLVg9IrI0f5
J8kddEOZQI48AtwQV1LNFClz0vLuOp8IYpGpZtQQwA3fkKZP67nHWj00koM4hgVXVBj5EhyqaSAl
5cZETA/eX90oWponeJDyDAAxyo0r0jSI4UtaLrPnTLvT0g/H1G9nXafTCEyxGqhGjrpDGlMbyMr3
fgtf3++eY2Oj8TMA8N6qmr/Kkx0FsTl1WXfIFgJU8tR95CqV8nbfFdrC6+4e6hsBlQAK2TOvSTQ5
Zd/VCkyBy+UsqJ7vnFPLlnX5LBjNQjEXaQdXtChJEyYMBdJaEb7uPZqiEYyj+HCc75Gghf9JWexu
leS8Z1f/5/zSCaiUSNHVGHz3xjn98u49wOFy2zz3foHJp/xIqimv6ZrjkluRhkhMh/wDcnE5ghS4
wNgiofd3Tee2q9A4eJcPjlnrf6sbzfKySPDRK9oIK1WUzSLChkXsXY6ErDgVFc960MWyemKDayvB
/9n2kX962kuq/VwM360ezvSHBc3uTs2wSqOtVIf4dNs2hyvfXHKsuQ2ZnfyROxwPP7ckfcbcbLb8
11UVB5NEZtRR4FNzqyjvZ/+1djQrNT0R6D71zOs2FM341v2Ma8gik9KzydCWOjcTP8bZefOxuDLg
SYjjMOeA5OXZEm8YbP+ZQkg/hB/iTJyoH5gs5AmzKm8cv//JgjqdpX/EOVeU++2bLZ+XDzrDQm/r
kGVDSUenqSxmpQHbpfllwy273kWXYyx86828V1mnikHheuDdC99HrjeKh2ey24ywFxQ5G5BPsmRb
5Hta8ckTFwbvJ8fhckjAgN2l40sieLz7ggWhEgB52rBRqhYrWyYN6gfyLYxzEeVMc8C7PTLhNCI+
IBU8A7PR0fO6J+5hP0DwRN1oVyQJs0vl8uwmtM3D8I6lcux7TltURaIcTYJGSlvWSe6C+Y6QO80B
yF5GB/GAJIHYBcP/aXsR9DJzQ/Tr1gwqmO6pIGkCOqNNSlmU/Er+mJTU4lxGrx2uZWm0g55PaDG6
fLK0Tz9tKr7P2LRv5kI2/NkoX1i5X2/dIpvyW7Nda5R/SqaTInZ/ABN4pMX3oWGKlErnvdMi0N+g
tpQaTuAoHDWsE2+9ewDUrhAx3yb1HPusRBJsht6UtVXB/+BKLaocsmHFqhanqbk9mYa2gl08yyy8
EZ0fjwZnZfqYSFnecv9ZQTRRd/STqfD5CejTmVrKMkYEp7KtvdXsx92ZthMGcpfMl0fEImItm3jx
ZNAwq8FcEyw+paF1M0g+4BMG/yY7jm38jdpRLLlGUco+gJBfoLIq2QHNU2HOVkhCAMZTcI4E+Tql
AykYEKJZtdHbHdFxIYBg+vDQrUXffEYgSgN86y9Ga9GU3yBe1+7uXb4SnVVVgJ+y7+4U/Ns7T9BF
Gj9YmW7+sApke8v8WFEbNxXDBs+ZEhrli5dxG/q65TEXIKrKAoGm6gbH3FdDixCx41DWPEuFKTrs
GTHxtXM9w41w5b8+hZ7z58U61kpMXcRkrPhBUVj+3N6FJ4USx5YiTSnhLsmSsOBRV2znL4uJzjDe
fWizcPGz6Vdgh0A2A4o0k5BCqnizXtSxce/r3OumbEYlRGIQzyBJpS65cIIb9jCgNthY4X+4YHlz
wmI06rI6PyTLgr9h2ca7WNRrEaQgDrmj6bEh/aw4tO1ELQOGfZ9Di49m0LEFAPiRJ6yGkfSG7t6K
3gtXWjDi8GfAhZpR7ACOaHfv9fWXkOSFlMZM7Hhgys+QwzsAjMxVy18Ud/wFMuOTpakKQBH2+3An
cPSGJ9qpt+ksiVZpGkJ9IHvOoxEjAHB7pkJiS8bmymwola+KLJ/uIWZrmFvvBVIAkSL6C4Axq0Kn
IH0hVp+ETcO2TQkChV1/4d6rvyPQHyMX2XhIQgE2e4kG374+tAl6f6he0kZJm8WSrvQkhWwed30n
almjOHAqIsP4LHbamRaC47+6GfNAU1LDmkjNby0JiELwN3gZWLYbUA/ZC4v+jTfL9EaWtGxKyr0a
5mXjeNDpyqZknqL2DOU1D0DwdoU+W25eVgXLbXRFPKMWFXKJCzaEfwy1tRCEML9/xhWl1ZJwzfCr
aynp/nKvuGb0Tauw6MZnpf6ABnfTw5Jk623Z22ZHmZRLlU1UPVh0LHQC4bR+qaPeq7jPX9X+/ITw
XwIW6k6rFLsbnGtQmC7H68BSbpX43/Ec/hLB5TVvE4SvDCJgrfInP9jNqGoSLccNIhypjxzjXFB4
KnmvLSmvZF8HgiWZh/LiHNWovreFzFRWPNwsI9/oY02jdwxlaAtqL0CygG5nM1oDlRNL/Ie6GB7B
GcNTs9UKlHH3DPN9EiRT6tjMxoKFSv45nYJotdKCBu0oM/aOHxwcGi9kj49dLU94Sp5DwNp2s4DL
kOY3bKYgqODEGsgjPh0oYDLBHKZO88a1B6rUS07QQ4Ou+5V5EzuWulurlOj+fmyRdoS6UVBBTJC5
Zo2Q+fPScMenwJc8RnWvx2WRbWGDzSZZ4mCskLtI8eK4YYmOkdjgN3CSgQHvyC5bVDPqhJthd0Ul
DS1gGwLv90jTzxnRcjwDN6ndVvnflm7OFaz/p0KiB517zb2GkqX3sIKZzQkjKKSfhG3PFds2MR06
7fO8cKYD+ZuWghXTBL93fYl0zn/H6lu3NyuDuNyLrQrErNzqwR+3ENXnezHPh1wJUhc9UBxsebB3
e1WJhYTizxCepdoVWEsj8FBZROBgWsjHMbBNmNKI10JdBqeKWwEou0bW/jCTBjEhjSnpSuELP7QS
pAc2+msVUDOQCbQ03VFRpasNP1wpIRCPVB7uXVLew0HJqmL7+6TaON9v0zc+DSVxiEYAIkAE7loQ
M9Ck/DwDoi8SxSJPUtT6BsOYh28n4h2YTWNEf8L7wknIQ+ZJYdzfppGoJSjOA+xtilvV6cJG/90J
tUuBLCpm4jtCyyMRKXSnbFrmZT+e75lljUsINRvyxHojATbfgWB4/YFL/unw0Mj11xTi+XFewO0f
WvVtVgBvbH/gkJn4LVqGN6llvrjx7bZmnj9mbRruT9+q/qF0/siSEpTQ1+sy81jdtwlso+fc3yrv
aWaCaP0iLxw6tpN1WAfey2zvusl3PQ/h8ifOlfPeVA5rokCcPOmYoml+uhGgJGTcpb9yNS2pknOM
nXIYKsUPJ2v5L4PQ0wXPthFyeLWbHTBt6tRCLsy7jQwbofQylarVxRrG6iRT3FCLZOo0KekccCjU
OO/MxvJRFRIlTOsFxYRc2zRoQaFPi8ONsPUFIggZh80njGXeNb9Cc1jdj0amVO9Ka7ryLNDsp1Qa
UrH/58qe5kSnCghvDtQe5uKCHCOmGdoPeO1U9LSou7W9JI2Y21vxQCtuqnobWfivJywU7j13+WyD
F/vG/0FYVt7uo84drMvX8MR93WMRo3rbhvx5HI6VYApzHiPjHRNzMoGhIlGaOCYZS2eWWz5i5+9F
tGZxYhdsVWz+oj+YtKSVarylcocQMqDwGkTYktgsPqg5tK5lzM10CX5LbCps6Fc1moWZpA1HTXmg
s0AvCRteAJ8eruuRh0aZbdxNhwfpu5etBShQ/7FQFM7XWMycs9FhStXMVuu5EjWIqrZjKstRuttF
KOL4eByC/8oyDG/53/R10SmnnBFH6z+eLiTLXfkpNUC4E+I6LmfYTCkaou63TnxN+XHPjUSPFd87
g/3OuZAhaBfKq4DDBAD16GicDhKGSXQWmERDNKIbcQTNsh/AjcLylsOUaa//VI0NEuLW2DB8sQ+J
gpWYf6viorcJpjUjW/mXUOinILaLmNkzcoIxtMr5wysxwRChUe0nLYvd9it4wtnFJHytcOFtjh51
VdnumUk2DUY1CWNb7bprHnOPG4fod01UeRQaGIehUx/JvAjW3JOruASA0g6DiAeNwULd1tZrlQdS
AjWhCCrtRL9Hx7rjX6GPgv6qKR64FuNIA4JK5s1D4oocuKXNHuvOwHXnki8vS7bLlY8ci0li79WF
FBQxLRuXKKH3k+oV7WVfFLlnoZ/H25b4C31PU3qmjCDLvwLosZnODd5qrETGrE2lw5vuabMNqKf4
mow/jbYhsaQ2MIsBVpTyIWECsr3NNUuNFANFx08N7no6SC0dznXbCHtKr7bQAhOvUgO6XernX5do
X6BT1yPnfWAFMxAV3xqzqyqRo4j2jQiIpf7SlOL1PKpH5oT9n8iArzuqL8fgkQrsi5Q1jLggwu7i
OIRNvh8ud9HADdmetBSR9N9hoEavs4pNXjcAGKmQbIzv0ao7z0bjZjcfqjlbI6KlQucfc4SRDvyv
NUv87yuh5qOvUDhy7+Cf5IzoYIIpM2yz2DVDBzF7B9m/wnNwB0MJnRFCi0JR4Wc+h4Bsim5KktAF
zzHdCvkgsYUWf99pfk0LktksRlez1TsIdGbQgxlvj6LILnD+nvNREPrx7oAk8c/hD75y7j91JQZE
l2imyykErgXj2lGCZ2yDiRhw6+S6mvJh4ahlBP5m8RJi70DHQUvkzRONy4oYFjJRaXWnU8PqbHbE
tkmpe9SRYhGwyyszM/vJbIYUNsDhXAiWUbwSNwdL
`pragma protect end_protected
