
module SimpleClock (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
