// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QntfCXl/rmgEuR08vbaGe59e6blW0oUsRWHl699WuYkRDsEb+BjQmrSxan9SuTcB
H3iSrIirK2GZAVwjyOzLjdc3Q23NL8xuhsD5vODfIJreKS7MzjP4PsF5Bxz9xU1H
NKwmfZKlwsOnJxNhICWXTtyGAizUleh2Mq+Tuu4IjCo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5328)
uj52VtztmU/57YQvAj6TH4BTaJlyXUFpv8YYwKbP7uWSCYIz/3RMuf7fP0t7QLJU
VuaZwgRLDdohob9OK6A3OlaKiulwrJuVY2D583xzkNoppysHOW53OugoDwNCj26+
zhU0XDYZRQHJ2/puOoX423FppHaAGXqEW/CzV51VMjn8qBX+lPHNk7nWkyHVfWQv
Mj5m1jsgaZlxo0lMwzgFIUbHhhkhjJgka7So9HOakjLmhAItOEgdrLAqVu7L49uM
WEtuU4iSiCSoMPOBTlPUi1sgGt0ChbLs5IU5ws1YdjaCaCG7f5u/3lpDeHKTh3A0
6psPvfOkZ7YTGsbHYSQNXOV27+e1Ott/rKeYlJ9TACjDs4SDiG7dHblITsp4j2RL
tN8g/skfPm4uOv32CvWyFjouG4YIfrpT6GpbSt3vrcGMl+TzzMSaAQMDdIuqG+dZ
ecdd76mnHdLcmUFtnGn86D+sGBEW4FwTi2YVnQZ6U/4xxppNfpZeAuiuUdyQXO3a
VQIE33kupsc8HOEww6zsIuY3/LZIr7HZmOh27wrwSw1OAvbnhQw82jasg1SZwfDl
qa3jkpA9S9GohoNdqhJ9PGRHeIAkVoCMmjdeIgrRwhXKvIzEZ1IRZWhlxIPZl2Zq
L/hnREVgMdxCC/LqheInO+fEwwCneOv4yFfSQlhtS5J4JqAbeYMyxJAPejNEPq+8
cmMdD1RMAZXwkD43bqoKQJ0c7gbUM8xoyegv4N9hj08TPhH+nIul7E5+5slXVJth
Yqw+hxcmZZGJeQyVht4DrJXa5KlFYiLmCzWrBbRT/8iUKMvutn89SFbIZFaQ0t1Q
X7DQSePX259DDY3l2FPgODALVTGuNqNJtUWoSQH/NZiP0aJc5qErNw42N2T++xtK
JnjyJjBp/02dcLsB9ATyyzFj7mFeFZQVEPEhl9fVes/5JvemWqB7hkJLyrsFFuWg
rBM9hDZFc8vvOQDbOPMe/XkBJOv9bNaCGuezFhubPgY+4tJkZeDZWksPdkGRI7N0
d0WVy72RD6AkSb2dh9nrGxKAUFFHh/wrv6m9IB61HrDolXMJe+FDkSB+o/qrBnDt
ToFpZrUhui3h0a2JYMcdUdWQTuWlR7ckANehCvU6+FqKSpg/h6ubLlsvGDTGseID
EEV+9ikUDVWFxa8+Fm5B2SXVGh24GfxLAkpP5H8MAIz/SVYWn6O3htDjuB6M0A/z
OKmrEIjYw7fvGm3LhpxjD9LeEXa1MKhTM1fgmWoI7GB2hu6H9SuV7sbdQt238GTf
id56rFOVK1HT4PX+RFzuXl99jqPB3cMVvSY5SF9WCKCQslbxIU7dsBLmGqNvd0FF
GSXF9ovLOzsmBOQfA2jtUYEwEKvBTillH+zIxDFrmWiK0WMIscmGF9T9NFxZwZ2U
3wlNH0K8m6GI18MvNp3H8t2aqa8+/7BkFv9d4kjwMXEfdgwyc/NlF18ThUqUPqES
aHQkxEDtI+1LJeCqvpG9Sbx7aLlGEON2RywsglW3xreGgezA+V6LHR0i01zUUpd2
QJD74El7Evff/77j2G1yOAhRG2fspZfUsvYAzgPKuExPubOJXuudV+5SQArmHWs5
EJYdFtOhGUjJ9GbFfqie3Zw2FcEjfoJJ3Oe9HdoinF+v5eKVz0QjckFHnsCdsPbo
HCKuCxAhTbmPZbn8cs8bbmtffhKOWP/XpgEDlTszA7wXD690hdolZGm1UOC5PeFy
DKjh2BZEh6S/AJ9Sh43SKt14jbVEbh997FZL6VhB9HtyYIRLjk5XQVeJpcg0Z37P
NrdRhSzOEZUqtFJNi/IPefn3qh0jVT+D098ivr2GodEfrgz7qCaRwcP1UCqaqsKE
igQFuabwouWxtOElQYfeHjGrK3S4H0pKbjPVGFBEel8nlr7cJaXrQuwi9NY/B4E8
ncb1f0PJMCwvNVwIPNyEh9duXLQ0K74gjJ9bzWqB+Y+cmXRoZqNhDbLPkYZPZyfi
ADZIK3tGrMIueuUJSyYpDjN3pGA8kD0fdQ7m5fhuiJlItqgYlp/Xz0qBJCyqNg5u
i7TbCQFJOHZ+jtw/+AmXplVHB8IbY8cW0CLB9UOEiXb1qfsuOxqvEPsSrZ246JQe
NuNxLq0lwS3mFZ2enNfdCtuwnNpCJFzJ2I6JZ2JjRmQaPzuFApZYjwJLySfjyfVe
gJkSRwd3Dn3Tutt6SQXQDrleNi8WdgGwUO8hyjCDOqHki2j/RhLJmCL94k/MrEpt
ZeQi9pKcPN83IsEw+ddd2wuetc56BA3KCI/vmXbxUIFxpGYIpgTcFvAwl3rvJhcs
NWQSWuWMf+MHPUy0W2TcnvA9wrP3oQFbKyURkXT6PGTU4rPPS1IT4Q9urG//7skB
ulk66wtMOdQxCk6yAGERqUfRTF3WODlJOcH4lfFKQN46IwMknGlVQjjjg3Qstkzz
BtIDu/PtE/XwprcpZYCrR47k7I5UnN8dwMFQSYDAQCjBOhBX9BB9seacAD0zbIt6
u2woGITwtDX1IGTgEECZUjzjzdF5RHW1dj/dh0EY0fZug5mDHMsSyOqj0YqScWto
0ppgbBE43nf4JYB4CQqI3oBKINuImPYRtLsCp3Wykbm6EFl+dZQ2mGzX8svrvKbg
viXZr/VvGbWhjOBy0z+AWtWRhFV1Y1HsGd7tKFmvpSVxsTOKxJFw7nsaONGMtwtc
M9Z4oMBckHACEt3eE3yL+jeOLb6V7eUFVQgfZFn7TabgDe18NiiYTB9JnpWVpbrZ
lJ2wr7SlXN0MwdNiRV4Ai8YoKNbjQObs2cPa2L71T/FYxz7Kp+F7lu1MnyjGedC7
fYd+A3cmZaQl78/Nyyq+Qqmc0xH3umE2LCwZvjO9I27uM6AUYLepkRM35jdg3CnV
WxiAmot5PLc+iIjQFBP5a2Qy2P8C2uSckVTB3GaNcW6ICH5HVkSymZeY22/fGyXc
idAIpf1DELrek/yuEDb8YIYDnH0Hs9xLH5uNVNEbnBBBy2gEPtxfAAzd0J1rOGWC
UZdZ0t5sX+Pyfwj/fTa9UnqNd7N1ZouwrHsie7RL97kHIRYsz7bweWJlbREV2JFE
YghN357ppACSiq0MHqrkbY4j1PyIGne5XXEU4dIFbvyOWYeuFnRHgP0pg4IThA/m
YTIBQra2yCJQgAGGmEQCnJbVzthwVY/rh0Qbm+NryFya6PUs3IXvzLTGKq8fwWe0
9dMYJKarR+7PFgo953kfZcsCOPjK+7NC99N+iwf6EPTn3CieJ90is+k3qISGQLbv
iQrJuNCouueuUhatnEfGE2s+j5a9B9U7Xb5dGoOSCJYOOWvkm/Ydm+EL6Oyrlh0q
JrGpJwM2PqIPUL8y57paGO+VIrAybH8KpsIXrSp+9E0EK80LB+xjhLkv/AJvxUqq
RJetlWFTVQuqVqGbDL1bOaXVnUB9pwVvxbr4QIHejmh+37Y2WU+dbUXH7+lIrl2O
e6vlLIaca124OZGsYsql/0/1FSzqUK+XhlYWzcDQPXWRtBHo4Q0kyfOF8NnTeadu
65Ok0KZkaQZstMkHYU7/ngUyzVb8hy+HjU2C54lkEVKD4dHsdCmp0Z29k1jlpqYf
PSaukyOQTkFkvGNPLo3NWYQu1Jphc+58fSNT3+lOayoOqvbu3ZGos80SeQ4G1Len
Hj1DFMzMkLozBtP6YkiC80RZS4wTpoCMt/YNhShx/+PvYwvE/Sjmy5bjY0Q5+DEH
wIwqU6/wu1eA2E/vEQ0NvGI56cR3Nd1fj7HGg4MVETLtqzurt4c5axiX8QSJPT5d
uCklghUo7FJ7bu4R5lJhoQW8Zw2fzyhpzIrnhlCs9wjVN2LA8G/UzRDsiUFs5+g3
W88ctEkaRdMNEPo2vB0v422cgRtVLjw7++1HQbaG25Sel6xeWD9pgFLWkir8vDBd
5OkaSEDiuMYOxzeCbNaPaVbXrRszy6TtzKI2HQww6URtynUI3Sil2N9Oi/d8lsNC
jRDt2NOCw0jfAr2qfj3iWF2y3pBpYsV8/AY2tSUGGm/eN6H6fFtLv4cLiBZ+OuQh
VFs2IKUmO+2g70xPCLu/H7yu5V2M9UOtFZJ6zPS4TBiv+QGB3+zOhUtmpBQ5FfH9
vuDYbeHmK/OpROEMN9Eb3Lu1RfmJ+oWo93OG9TGoqWXuTxZioQ64pNKkPhhsFYQc
8cfWZhyItvp5yDqEmZKeu8EvqlOSbxINC8cnRWlCmHOJOv+8JZkWSyih/AnLmKyy
DSji38N6DTn7K0e2m/pIyVdc9pIUjDYZEP1YUNmKBn60I6t04IZxnKruufnvQzQ+
vcdoHPXmH+Ji8ZfmVtPGw0pQTEI4KsnNWgZx/3JQHIuNHMEOgnw9yvg+ZTwW3FJD
0dy+qoGVrpupn5Kk2TDvC2zfcVsWG+bEJxsu1Ucogzsaeoqeye3ofr6i7Rymf0oy
rW1fZkZ1mhyLZU5ZndT2bkWBxhqqmtP8FXYUs3eVMB2MqExHaTzCDgaFh67k8ckH
GcT6rsWF2SS0uSXLOIVYTAYQBC/8+sqPHXHXat78h2y+0LIm73Pz7rFVkVVyQbcL
o68p59QQzn8b+DZ716iZaHWSxqdTI1J9EXgLXVv9kVpgG7vHLobbb19yFgmsmly7
vRM0ncbq4le5JDL3UFqPY/hLSHDWGAvR1SDloutnmpJNerhG5VokVddC1SaDqyG+
zzV+F2B1ISN2TQcNXgDKiXjGSERr2eT0UzRvZ4Dky+AVqL5v7LZMHOMHIf2PsqH6
djBSiwHMs6/iiLUNacikcrY8h2nAIYUQlGGQPOjhw2YCRQU+0UArGVYph8tlCf6H
Cuivws0wNi/qf4ijYturpkoj8Rtrl6CeIUK6xtKIBlAVwWDKSXvPYOxMZjZUvy2R
h9lsgJ+A3yP1zkAJ0GDSuc6MAXR+Sw2dBQwzByJWtmwmYCcfjpAhxHfFqnaejQ2Q
N4cvzzxBt7Wt48dsznHiIhNLol7s+wdf3UTYGeY2u+ZesLIXwvNMz/zUMW1i6ybW
XCGoF8mwhLtjcHzR9i+OdHGjF53muxW2HPGK5MrOXzKOvzkRI98D1T+jTOceyle5
hra1Uck47YJVT/6sLxaar5ij58fCejKejPFIpvBlnPQeyiwUaUUXKaLiC6uVuaOU
Slq3BUnbplhrllJljtnvdGQjLOj5XuPOIzOjWsXKD5K68eCqIwX6F46uMT4ItK+Z
rifhbGAbJD+YAUFz5RWD/4mgiuyr1DzN+BbgXIlaCf3F+30z0OSQw3pDguH3z6J1
LNctkMZ746Jacu4OdpZawPPv0B9QAFKz+hxr7xUenvHBPDithsrPFbm+uZzjyGnI
8plcEL9EhOh5TI3dNaEhiKqfpQ5SusjG+vHBnVRRAtsb1pJw6T4m89VKqPsLcEE8
UuZ72alTV3F+ihHHW4ireh08UmuKizcE/eXHDEmzO+SlHBicbCxMR5K2B5XsmrMF
FyjamDX6kUXSV9fnSmSNn0t97O3TL2VydviZ1ctvHvC5O3hAVaAw41VspuP3nxv7
fgd+64s14ygu/YVrTnXTTueY9TkCc1+iu7+1mcrli62IZ5rTrOeUGQKcZQ1kxmmM
EPWIC0YseMBXVdAG46SSbxRczsiNzchFPsbOgAwhHfM5vnmbzyb11soimd+JFZ8v
5UOhCrfqLG5Sk12JL0351/6m9Krdl6dYw8+1JYSCpu/5QiAzMXQMH+2laDKenDGG
5VxzAraBA9DkF9N8zd3pD87jaksP4a6cxV1zzh7sZQfG2Bot26XuRNeDVIlFS4Ze
enbWsg7s70LAXg8nick96A+SVTzdNYUqHVgeZHIsIiVK0nJDCNulC2xBu9JRZsoz
YoaJyBuRDe0el2QPROYnOjT9dr2JH2DL7b/PiNlRK5EcJxkrfeGRp/6m7q2tqnML
vekcoe4JSHRC6SEfSkjhD5CHLq5XmxcGtADs7eFt64Rx8uNT2NznV7q8BGhwQr7m
mOLERMC7VklF908JXqgbwcZmyPCAxCT01NaqwXieSyRfh0zHWF7tOj+w3IFtF+tr
Nd4huWnd9Ut6QGRrQxiMSmvcybl3StzOlsTBQxDvRC86B/YWu/DLezxVRyyh6O0q
xD5DzG+YbJ+OTbrNKBPNCs0q/ywWPtm242h35/DkXjUnAPuTPvjR1kZ9EUbPh47E
Ntg8uXewpd+pte8AMK0+3//FOBflg9CoaIbbMVBh7dM823az2Et/jtoUoVu8nNW6
a8g3GvB/JXvJl4ruIReW6C9C7ORqAeu1xzbg4VVf9xreMzsX4A6Jjf3Funn3aJH8
75PV3UhLmutsxoG3vfOSk5a1XBH/+Thh9lR1D/OixA/hAhlCS/oWJH46CC7FmXYP
CzW8k0nwUP8zNgoT+7vObxRi5QDhuVH5qWGTD3n/tcBur34auj79yYL2I2aGGB8W
Few53KXwxGTd+/2EIER8n/PTagxbsUuIdWosG4n82frDUSrxXZ/GijpH/P+7wQDh
J4XmRzmvz+AkYiehbbPSJ33YEe5F+0pUfiuU8s1KtGdqGzq+jnjOV3BWU3iP7ZoR
M8i4TN0G74MWeL61TD6E1dSQfT5lqNwyk3oSJUULK5gM2dv3iJk2CL/6mGF41PF9
/pEuupuh3ZiHx6iqLs9/In4M75Gj6L0yaAv1/XuIHc68XK+BrCC3flc9LijdwWa2
0TycWaQDuXclchCIQq8XZDn1sCDxpmWiwjJ+gzoPkvPQf6+nlMvU/tc/zofiMBSk
Sq/3uAdXSC8hrcaCLXjicmhQkqBBj7GlWzBmVgoqsga7Cevy6aCYXA60O2L4g9Ri
5xBW1LisxtMc2NkQTjOQxzx/OXS7W3/tsxX3SdhGkZTsy0zXM7LOHn1dFj/zTs6Z
4PGRPzHpdX9uWQ4d/8hP9B7RXu9/vVDcbkJF3EcjUyk3EfDe5ejgNrS+L4m3sJIH
peAgVQLgYm9P6WLVqnIVsenzbRVbsMEmV9CEdxuxDUc6vz8djEi8LZaCsgLhsXwh
OW5DjJcEHAMtNDOYHvjIcUvpDrAuEM12Ch1LHtkR0mHTwXWxetVDkODFuMaTlPAl
sxL3/xeJCubt2lRmNik+pLeneYkQn4Av0y0dBVTVp/cGxQLioDiLecWoW2oL0gqu
`pragma protect end_protected
