// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A+a7obd4/VPjPqkuS5NbqTDl0fdKrzfNTss5ISG4FxEKOdVw9gG9MF01ooAonbGy
632Dmw2A03LotpLXDyPAbR/oBNO/M+38iOt4bJ+PboYDaJi1cHAIn6O5v2lm8kvW
DIGOqKyv5D6CxoxsdiUDJLv9CA/hrMgU6FbF69nLMW0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27680)
SCa2nPgwedWDLE7p+C05PgkRyvkBsu1Xc/spmViN7JRNsHQLf7kEwMXuVqajvzUD
iGPs1wVrdC1CblGSYw0v0iUrp14u1ODCRmCcMX7NC2Kjqtl4CMDb5rV0qd+k9DSd
wAxbAf45ezg54MITQgbSXnmMdNzRHXjRjEvhPY25MPZW0URPEOBQmm0IXfMTlre7
tp4FCDrYBF/VKcj04K3q+Q/R15SgGcxieMh0vXiQ4OeF2dJSq3hXSg7RSY+Z6HHJ
ImdISQj8c2Lvv6dF+rHBUtQsqJyjX6lh3BokWXVAwNIGzscWZjw7/6GtDr5t1169
Mpeg3CPzAnSFtN5bIwmbhdWkkDoPzDK1DxIjo8Z8LHaTSRiGRaKA/dTtgDkvyzke
k+Ib01MUQ6fBgWDDBss9ux/QvN0oA9qm1jpBdcWCZLmeQ/pvJGesEVUjCbnn+e25
Afj/dXLp34oAeV3zfMiSOxeVMlsQKLdngAiW2GLSybJ3OfEOuwhxuAZoT4M7Wiv9
uhjuIolbcmyACAoMtFvVvKvK6XlJZ7A70+jWXJWoOAPgdOjHsfvZwMK/T+ah7krU
mxZrYMzSPJzbNaXouSq+c5Rveruhj6Cklc2kUtCtDiE6elKYNk7N+/fL8+gqFxRv
C0NEgky3UL+3HGxRIJ3Cuo3/p6kBpP6xgMVzH7NdpcBgt9wB9hFqXTwsqDtL7fnb
IbwwbO+lsuGrnhezHvAp2/Q7MXWtYWaPqkppEIwUfEs9KdahyYjg86EByWY4rnUZ
epYfYOs2CqqW2/I94taXIJu+F/DlhGMS30ORvWDh4UyDgRP6sI5sP9yyWzfRsgl7
8UjsBtl0SfFrbIEco47wAy0tbjjX3zH/qWjHPlWfHK/kED7RIEAhq8QeNjA2pDd9
ywwvKk1hlY/Idla6TofL6PcLKgwkrH9XXvnDYJiGSnW0t/BQHINV6NS9naQXhkml
UpEuP++1YgrGaIlKrxkVMIVlI9hcuNqrv+km6R6cgmW01fnWmXOeaoLbNBUXNBNz
Jy7ymr3SHAgypIFF4XMEz2gFGjeYcYyPruFiAOpEFu6Spu3t/A+D+AqqpWCf+e6V
yMP3JiFoEtubo1l/aEdrl1BD/jDsIJ9aCUD79xNSnxoVYHiktH3mcbOZaPhJCjKP
GVMzUZ301G91kHuy79dq5afF32oOvzjGH0HsH2baZy0o2D4uFMK06OwP3d1Xq+RW
CCQouoTaeDvQD8K/wfOPUZkBSRJTGXDXX9M0ByHejF+ApOT76COVIZHMb9QEppU9
CbVZkYbpFRIVrx7qWXJ/pBgCiragPOKYV3XO6rN+yCxlV+P+JKYezAWCm4yP1ARJ
6CgLQt7BpzURn/DfUfnoahNil9QzYu/NPOTrynUJJ5LSqVcLopJbO9aw0fCGZMFz
7aFTEeB7ZyhK0m0sBwMgu5wDSi8uAAVnpPegB6RHTiUjM1wSMGqy98NG1phG/Z7J
XEN0KG6Z9/9uxUAZMZ4DoQq7+5wimaX6ouDxnGo5YEKhodv9ICMenhScgAP93iIx
HO57paIhIZkS1bnjUts36cezbna9aABHvq+vD09wbAdcLOswpXonyvDdSIoOxu93
ozFR6E5NqhQlsW6FyXCYBzGrh5zrQrNt6Oak2zqqQaLjbBjIa5cjB6zDvnOc4jpM
4qMSYotjk40/nyRm0Cb8Qe9Fa9servLh1tEiSNbpBTTr7JJSJ2JcTc66vauPTEcA
PXm7C58jbI7afzylYQZ19TIobbyD6Qm0CWO0Vklm3L+wbVa4DZPBsMBHYk626LUP
Bh7+bvI1wtZTjvQPA3W4QxElY55U5SVxvN9lh2d4rpgtpK7NTc1d0uZ4T5TOSvVi
zwg3ISIy/xUBq3CcGFUE1lGjI52t2doe/cwV6GYgsrnAbWV/Xk8a109PS4FGdS2J
D2FOccGeVmDtizT2fs7FAoaQz5oXFy1lGdxKjYgy8Zb/AuwNYj5Uka6jAWReAEwv
lV3V7Cwbatjudq3bBoDcT/rM9OUxQcFSCnWa1Ulcin7ynR1SOLnBUqXryigrcERP
25zYudz27JxVgGrDUTrIhB8gLc0/IVVBKr5o8AIlmXGMZUCIoYMFPJVrA/pu5NsP
KQIV/y60KPonCtjiczNu0cVQuKpuIOmIo16b5LN66OwQn9xn/p3ALZqRoqyhdRWX
DzFN6D4xD7Os9u3qXwx/K0k5//8YdZuJ14nPgsFehiY8t9VDCN/MbbFdBjK/CDXu
62XZIoSXbtAUYKytRqStoN97vHxY6arogcg+x519LsUqHQjdABJfnCkdctkHGtw3
Q4UyO/t0eH10/9RMrFyS9f7a/S6XzM18uG+FHw+ipfQkL7mTX2bLXSDMqyiTXGv4
OgHsvmIPS0+QvsDRu2cNi0XHmEIsy6Lxy3TWm16bnfZ7J56h2h0E7fsxlpcNUSWS
dZT3KfUgJG1mRCBuxZ9odUFGc2n+P+dKw8QoD9wDAEdCirLehio5k3o7w/OtG34w
1//aqDRomnH1qqRDJcp3e8Lc3zS0+siMQRDxnAYT/SBRG7VFonZvs4jU0HpCtL+P
ibHoR3AznkYK1NGl/WVFUEpvcm1l7JZlFc7wBSm/k3kNsn6OOBQUXQiMhiD4FB+J
xOcxF/i1BWdtwq3+wKfedqTyAXF/JHcYGn0sMVQ/M3wiCZ7SDIzB1epAZws7we2H
kRfLRnN5+/mxpldgMq9oZZbXw2+XaF4skXOOd2WOI32TDVJxob54X7ahfnBNLG2Z
HJq5nxIMVcvNAq/mFuFdNK6lE6NSpFGNfu2Zbb/OfMytMD06DNT3bEk0Kp+A/z7A
3mroVQ5ogbPOUMebeTJd2xFdK8lVBW57DORMODQNixrgZ6oL8S+v7k15MJmIo9A9
sMBQICARGBYQ3WaGDPw0rvClgUMTujx1IfTufyilYwdFt7Vv+lASNzJQOJAAs0Ue
ntuXg6tY8f4Y75mmLYY1sA0t7A7qumfUQ6I2nTRn8Mhm43HH5rx6VZni/4u0pU8x
xurksnGrBb7iKKd65BgRz1N0MO4sJbnVF0mrdPctJDtZmLEr5t3g41T+lN29Dl7X
8Trefl5bF8oukIj/PTeN+k9cePZXFAQC0yBqTbfJjepJoYfEBX5mIH+6gqmB1k0E
xajK7SB5drMD/LIK2rOYFDUk818hk3TdyGWd56nYw9HwYyZdmxgkmlWlKb5iN/AU
aU5EColfI4QmtwtlmZOT4kXL/5prvi5rVCjeBEie2pcOIuL+LT5OzsJePc7q3u7Y
C5g5VIPjf6DeVEi188MV+01qhX2tCYVSIZJ4czsB/VoeSfXj3QlOaIGvqP7yCbZz
JyiSe1Q/Sd6RXjMEXQjoQTVnXcfP9XxozSfK+w5pB4aioVtbT8ZSLiME/T7wMoqs
296mppLxQ//1g5QnCR99qwOiJqiOqleKIP7zfLNz3B52PzV7cypB2O8BlB8PN9iB
9iFFwByhjjQdViILDaOnVmDTJhKaARqfXsmCu0LOANvVClB7hmDNier7//967Cmk
51EIRWr/+/mS/4pli8tJzGW8xIqz/84itPn9KkmGmr8sHJkcBeizvSnyn9flkkHR
+XOl3pSRQqMM3etIhZxTLgccoCE/yHMC6gtHIesPeR2LabM17oj0QpdWVmSZ0aWo
W4SJCv1iOTjbnjgmpBeHmKcCMYqZlHrgFTRd1PzDdmr0Zp3CZfRUmt8JzTmKDBJ5
SYNh7zqovkp2CVek/UrqjknBK0b8F7RqPKhVOFX3BR3kLtp4ITinKODNechkdWl4
7bdfn+ZDqSKc13wGaa1g/2Ety3p93uamGFrBdbTXaoluII+U4DPXgA5pTn4js7tk
KmHHpsM7ms2J0VV1KQ14L4wC2Lxz1EInuracCM53GIk9t0hXOdfIPtjGxAv8oGU/
+l9pNv9BksJuZt9YWNCI2oITfKie3Xv8Gp+Js2gXjMAk3SUKS9v6q6oVhmCKaMy9
uUKIEMjQaa0gpcx8uIRcPY7a4OoUQMV3QpJRDSAQtwj/dgMxxVG/XheL6z0cpylr
OLOmLZ4FT1vyC3kHu18PD2zjqvEk0SnY/tdDLIb2/VPXvoKjAhApmDZY01N58FDf
ZeOm1ZUmg+uWZkpoOMMpYnJo5kSiMh0tk5Ov4VjB3GTuZ4qR14HdGD3K7VHwhC9T
PASgYsD9u/WRVo0QFHq67b9cGiA3AShBV/0JvR+tPiJzq7IBm2qXFq9rHpKcusot
ME9ldLz1NRooeJ1+thy8eMutD4exHXA/z1kPMLjZQTYK1uEefKDYIL4jU4DmANJc
E+tJigbuIPzsS1pZlG4i2PygMtmwAR4u44XjZkZlpBX4xXHMJa7UeXw1Yt5AekRF
AtDmAu/3QfnBo4LlBA8FYOQXpVCRd2/6snirfOZT4Gi1xGPjqnbQpJxxjBwBF+vS
Vog8I21gsKf2UdWrDqIzqLbGg9ieRMIqCXdWqr8XNIu2tZgocrPxR7UjtCmqYWD9
ORWPh/rcBMzRIaUDU/hveznvKtRNOmV1hF4goL5kInn0rSdXX82arPpBIOscq4V4
3A0jc2WX41snbXWuQQ+Llpan3mInVWBZY5+CeOZfekGnEcokA5c5ZW+TdazPOo+k
t9gds/WfbUke7U4279/lXrSueb5IcYFKlOdVf7hiUnfspxCyYMLRM9GC/qTPOEUQ
3rN7fxTiWzxAjecdbFZVqqUNAgsYkzfG+y1H6daDRTdr/gM7WndcLvH8vV9E4si6
GPmnr4KPBQaGAGy1qLK3rhSLvJJmYkLI+7F6EA3pXvqFjf0LYO/dIe8iwa/VbLCK
vWqzwFStqHkD+wP0ToFOC8XOTdC907XhXaYWg1lZCxvnc61cw3AGMrFKrNjpXC3b
AwkTYSu2mBg7/pOH6NRIjeW9qtFMIWcPzIOdU0KUX6r2X/elwkLmTWU4zJ9MrALj
7P4FIEN85hBZ0QEGWEUvyt8EW4Acfc10TLj5hQOpV7/Mah5c9a6feBEa2zORuyYy
MKCsi3IR9bwslSZqYCD0NgwcEEYhBcxNLi7GmhFfCuaA54Mhv0ODcgRA4CtWDFN7
xbuXvWeCTd5cvXLml2Pg41FA5+SdcpyzD2ZNEzQYCf4kixccZLXPt5ofInEm5Ki1
1rM91GmuOmZN10cLjteN5Lg+huptUNGLRzZBuNF0hPePHH7NmYx8IG5Q6V9Q4/TQ
Or2cgRSemLJ2Lq0HxQwUDU42qdUs4dea7qmmE8yd7RbEsPKECJ9H8Nun+nMaRGMg
r25eMdJ8e06ZyOfPGUi+fR8bX8rCxjMxE/tqbQ7Fcwy430Sb8gYbGyFG44Qn5Ljr
kD2B1Llbhr0LhaWL4yEcP0U+h7J5bt6n2RzS/LO1Aljb8VCWBuSt+M/BQqswMLoI
Guo49hWHZ9dMoVHXv0Ai1quiwhE+9+geFK8Ilgo2vuWkEvNbsE2REG5o/8bDiMwe
pqtY/JEBbZwOI1gShUJL+4yELQD3Ap/eUB48accc+DBboY8FIfcKwHNYqJK9tH5q
RWxpJSOJH329QV6+5wOJSWFON119lAA/weC3z8rZKkUOp7/XZSrN2+pYxtmqZStv
/7ilxt+DtJ+K+DXH1suvh8NmppTPAeAfIIwd2W/1aRm56OBSkNIctRRRhRhgdMj2
Q8KPjGuNf14bSeRhDH0R2TBWK5233obWGoosd5FDS8/RrW8WNYbIYQB0WTIuP0Fa
X9cYJKcGtbZKW83GVhYqesZMWCuUfYmQ6yX0ERVvkBOOxRFfGy3DQSgAb94C5FhE
fdKt+xCwaNfdk5Yyg6D3Gt5krwB3ZL5S2ldrPvzCmnHvjsaIfeaJRWLO3mVyEfDy
nVhFItOUPVm27o9BAdILVz8riEdxWJTuWT2Mliy4b97TYYC4utVed5xCPvZID2ab
R1nmcwAmLxAHAjv8ceeUaEEsJIfS+VVbm8ElDtHu3f8TY9jp43SufiHz/9XOdgZT
d+3SaTN5qMOZunhJydG0jpiLwf9TkQ9vrfx1IjeZdz3D4xAT6PfRSZGgsvLOO2VL
Y80i5Pg1En2mdbCdSc2TfGc2Sr6oSr8eMVB9my2pYJ7i6y1rv6QtzNsNHy5+ZBhf
m40Z6ebhNb3zubrVwgtD644WHRI6SyM9El07D+dQy0k2upQasEm1nUZqh2mVAPn2
UUk14j7JkUAWGxng5wXzJSsshZ78RHE1w+3bxGEPwoFp7X7VEREYDN+07Rpth7Kc
Yk3BVgqTubIUV+cp0ymwUXXLKujh4wibJtJ/7UU92dIy2MfF2MWydBmMqUX711Mo
QfR4ucVNgkXrKB3T5bPa9fnY8rH93Pf7LbkCSEg9F/Po2iRpBSWC68PrryXvvFGJ
MsZsh/duDuSmPlTfat1MG1lpDj5Pe5Xk/e9FgJH05Zdznbod1SNO+hYrIIKASOEi
u7RSq1c1BcC3RH5pNENsNGPZ4qR1igN4LrWwzmjtmqbV1RHNRsWNJs0eONAWMHoe
zXmXFp+PUvLtdCtGJBMnPrDN6usfXCZwRT0EouU4rkmu2/tdP8v24kjSqQlv/M1U
VmM0LFaN51hKvLiOct1uQ1IE7EVSRPF66T/UmJTRVoqFjKS08vGa+RXZU8R+Jdrs
WREPDyqTqEn+D3L7jjDqVBd85B8shRnjgoyQJ/RBydwSzII1Xvoycv210KO2RG3z
Gu6i5zBXC67E1D2fn45IiTnJ85sDYqbs6Jb+c0r8CLgdJmn+Nivtoyw6qHDbCfCT
fnReL6UjARrtG3WtHIyrDrZW5b3Ry7NnuVUCPqXE9TkeOL7xZzpcKg7SjQjr3EIY
xbiB+gJbFMOe9bZl92qHPtCOnumI03cSWHvMRvWgBOsyenYCBBI90/juWfF+pC4z
uTGwKN40uu8t0MKpFg59VYPd8D5EK8uVFHD45R7l+NeIqcLarABke38n//ENAa+R
sW4QEKCzve05hPZttozy8lTlnljKgnZCn8aY/S8sGn1QPhqlF+h51sQFVBPk3xnZ
+PsSUFUkq9WhXyGVCdtVMkl/hl/j5YBl603tzEuuyf1v33LCCoMvZN5rani9Sy75
7OzdqlcDJ3t33tBTIKiPKLH+03HfMn8m6MDDDiThs63Li4cEcvcqDUfNN/RAEUrg
dtzr5KQSBIkIfUsu2hQn2YG9jYCxwlPuprg/tFloQcO+Xx6PUYq4s52tw71Bp5Ht
rmvdReJUjD9vkThbnpzPHllFkfUbJgWzF5SHi36cKGzPvgRbrIDZCjCM+2r/QkvH
L0a+D8xV/eRceXXPa6dYZvIKzM1jZmxsWPy4wbo3AHQJlUKHMN/NHmpOv/WIYeTe
DblpbcyhpmmG8KPXBuxYkAT3a0qjg/3FpnSeUDqEBOpr2KTq9elijVQ+QNFdKy+d
1LUuCrE6jHSSCLa5kp25SH74FedNTy/IysHSNXuQsrJyc9bs5e5qXAZ49u85vfaO
q1C0ibjwdDGVDpUADe/2jVG2mk8uRMOVLYAnW67kpP49u6M5nkaM0HnU0xuKehWL
GjSta8Cax7LSLunj1oqppaYefbRkNbXr/BlgxCCCiQ4stl4U89JtSDbJeMRQAjHc
VikIO5ozKh7r+bQPE0BQlLclS8vepWutiq43tLZ35HIhVIto/R6NQ/3FXZGVBXRK
pE1OnxXZmXupNXAUyrKOZjz9c9Ud4bCMPfBlfFS5QYreP7lXa5V8L02ax80hZ5t3
oCM7KMBybc/h0RibrFKAOPh5TQbuOgq183YnhuuNo1jHyAUzOy+pd/L/9+rKYT7T
4cQRPoi/Yt1zfI7/wpXCojK68dJRaKzNz6cD+QpdV2z/P8hqmz2Oba+xO8jmc3HF
RVkutXdjMOAa+D+6GG4XJr3nEOlP8c/KM0DgEXag2ACy5hWfHyEfp4udaD6VwTyc
xdsZNuT6jjvgNlZhUldooTBh8ImN0WBUx8BGvBrhFL3mBgBlGH8kfcXr6brZZypL
+/NwIirkpLZ8H927tlptHpQXg388EkBBLraWZ6kvgmgXbyUo5Px/1a0qd3Wg7bym
kDz/7JmiQuGx1u1T6UyfhdJfSVfGNGdsO1aM4gWaDY1y/Ce+pdBzm/DMS7Fx2Vnc
a0SIpKt5u7fyJLh/dqy8+7zlZ4KmTgGRJhuqol27HMYVZgP4yvm7T4b9AZvV0gPP
WlhaYrJOR7PB89l/pAsDhBt1CoSwXDIr5vsYrq1jqQJY90Vg4cZaCWx3gfAQW0Cm
sm/C09XMUYjWcKH1YM1XXm9LdRjBDdLK4rTPNDayV4nLEqn2LuR63QX1Hxe3/ATF
iYa29mlwPSC7OvW8/ayO8J1PO5ekbzD3LnniJixlSCp9wi4TDcsNtQfIZDjqOqMN
ZAWUo/OuPXeJgZTZB4Ixzx/tSr5qdVitiin2d1Ib73I94U3vlbqDIBeRT5or9sek
17j1YPYhvidGQAKc6fvysokSAJ5NkG26WQCJ2Z0l+YDXd/vhRd9ykQYGXyK/k9N4
16K869QJ0ILjdNzK5JhZKlLA+LMHzIBeiHiLER8BaZ55xOcozo/WH0wAq35J/lr6
JTkSqEu/17oN9xsXgYzuyFEnnLxRbDXj8dexW4utYrnKRHwq3bB7pyAniJhkz90x
snYz4z4Y6hfZAgL73UnUQ7mRP/qTEhsnHsLz/ZsdpYPyied4PPiqvL+05kR+xFOz
c/+X2nwtZe1tueTR6SHxGuCZk+C+wYkRG0HQQ7JesHQd+KF26YjHjw53T8JjnDab
yFt/6z/d9DllLbmLgH6FkKFzF8EHptWn5ijapvww1Y5bUFQs+x7ixc/4hxhdfZdF
jELEMu4O9/bElLS8JhYFT8tlgoSDU+ita1fN66u+XCGuwL8A0C9mOOcswUT/B7QP
PF1MHZY622jqDKkWAWXJRCEet51td4VYcx+G3Q6PlfVIIztx+PuD2rEq8L0tcBgm
/kVrDWdAKB3Hi9An4B82Xo0jK3he3zWAmpKV3dtljtYMjpLRWC9xGKT9Rwj13uWH
m4PuWdJJUvuOy/Uu5ZN2PqTohThMzRmhGBPM8fXlSFD+NpNutlTwoAhJlsiilhaM
2LblgWTEdmQNBF+capt7hI1RH4PIt0Opt0+trF7TCGsvh5Rhj5SWEln0pzLC3A3E
ZYHd84rzlgeMdAu3RO1HMNWe/05XRSNgnxAxxWFGCg7hqBzdNCyiBqfpQqIlyrjF
zVVDiNJNwfNPTTbZ2R4mpgsVryl2UwAVW1XoYu6XW8qLUlEcuW465/hXWnBdS5bw
i5+eXxM8ALkKzhQm86NpCQd/vHPXytjedgOrZvcYQTG+snJi9iwn8+NV74z1YZiQ
poIeEqK5YBgbNH0nrpsBuf0odJGdnGPB0lsjOALujPf9wBZRWuLAlC8IiZOnpU2V
ANj+RRWF3JPRlhYNDWu20RYbA4cRmybrqFi0HyIEAaPdFIBNSxlJZSJ4H+TqdJkR
lCO7vD6Q7vPla91vWoyV4vyKfMFVfltHb/4M0NaOeaxzKlUXyGsf5Qh0Trl73zic
c/X6c2iC//EL34RQx8EGOFBcOBDUZJrkvxwf7gFK1zajWPzOOpolKucKINfa+nYo
RzQr1swu1CT5ZXMzfODQDdwhNDS0mYDeab/gRsbfjjJRiW0fc8f605FDpl5ExxpO
pk9zjPfb/OMr/eUi3E+fAqd93RjxwIBJgSU17cGk94rMLAKer7PctE90iMBRy1xv
hKchIFbgK1CKaBkiGvP2rqVgCpobkWs7pR90Am0hS/v1mBW8Rq2ltPFKvHHl7q+8
6GTvr9u3VoJXN8BEFzHSGbDUG5VftBbJ4TpF3CxY/hc2MiUtzWqf2DJ4aU1vrMtl
Abqq4BaHSWqopGXe0PhjSdsa9Xj2b5wypYAFmuIUpKFR/bKi0xSUYYrdUwLzIqBK
oCcjFsLeYehfdQKthP9uNNCIj/FzTL7FhZRHgFH+zpxVWrESDzrXvz6aUVZ8heXV
cbeKcE+i/57+rSitpQMV8qHNdP16fjvbZSyx7J26uuLFVMC/vrqEbHZ5qGQOHhro
72IkDHThvxQ5NXkWJ21ht2+2wnw1fVZkStJ0LLodF5lpClphLa7lUN7SWLP2R22i
OupxAwiOO2C2g3fOYfdnR39fiZvOUFrQb6Rv1ZpeUgn17eUXyWbXwNKkNcHUCZXE
aBwtPWh/y3jcwqdt3uIQ7veoS+z2NfEofA03qUWmUfp8W4p86s4d9YyHaID7C6Ns
VgmR5d4Cz+eGQZNceRInrNfz8Px5WYVRPwjY7vK8Fxmjnc1ylIp/QKfxuUI4dECB
C+P5Nr3sy+/BV79WhOdgEaFge5zUPkgMnKVBgyDIXedjNPElyyDWNsR3havL/fOp
9809ztQ03Y6+35pSAyD1etWhqnsoTcNLbwaAZ2bvGeRzoIPobJX8hcK06GxoacPx
3H1WqiS1KP8IHtrvvvN+XZUyi4ApHpgmiTEt3KvdyNhqIDhvTqOIHJR1aoRC6Uka
yeFEtUT/cv6X52LMZQZSbuAiolfxLrz2/NVpA8WYUVlJPf+T2KCsR/qYpdpVO2ii
IGc9Zv2sD/O0q2LpzbUTSZ3DxEDo18CRMbgaLrYqzvPv9pQJhi+LqIX+sZcZv1zz
s1tviJtuuIRFvrSrMzaAMoA+UoBXqXdf68MSWf2E3HOWA6qqXNoVAWQwb2okQoQt
GYhhTrY7ziuUQGb6ofE0CRT0n3DW/p3+PUWgx8wB8GQZe2ar/lwMTvVSLO5hqcma
2wMljkaDsNB8sUDNhM/6bi4aXpmbY4yWqpOInck3LkkYlJGNpwKFCranAPtacGbh
x0MmvZUrv6E0J41+Hr6gPy9pWZTl3hZjaN1AARvA5E+VAFRx11LoYuSTlkUhOmHV
Bw0F8UC+AnRmmrW9b2jPbJSJM0LO45JiivFbvCHqEbjxNvWUz2hLgqDG34Sk8xQm
U1wJkNwawMDqcZXWytAs2epjzFa88jCSna+kKSJZn3IPeFRyRujOvsF+1Offu+e3
Qgdq7anVWt9aLCw7nhEMcfbMm7RKdhkY9llvhsxUYveUFMMXLPvwIEB2hEHdHuDv
7xDCpvatgIO68PptVwcevcdknUkpNteML4CqSM2iSqKMrBboMvsWaMBpyYxYrgL/
3tsd+YNufnRLb1KxiiuqzG19tLvJy1tJb7Ad97WMcZ+3n5U6u8wjBOVu+PbYGhse
FL/Q0mVHyHGULWunhnF5mQ7Vr+K1dAGne4ofYjWF3HvD1o9hTfz6Ektj8Ug2AKd8
ddM3RgHL6MpOzFdwyl5a82kTMAMLXz4As3WExf3CI8Epnh7OlJNLFGAKvfzN1Nkb
XDW2ZECOfCbSozi8P+FGYK2aWhkKcaZuYZTh8OEqk6QC7E7jGfTZ4HIG67Xlevhl
+YgpaBoTktLzT5e4QewxyLAi14C5tyrviTdYVehqiOA9gLcyHRHfIF6G4LJUkAHs
wjhkqbjZ2o3MgNo4J1EGs4+JhENx4yq4I5xLhezwX0ZWo9DYzASvzkcgvihbDafP
qNwXrkCYtVZ5CwU2+Pm3r8Br999uphtgaTV0V/reYJ3PRIM9uFdwSkIdjHtrRn+/
BZW7iutWj87gPR14KXVlKsvL5jL1cqaOSisUvt92t9wxTvUzXZKbJcbEYnNtSheA
rd4+deatL7HFbBOFJqB9KSUVqRin4UvGcpBABTivpQguXofNOs5STRYFBDlIFu11
V9ryDSo8F9z2Km3Yf/otlb51tZT7/+kj/mh+BsRurfSW7/RxcO9nCodGUG2qisuy
teRR5Rhzkc7XwFBoEwmbuNpb137cUBtUl6pfynAw515w1Ijkv0evVpbza2uFuqqK
VEjdY8yOHJpdfbu4wjZHpcxqEHx2dyghAeSktqVWjcyb9+HxBihsaLZ0QlCS9bKB
WgJud+SBCamLsDjFkIpBLpEJcGKm/UgraLacgNiVD7OlWPo/dVMhoH6e1sWjV6/c
j2UyHgJrhxna9QiwgGkQADHfEwotxAj2wzftIqopKd80zYchqMDffarCaMkcwXfZ
R/GFDySwZuGyf2b5rr+e4luBo0/zF8ZHniaB9xGnH3z7ilt1VzIpblc7KqKx0OdM
c3F1XQJK41paIvdufxP/p/6ZgWODzlTU7sfzuUjFp0pdqfmQttf73jXmXm+bbwYz
P1DtIFTvyeom/31hT9cm0Mp0gz8v4ka4/6nB53Dr8XRyrvH07GOhZ3FxQ3mLFGxt
rUjJcqRTAXzoeUSCQ5s5DYS/+ixGg9nPHzRnAnfHSbomxLZts6RUipTSlPYiPUqg
qI/Qr892uKHb0AP2Zx9F33ZxMFEc7Q9HJRk6UfuzDt8x8HaOjbAqasqeDTvUql1z
SAW82R68l/2nV5O7dIznu0obeJNHgMrOBdOLGsQg+7fFi9pF6Vmn4xCC/tfCwBC6
s/HcaFbEx0Q6wVp3QOyzSi2RhCd6MJICclJamyG/XS3IvhB50fMvgDPm639If4rm
1wBbuLwrqjFIyICHaymfmCio8S6q6eCFSRq+C0TfL/MOKvgq4LGbYyOympAfpkDX
30EC3w+J3zhb4YdgGIhdF7TFgx/0EkpGJ5uxgpQRG4t785n/CJ+YInUeiy85ffp4
RolPtGxd+ta5q3g0tTQKXeK1Hthcof9zbs1ISgt2Rlm9o5wImH1A4Au1lWcd5p2d
UZOfJ/o2JbiDuTEUpRXHBwgikkv0M4dhw/EdDJC+45K61i5Rrazco7jjS3JktgpI
PcEUVK/bKHCKsG03kVtMsmhsL9ll3ZSrgUz9WDpCRY84DtMZZEtaA7zCDg2Xa2AF
4PoD7b2KWxM7X5bwXxSKPFHsxNCq0sm6ClZNBXtSea6ZVbmmStXvCfl2KXDuVisg
Qa2BdF0/xAyDHdy5JyNF0uSgLN7dMOaitoP+dixxKm6/9PC3ePklfP6XSlR7V9Nn
I/Wcn6k/EEl7hnNfq84VJvM0MuQy9Rf4/wvXyaUWwDkrnZPPW+blGupJHjZvCICB
acxVn0NXFZ6K2ACV/XeuH0bszaEnmNiB4ijePtxx9ZlxvRMpPNAJRnQjZvcrZqat
OypvtyQUVDQEvPZrPiRNRN42WK4LTN+SSnEblIwATXjhXKmQfNQ5hDAXFY+fOtsk
M7iOULvM3p8IKVwKcxvczxs1N/EOESj7Bd/5umU5XDIiU5HSOh0EDJk7L1xw7mzF
qHtkZL4PSGj3bsI858WgiqXWaRvXxAAfEarpzBdt3rRRARn4JHyoUx8iIcRmXqWb
LpHb+6kQ9uIq258x0vBk4VaXZlL3nwbxFUxKjZoDImTVrYlT33Q2iyoNe6ALn2wJ
UAbm8m1NuekPbzyrdLVw69VuxrAuofllBL+3+f68txp5ViBmXd0Km4rec2uaJNlk
M0vEMaav5m+2/7oV2egKcqCOkZXU83jAMlRtmTuLC4ECL+IRxX+4iF+GQ59BA/aO
7SJQ/lv0hJ95IldAfLsioJOiKefaD/Wt0nBoqZyk9RByZ2wQyrRe52RWCLj9V1y6
i0yzwIyGMP9YkQS3MeyRBrsKsvaHxiwNBJts4+ridpISB47TG4gxna/ULt3188vg
Id3DdtbV8draBX7TQ1vWoCDY1+l66++PsKDaFQYwOM877bi31oL+2Vk4XjTT/hP+
PuAdvZ2zkl9iwyrryXfD8ZAXV27esN+d2THiKLEZDx+xbNmJrCgyyKKjkvcyecmt
ICWbE65R/dBNAlyvKjRVCAwGOjpa3ZSupFZRw58+2OiCX7QGw+r6gifWR5wrslrg
bTZ1D2GCP3LRdHLyKHP4aiW0/e4pNLJTo39eF9l55+qUI3KdehvsDOBSuIYSiMJp
TDcJdNHZjnESCXQuyBhNrOpI8RJxexSod9/XpTB54X/h7gKEjSSjJEiCyiQAgb2o
cLemrrzqI1BugfbNTzF4pwecVD9jplX3OjNd+IaxaQ+GxFSaBCpqAX0007p0nhxr
Vz39M52ItMXj+zUY4GZ/2zmClrRL9xD/Xwg++2Kbu4SbeQCA6AVcKQaurFk4DEWX
z7epEut1JbJzFF/a4HXwUHAphKsGvQIdZTYgY3lJdn5XyfbmoFtfm8CTkNQlmZf4
TO84KiSH+nQTVUBa4LuNtVzOyFwJw7rp4YkAIhHEhSXCa+hVvmUA1nU2JtEyBmfu
ArslD+BYhtiotJw8pOQlDRJn3kVBuKB8OZjq4SC9R13/VpX8o2w28E7NHGky0uqz
p20XswnUlWbV2YZ4FgyuxgL+SbFFahDDA1tV1w0tlwHfWbmwMCivy3YE/TBv/Bss
DG8JMaCF1hWuX/gnP6bSt2tbYXxmC0TqjbO7qbLuUEGuKLUiANfFBEcHuUoXqE1v
z4O8gLgLoWkzUFykQ9HrT8xqj7zfDGRVBsCvBRFqFudLqiQ/+lKFNsNt+Bbh3HKu
LlF3bO1G6iLHxEvSEOvHwGcTSCA+KcU3UMHGrdDCLO5WRU+wQz0QMDOx6FOyaV7L
R+5ezriHLtWtXJJ8gwa1cq7qHQkJMEcE2lzERovWBow8YH+7NISZ+9+lV/LFFHc9
gBI4f1iRGHYFdd9nJjDzAn1SUTg0qg0yWhNpHTelLeCCaF1mUiwBdhmETdDe9W/g
LockIyndToMHhMCbjoWX3g3ySX1Mg079rnRMlxLh5GXZ6DcpaVTJfSPje0evEmID
Frlt4IeQPDtt8tw95vd1KycZP5ETXNl8t+XJXfhmA86eUBqBzeLdGOZnMw4JNLZO
vQIPIaa3szvWUljVZp2+7Sn7/AT/Taxva+4KwlUvVjqKhGyh8Xonf8EoJQefJxNC
CfXWy+NZ8zBZz0a6XtVh7RtYf7Sn20SpUIevvw3J4q7aV7+oQiISAggwqCegEpcZ
GX3b+dWZO0QBkP4YssxGmoxS71ll7V8dK1mAaiQUkX/x5WdoyY0c3l5QP2dOmO89
mpgR2I1hhV2b5NiLb7W4APVCHZW6M7Q1aGNW/MhtC86OqyxqnN5ivCgQCt2Y0YHq
oK9mQLVk5cRE5f8ibNo4lri8JtTYisSyJ5WHYmiOJXd/KbWu6fhUoEgFGRMyBI5v
JEnaeaKpCFeRrpRbloN9DLUh4Wn6xiZpG0678vo7TImG/0Umq0elSHxcCogimq+V
VwrGDwYD8CzlX2pSJ+ChRErwPeYfaW7LpbDq+SdJAmvcPWKfbijLu+muU99DsUPD
gkp3knHinOxitNgPHXkOAZ7R95tI+Spc6KkU0u7RY6rxLfu+njT4ebYl+yzGsvmb
rBqlzgQSbnXq49cyXLZF+fcLkQoGo8WBX4X48sP9r6ZyDIFAlQ+vmmrMkCZX9HxQ
fKHmN2R39pLWnAEgMJaT5dcwH+bxe9BbjunUacLDTPQLVQszhjqQcTHRwMv1flaY
y+ZqArFzhcRTYlSBAZj+U5XIS3OaxA9ZjuuTVdBK61QWXud4NSDgQgShK9r4tg0v
i1cI1pJmtUMzKUuNf+llM1GSML7/wuJFVsULx6MSpD2vo9/roq9MYIfRuQjJTJDH
F+0Bh+cg1he8GYqTFN4XmTyKlpcNgps5t7d/+Nbs4jWqGFLQFBF7rFA4Q/g0R+t8
FrxPZkRHYHAZQzMaLcl0s+yocWmewWJrHwfsZZ+XY+e0aaQyrRgR9rCW6SCilrIp
ORpwFizFfB4UxoW75AKZs7+YuvgUpBXx2iP59GKCl87F2CCzK1MEHia7gjiXoisP
Meacb9cKXvPnupdDgCBSQtkZKE8M0/8iqfZ1HQDV3Q9fE2TJnysmmJS9UBxhU7FU
c7PwVWoCl1fkiqtp3WPu+ooIQytJpfk4nLDydMblzYKyJle6rvO2EMfisE4SRWrt
TGHuvWKaUNrTzDJeSUITRxNwBGyMb8JFfLzv2Qf5EvZcbaOsFFHh2JAbcsueB89g
ucVl+aigCZmpIAoV8YYBkpG0+WGsoqaL79sZU0faewSuXhLYTQwl5CTR9jAjVk90
z8ehoSscRFs/Py0DuTdFSBQaqtB7wFSFfgVZPkYQMRX5fnFAB1biGGMzyZa0+/XL
UA81q0HCmFb6Jw1+zRyJOMMmhqyQh/8CndCSrkSZ4Wc6oVPtqtLIrX8S6RuEraL2
Ysp8r9Cb3CkA3YqKmbTQvlT+I+Q/zOdl2PoS4n7a5RM+fTIjbMUvoIsxun1vpzST
9TzTLSSgHqoFZrxzoPJrfXD7GP8vYkAmB/VspH/yKmtFJMbzfdgxVpCDaXk+D8lL
JgXaPXXIAwpOBXRCEgaJKDrLL4rJ+IjotmS6SVbISIShGym/sZ96M+4hFimdFUk/
eIKz5qdttmzzZ6FcOXTKfySAjKjzm9l/izsCn3UE2fnV7Ts33ooagWlQnSkVdd3F
aXNAqT/I86O1/tqR2XMx9L5sE5qfhaUTZtSQMhL2TcPiBX+zYU29h2do+eTovBl4
L8JIFNXkDIx+jSRVQd+fza/PCRW9L5Pivv/rdGbq1gUyn9hC/rJhoB7GB13eRYZa
cjvXI3bJKmB0kdod8KI0844dia40bUA4YOIhs81TA2asI4wqVyt/PKdVk/6hsbCK
gdeFvEWF3EmbrSe2ohE9ke2nu2WjGP4NrM8Yrs68Qsp5aMuMtkXT8Qdwm/1HGfb8
po/XLXzKtUC4tf9qbqMutbPZPpIAN3QpQxrML7foVk7rOYz6xRp8r3vCtoqCTU55
lrtPn7jytu0ms00hQP6UDBlfKzwg81D4wjPrUGW1ziRlmY0/rMrkaLK+o2gxmi3j
e6jc8GQMGRR82k5VbxqX47bcpEMjRMUNiCnkeRgfMzmhOV5szfUaSeHVEfUJEhJu
8WeuDkKmIIyN8Zg6Lv5K+9iQwuPPfYU3WFDRRdOseHKZjPM7h9uNHeT7PFwbUFyI
4qYgHp6D2s1HuxTLGbAk98LOUnPUUzRUxQxHDGb/mM7Qz1uHdcFV6/V4strKLBD2
I6a+NW7pUflMk4LqSdZUmXCEAz8Y2qmVpc2F4rjRgt175ig8n2++Uvwfr/de0XWX
L2u8hd8F4p4fnAGXONJayis/UMpiBzfuNrciHN0GwkmSudLV+yq29pmfk/fsDSKu
O0rv3+6WZJNMjl8BYetxAlM2T987wBX6Th7o2b2WHXuIKXzKpiCyvaO8034+KZZ8
2PLp2sWluGWgi7WIrZ/+QIt6E9leTKtFgByzcMt1Po5jVMfYFP8uaX8v7MlnsqtO
SNCxzs+QBB1jPi116XtV/ExMAjTpppZOKd8YLl1nUWtlQpDBitK+n1Atjt0cPGYI
fDGOobLCXMBhhqJIWf8FTpnrDuDjUN9tGXpcnB8a4iQ+Cnt0/KrKUtv+9iTBXQnL
GBnx++/TSf2fK6nL2gZ+Iye2qSf2LmWgvopyUmuPxmgi9oTc7KcqPWPbwuiUzKoy
JfhesgAmsV8QML8uE1BIQ0tWQ7v2gpyCPzFhQ0gPe3+6raYKWjZ5J7If5ZdB+i2j
gmCQTX8KcD2IctDnmAsXnW1YioBfcSniOTFh9Yl08iPZ3TsrojMOAqoVMOkXKzyB
q2kPBnUNo/KSu4Fog3QBGdRuD68hk8JDp2EfFInH4NMbEQyvFDW7HzA29cfriXYX
i4f0zXrVgxtkgfduRa/q+BBemJ85J+XqKsElMAM5/Xyr3apnZKdvIGDSUUAIwY7L
4DW/tZCTD6cwsDSKDzZeA8qXTQD/zDl/jSf8YPb0sx+tGeEByiVTke2zxUCbOL+T
/5cRWtXo+ejcv5v4MjDynFyzEtf3WBgsG0wGmxmZjBwkSVHhRbAvNmtzlxk83jlE
1Nyf0QclbSyhVrkBY498Fid1HCVGoqoxVbnsqAktAvr61IR8Y9NUofqseG7Jqe31
unmLUp1iX2nS/E9W4DXc9CYx5aVERAQ9WUrf/MzZeZdodHJ9txjpa7/8KPH0cb6g
aIe14JomJL5loSzR2tGKrs6KmhcNlxVB4FWXSUG9RmW1fd82PVACVaQb4EoBmmpR
zQWu78jcaXb0e/c3v1jRX4T0Xb0ZImVGnXKUeo3PVdpgEuXNAn1xTbRAjaVShILq
u+7wfzi1Fbqdvt/1Nn070hVMH3wwfeS0x8dc3BtcMDHKuZdBF4BaoijDnP4E5T5T
NdMPGIpM+nx0y/tJNCuqHOYxb+cDfEU8dOe2F5sM0XOkqXM8WICOrQvq8AmSuhrc
ZeOgXhA+Qv3DPXnKQmlw1va5KHCazA5O9PgOap+vaYUBDuPLX4zEh848dwB5pBXx
DZGh/Zuv1lZL/J98b2NDQibN/gZ4TlyIFpjtjEBg5hDjybewiasMdlBF2dDvDjdf
zZ+4/jVa2fXGkhNRidX3D57Wdh+tbqacAnllousO4pJyBMB/mcxx/jiqeiIeDLjs
zM+SG1SMhbvKwxOJwt0pVmFAC0Gm0H+LgdoksCXDQMUS3Bfag9PoUMk0xsfC2oJu
lDwDXfgwDIAU59+X091OcFe5uEz+6cURtR7HvkSOh/kHOyFjnyqw8wdbUJKrzz7H
0mI8gmaHR75w08Lbo9lBHvTrkqQaPXX8cMdA2r4yduOB7wkgVM0Plq7zJbG+RQxD
nUFm/Z4FtZW8VUwyvE9d1Z7eqQQQDfD+7L7KOamaHyKYfaxHrBZ49KHqziPpLcdH
p5/o/xsTEDYaJ1I0+jjvjF2JwVcThFiTvKll00jkA2ZiMRtreeEQA3S9KITvcNKK
O4SAQwi7RPQoxT/D/2SmMO5Gmwo5HXvjt3xLS90qKl8wmN18ofXc58M094eWoKPr
NeoFfsQrdhCWHWjKgwfq2RFmr1qj/PX6Xb09h2UYCKivPyyQEDqCZsM7Uo+ju7ey
8HNC/Itvu4/brjgkM32n4qqrkE/f0u0UXwPn9Ie/4yn1xmOJukSUPTxa9UIrvViw
QS5GXSJqNnsv7o/B6979/5txvxCd5kq4uSSfu4J12cvySfcfdvDQSyWW8XN4laTl
Y6hU36DzTCLYIPwSO1vwa8lc5yMnrNmktVM8Gmfr3F6ybsVDm8S7W2/yI9PUlAzc
6irfiyYRQhsz5LluRDriLKVBS+BKPtAIAVKHR1AJvDJ/x5fpIAaS/5nUUq0Ycd7W
6yECXmT5+TPqcoOlxyfvExIMpjpHGcY+OlonLKIBwcGfcQlIKdJDT1XSqFiXng8m
TQ5zLABJcz/f2hVmcg+F6NOd6IQtUOhUKtjOVrTUdUiW7suxtc5+bCpCagmRZjUj
A5Bf1XMiC9s1thgZ803j60/QU1vVRzVofPt8Vdma+oNXQfKbfOX5xUOKepdjBQAh
FIABNUBhhiixaU7sn9B0mCTEzhTIMzHwTK+k6htwOZpOKAJK3DhB7E9ElAwkWrb+
50yDSYjMrHgnpEk1rLd6YT+efDG/9e+GqTr7de+RVbX0nFatyBbwdrCmSdDLJdQx
LXvKn6Ay9YPQu/JXBA9hUS7JPSuMFHx12uMILSgd0uwi81S56JfracbU+ggTt9lc
tS2u6fqfTv5Lv7KNZdtZMFmXJVhuDYNmrkT1mYX1yo1HGVo/+JMlXWIWX9kKUmxw
2mb2/yX8AfrpIf8GTBxkd235YJnVs7884UopOxRolgGEqMj1uRhN5P+aHj5VHU/G
oyCVX6MzbUWkYz76l3D3cpMTpKWIVzhByYqHG1A2MUZd8Tm5EbcfiqlKV7yannuc
4TsR6RWPhic3n/VT6bfcWmV0UPHzo3blxZpLSYqoYxESy6dkc+ATB86HgsgRIWP3
atuShV0mA1kLxIPHYGrj0i8dNmDuBbc77Zr9EMkgcVAH76sB6G40Gyl+mvJAtEDx
XBfiS9C5hdHHsl3Fs5w2Ld5zIusemKTENrAqzdqaShmvQsG4Igz+cr+ygisK8ief
AOcMgH4/z2oHt0rk8TYKdMMgZHAkhOzcDCOXLT9fvvdV/Kh6XBK2UCy+wqk1dCSn
q7SEOJI5eo3ubuVMnTt7esOD8kQeJTFoDwoIIa5uMsF5wxSmNJ8asfiLWMLeqIkB
A52VAzBcAZh0sX6O/8MyvVc4GHm0qPFGQCcHY1IfzUZ1rE3zADfPJrh8ihDr2Cxd
moPiWVDo55xH63TuBFkS2dci5QSMbzSSnAiNJw5BVHdDAx30IBYb14H4JpkfgBBE
rUogiNTg52Iarlc2BTaiii3UI304IpRtQc83s2NyYc4WyP3guDd3VYIkUsmToc1u
gmR3/QbTTWxgl7HNH0L5z683rfwb4fnn2bWvHysx63Y/QIHAUClKi/RWOtVuQNyn
KbLxFiF5c+R4P4CXAVvbFid95Azi5/1mPc+tgoy5m+57vnNk6jDyLDkVWTOrw4+7
1H1y5EPAJiHKx+/juAvg+4mu5GQQhGS5gyIFJsPko1tnxq6hfmJhDM7IojGg7xug
V+/NQg0/Ic3UUWzf13zU89GumPtZjAbGyxvRUwTNNhiNVpGT9CiQL6dUJUlZdyj1
rDIrkGGDjintFmJQ3TGOxKGkSVNEYTGwvBu3LjimkHTneTyVEH3JkvKJ78k5UoGd
Xj6vjU8W05wELVA3uu0wr5rWwqTl7AKqlokIY+mGtXSuAlNjBcgegMSiVnxlbCbd
lnFfp1PyZ4PPBJi1z9rSgv8thn2ubVE9J5S5fBpzgV3hVigoN/L+OpGHduXJTAKm
Ko3RSwW8/YMcqLn8Phlwc3ZLLrDWJVz6gbBPwEimFxYkSmHf3WyGVv5QZ3oY4qXn
xMbhIyqNxDxoEeB4kkhdaAQuZOmL5B2yMnt/Q/u78oB9+CTkFGRML58ygdke3rZL
F/nIg+ALHcUe9Rb/iIbV/YqdxzFCkYzogUp3RxYVVuHZmt4KxEIPQ9TUrk5ekw9M
utr1lCAvIaatuq3tGz2tPOmVwbqsXKzAvVai0OyWCSEJ4ttWX+nZpl2I1plBUDsf
ZGgVZIxl2fL3sUztCDLDGU0BJKfkmhyQTTcarnnb9Eclz5iHr3a5MSQY8gFfkal3
MS0f/4fvgO8mKC3q0KtQMD5vSBGmWhSFk3/ValFmfMKCqmOv3dyTP4X2m8H9O+po
cwYUkpnmraK21Pvrf36kjtguvDLdQG5Of43WCQ8MXRNpVyIqSvK8/KCeXw9C/Yk4
KIrqMVYS2Lb3qEcqUZ7CAp0SvJ1g+iLWaOy6SmfFcb46ypFELx7R9L6/1wdrK861
LRwc7B2wg9aADD8Zdf8aVUczA1FxakJcV29QFa9IW0+4pwyM3hqjGJ95bBOIWJqp
j7yDXVUnmdYYeHymOfQyCXLw5X4z6FBcLHrWZ23+5GTePxuhXuSQ4TwU+eJ/B6qQ
uUaapnZO5m3KZhQerGLKqJTBX43gpzZk5YJjz2yVdyXn5VD7JcDba4TgOIgqTExA
HseJ02L5oP2UKiWEOHNq7riIZ8oANKm7dznXel9LJKKG42HIqo0cG6jpZwo6UT9f
QS7S1N2U34iTqnwgFTUZePc3FaVdRiRyQ6zRs23Nrz52ZITj5L8+3F9s3owHvHBc
M6/IfcZt0GfjTE8WTNLqlczqAk3McwI0RdFIMx2ceK5o0KgMtN7/LNE8VTRekthT
j5tvsFj4jODJpuDCeCpl1Vhi6DMDpad7e32j0qkRygcJDAPwAfIUp7ve2/E+SVQ4
TtHk65KuE97zjkT0VRnjl9gB4RyayyrRfmvrcSBjc2cNe0B0yVuhUIVV1COUMYrk
4+CTd4ygYZDQ5aVbjSON++T2BBa87jSgboTELMFrhkBNwjiRs4Ulfmgzbhs1UmL9
I3hEz7UJyvGtFqsMYhdPuvMobfAytBuneNXd0Ed8F7O0KUYdrCzv/82BBMepBljh
llHmGuZh4GTFKAtp/fyDKkiYtdnT2fRmp78RSTMecBNAhFUp1/xzKidb4+CzMwoU
wbw6obnqjzrPvrGlDAxZx0ozHnMTiX9uKwhV+o3nk7TaYQPICcijGswNxBf13cJ4
q1tkcbYzRlTH5jABNW7TuXezeRxxF4kKu4By3TAKyNJMYpS8PE9Ofg6fRePfLPN7
/2/VIFyuSs1iOyjnipMMMwTM85s2UlDzlAe9KUBTBI2nXG30cJoGB6WbjAurXqDv
g9xdCG4sSOkg7hOUPsGSrFSl6qaWooED/wRSqsERA6MJLFdiPvSV0RJqqJSGYiEc
ihxTO8RP7Vwhpih5g6ZeVQ8MuVLwx0htGZxmNlT6WkJTS9EttYTiIk6DooJ5UT/7
o0KqbHW65LWkyfagyUcFtg3t0+BUWjS//ls3kW+lkvC8Q+Y3R4CITzJSRLHcPs3f
MK5nwyfuDei9bRR6J8WGboG2uOVBZPcVSwQRiBSmZV8OoMRe6XkoaRzCx46kVqzj
2G/1Y76i5uvk5hYnSnfVhm9wL4AKySXdUftDBcCnJSxfQ4xj7OQjX84wRZeuLr8r
nRCy4FTXLkhAwRMc//vaaaVH5SmgVscHOkLnH1Gxm3UKnAXqM1bHbp1oALEB+5XR
scv4bWjP7OrF7dnRBM082Ig2UBzqEb0rGj00LoGL2PMilclaJ7J0CEbXz0y7flv9
yp9RpFfo/SeHLUEJLD3naFSzcCTXs31IqTZ46Fgts3JW+1uZxyFWPdX8RvWTSqEZ
XDfqJGdOiZxb7q5Mu0Ugcyo9k+2t+60feieBubjMvqXqvCaMPi24EL+Bvx1t+QZF
ozjomYsQNsR8zkeTsnN3v8yYV/VkTXk6HQEyUdvKVBfxuJdk8vmwvVLo9MhRzR0m
wrL1ezRY3HiNVp6Gv0GL5F2JkDnBW9AvXHG0Zo1kkXTUa7GtdjVhUY5umOB8GhdB
UZIKuGSs35L29oZZ14ZjZTM5l1vn1hjn4xcbUo1cSNb9OVrrDF6eVb0J77h78u2i
umnDtpiFasiwD8GBtj1uBXjrMaBw5q9Cd/6rAqZIxCweDKWC2LLWlGS1PZrSt2XP
N7dNAjMLe5PRu3362boPxu5PD/5/FRmUPqUXzmLrvnh4ME90lICtjlu1eEB3Q09C
CD4ZzHmoxMxDencSbz4m2GFdPsYCTUC0aIpQBqIAowoDl1kC8u+xlt7Wgqrtb/TZ
EoacIb0/Q843nSvjwbnRcHcweTM9p6y0zEOmzy4O3DwjOriE6GWhORJJgoLJjNtX
lDlgrnf/BbycADp170WgIJwRjixNnlWDNxOpoBaGDhG1jd5HsE4CJLVcCeUQBrve
KsD8ihAhCD24nO0G4ET+a+9uSk1eXr/jxXxBiczcSEbTw1/oTvNUyr13yI4rfUZR
bxbCtKXv2ELYNOcs6Z6t1O501uWjwiyJAKafjGLsU7+a/DgBcxDyh6QSyVGkI7iD
8/8tENYfKV9mKZ6rBbc24sdeWCb/xcYlXS9zSs0gHCwwgVcQiTkzabO6BApvkXEk
u5hz4i0PoG8to6tqCj8TuUZLaRP3LmFBl+R8VYCd6FCglucKfmQCfwr4p3dMQFLx
HKr6Jhq9ghVbVqg1mi25548s3iRmhuF4i9SLzFlSalf7YCnb+DsfVach2AvRko9Z
4GtD/lm6Y+ngfdz8REE081Kri9SO7/7NHVgMkyJzf+YteJ5v3yHUFuSeTi//uRNd
IfAMAaKM1IA1qK60ZxLtuQsOthyhXo+pH5rsXxVfJ5PhIx0kq2TLCW42ZPZEUR0+
xoLZ+UNJafObW4LLpJWQVBx5kmDnKhBz7cjwVdgDoR1Eu9QY7CRrGERufqKrLI3z
92wY8fG6BoTKRW5JTMx8n5/t/RgcJmQrLO5NIGzQlWso4WwoMij3eSvBZfOTwF15
fOXsXIzs3QCEnqfAXeCnq4F12UEWOFH0/uUBm9re+5L1fLWXeff2nLWVr0R4a1AB
bqzr4uEp33EJqlJdv/YS6aLjrhGqGLi37JHuMIMmete8PGHU8dekWHiy3iZ+QRSt
6benrlRrpJTSIeri+7+pdH56cx8ohMHs1tZXDc5Llejz0Ve4jRr595ubS8IWuNUW
6+OJbz0IS0bzDamQG4liImaJ4vSkeqqNWr/Vj9FYToM6OM2Wv06XCeUL8tEOpMfj
GjZfKA5CWrkr/CQFyvyefMslCqsCSvLafC2UjWMxkcaIUD7Xv/WtCA7+LTp4qjTF
hb8fHhGnyq/y5IbkIuOh5Wse3zZwPu1wq8kKgUs2GA4vU/HNkmjFEI5Y04rxERNr
rIKMMBZ2orRv+0B/nXEUiCPFoZkgk3nvJMn/NV1JRlr6me4oi7mQ9lxO5PiFwFYA
SlHNl/c62Xgsb307sNrvc+dLluFufGdc5C0m2xEJu3TCNG6Zc6Fflrcx1kjQ6AvG
YisjPDVp7APJBSkS7Ff0+rUdONjZF1AqQV08rU4JgKT6whub+VVA2tIlsMsUs8Ak
x9pcIAiUneClSedikRAvIraVQadLjtw3ruDq9QxpwTNlFIdhlIieq1SHpubakYZ+
ltRJgyP6iGlE2KqhYJ2XT9zvE/1WM9FotJQwBwby+wvzKzlZ7er94Aalei5He5P7
wNOVLxmITAB5xg58Ah1HfgZFnQ/ozPbRxOr99IG5o4Bjyx5pEqXNNyxxuex2N+s7
6Jg6nqe6Ve/wqe77P653E+3/gqBQZuRWU0+j8g7aK8EMXgx+DHTL6qe9HBR6N6YB
Y04G8jol4cELMBOpzCi/TpSXVpr79TcqP1T4/Y/3cDhFLahzhL9HNVczU65OLLYK
H9yD5AUY+uGm1ZRIKka5NjTiao5pCJgaVzh7fcp8/g9JqxGcLSTTdaW5QDhzX7K7
Mz6DLvX/qArdd0v36FCIwrfnzISaxV/Qbro2PMtrunFG4km3Mr3uObfRoOKvcU3+
Kfc1gQPdhiAnElfsuK0Vsg+FwOLCEMisHgTdtzQ0MbAfSa8IXERtddkHOP4U8zS3
6mc+wK33ZGK2e6frl+GUDWZXEkD6k7hVbhf93rFbWAdgNL9ix5o8rgL6JuhyI1BI
TE1riP+ALmTDDPdM6PCKmYnuBNdCzhg/HzeB0fZ5uvE5R4fhiZ2ZSlu0saJ4AVpq
xMoGxLWoV+QRh43SEgeGPGnK26U7fawrv2gL6DYCoeT2YUvGFQ9LJ1eYaXBbW81e
IanhaT3LEwkFqAc2RUOjE2eCi60Cd1KUQPQbJxNxZ/UHwLuXhKnsPI3GthviXYDK
lg+WtVq23khI1sM9fy+4FEhJaXydvLufj7wVhTxT5IdR0tkRMSQKQ3CIbwptINdS
a0TLIku37DP6jZgTB6MLS5CoLTJpCaD+VGaXvYm6UoJ2a60hx378GrukuZnZVf57
EFPLrnHjwFA2yW50J/SfvWI3neuvCSWjuZODTDSDSnJCpVaKF7djdwR4Tsa+1EK9
XZ3iN5iG5b+dZO2kT+e9rETQu9Y6Bkn7j1A/MAfgYiOKA4FtiICvpYWolYGGA8co
CmaBaFiKFwzztO7L1yMMcMVmcawyDi8vHMSyt9vv40Qp71TD1yLBR2P3IqQ9cSaE
QyRHNjIopRmplAoG+DlI1s42HIC2gUOpmjEy8I1arbYFDHi8+swrpRzEAkY8F0l1
XypZrW31ZJ7vH+zlXoRlpF9P5NM9eic6wjDkEIwQmtS+ENiIsNGFvFU0hoNoGsbh
jp1vTVXTtPjeHPtB+UvKIEOQHsXjvbo+Pn6TF0dtcnxLzuOzZZEBMWrMah+9sYSX
bLN66uUwfNYLTaktbd6cy/P7FEurd5uycdgwi7URapy14zloUiutT6BWuL1JrMI2
FbXySxK1QtTLdR3UHuoebyxd3NaKN6p+s+afqvLC19uwbrNT1WCmzz4Hc4b9oQ88
Bwe+U39uzJmghFGE6NfwvNPq5KdcKE8Wfc79cE8jtsXFviWu5R7li9j8jpRQtsQF
eVqxG/aHTqw5gC+9QdLojK5d65RGpO11j2FGdjWs1rjYDSNmorO5twcC4rj8gp2+
Ey9IhH4PCthR0Zk2urcpTE4qCCTAfmaCJEeN9YuQzYFC93rxfuIBrtRhSayMLSd9
QTFdz8IRBqkjy0jcNfi/F0VGtwIZfnzL5kbL4/s0GTBRYiPRFI5m4QthqndBGxe5
Gg91ezy18LszrcYLpH7hzFEl8JnNwvZpv78wx5pkeA4Kv83yVHwcMsr+YVQe599/
tw9fhC73ypNr2w/Mr5fu1dN9+gp1rDJkWZ1upH2VByNORG2VVNeWNnp9BOeOjilr
Qd4u6JhHC8yELf6qE8di9WaGkfgAp6mh17DCGlroqWHQhWkXHvsfp2c71PEI8tKI
zAyR5J7t2/yEqKUIzJj9aNz7CX11FJbj4yBVcm3Pt0SRZEmEm4QSAkKH9xzJDVxm
2kgjfgT9wh5+ukjOeWrVlx+BuGY2zR2frPX4sNJbYYBqZFDjlS4A8+TjqT0a7SdW
ar5s5dKiD5Bt9pFmLki4ekpf9PXmm3KYYBtdCogndVn0u/aPyzC9OHC4t3qyLrqD
kiiTnhpL99BWy1pbQh7udTvo52QV36JIx8i4yZjT9ezfBfeA1kFQ+36mGsWXu1FJ
4tjFh7pFOtOYvBnR6MLSMqFEq+1pnVbNX79V3Acy54uTdd1IpXKxlfHLInJHLKbf
x7sAw55+LGtK4bJ9yrXybDvO7vnMaZi149Scj8OIo2/fHlPh+YDQFvDgDzqZSYtF
McJzuu/whvIgDzxgEpQmEA5aDXmIll4Gjs+lbNIk0SU5BTbGcbd+xSmxRAj8wUrz
hR7fVdkboscbIpvkpDz97GOqMHuHdDYaggX2/UxPZ9axMTHWx9ZWaM6tuegHXXj4
bEWG7gXE8xL2KshxXEk9BMuFQW+j4Ezz+Wp0c160/l3+02G5booT9jsWXEwvUTXB
iasC38LYaCQEMrBGHAmCRwrtgeevFDx6uxrXMsWV+1kG7HFDI0qeNNR8dRPXZTaO
h5idrs9GeQk0UU9TDEkOtpFpW+vbh4MlH/sJFJBbY/ZVaKb7G5bFB3nGknbkZmb1
EmvZp9YSiQxVTtCPBUxr+k+IAIf+5eQzYlVd6MDITJL8LEeUeLuMJqvinkc58oPy
wPtR/GqpUIozkk3ZeVOeoxA8iLxrUurrq2s+2Ch3NK6HoiUp9kZKBcE52eb+IG/V
mQ14/6TZtRxXKMHHK2KHobM45Jh7AJgND9Xy0OSv8L7iMplKnHUhNjotmPBJ9U5a
wvndHHN2RrdpYcv8OOhfCE5I0rEciKAHJr5JnWwUK0IJEXtVAjFJzmH1UgX9qwMl
YhWXQ16X5Aw1oBPPg4VVSoz1FITDSWB+vw8u+QfDTZz1PDgbpx9IS2/cnOXuNEN1
DQh43j9SxD9z0Y2Yh5pY3+56ICOxgNDc7lgftRlkh8WRa2ZbFpwsUelY0NgcBv7/
LdNL8eVv4k5oXdY/XZBXg5TraPItIlDeGB5cWKTKZO+xJCI/4/rKoM2Qc3HqTca6
JheV5Dea38eXNCLg00Igdeujnv4D8etB4uOhsRG3REYCQO6b+0u6WygsFq7+3lCH
WrbA2PAguxGAt6a0SeJ7SDOmmuWNUUTIz4t4e9MdosQDDHtpk6kvMQjynTFvuVQn
94vHlXxO7CCJ6PbZmY+jK0HvFNZjziM7Sbbx7uDlGgTvMXXSEQEQu4TLdT8fqHuJ
ReJPNWVPNR1hPu8N2cDPjyc8FEQs8ZNpVlToB/94VBzO5xlH6nK1kNTyXMLPL6ki
kQ/2sAJkTXNPUNgGylFTtQI0lQckFjYj0RONbfgSZDleZAa4cvWG6cCatAMtVLTH
cj/UoM91zPRfaMxTeBvG+wOsjjBDQLqK3j+xK3BvgScfTi6wDBwsSb5W92oRnUU1
lrZ3zns5JUduCqUiOvfOR0GoIHWShesN+rx6Uy2US73vXFXIE2qi4CVAFPbjEwD4
nWXNr4aARjPQe8XyfOqyZR2eIKsmLXP88Sl1olG7q9mMOO8GOIx8z62x0/PB6Bqa
+inW2pwPlgsDP/7ndtgCRr0iEbw5gx+SDN2jYGlcpH4pJjlTeI/gxV8lubb/MQf9
ky9pff4B8bJblrc+MKBa79nJwm8j+hZyb3UwoE6sq9o6haHo3SU2yyCNYO2llaDZ
ztZ60AR7ZecqonUJmM8F8NikTaMgud8Xj8fgE9DGQxXnv3BF0qU3Q7UqBTddoxd1
F9yup/Q7kffoOx1ceGGNZfnnLVbzVttxHtoiZWof7eaxSuPI5515WOKuiAk/QsPq
uxwwmSQUuq4FPSfCN+2j1XbRqUWr6RsrGxFxNBZbFkfw4wr8Tucpa5Q4J8Hd8dcy
B7jXmWsMLBLQR3TBul48XyWg4slaACDofSQteFvHbWnVSBXKAEvEpPLtyHBF+4zW
C/ocL5irrngzfs9y2Xe0uGbk+MZYUnS0bdAA4QKSeMQ3syabfUY36Q9+LsSu9BD9
CGKTGU3FASbx2jQ7XedXjSfA0Vgendg9sd5ITi6KHkrmCTDBvy/agYMMdboHZ4Zq
ChHckXCEdMFq7Zrzhz0jUATY9mvFV6RBIoZAOw85LFoKavkrf05ZR0jn3g0jtCgZ
JF6OBW6C7f7iNxWYl/hvbT9DDRVA9GbJW4PxvzVdExArz2Rv+zx99l273SKYRmXM
80jQHfTBuEL4+Qf6aaCkhQwOClc2GqtVslRU84ZH2BLvmZ/FWo2Z4cVTFDLCRvg9
bUY1TONGSoDjpArptVIjEv5Kg5KPv4DdE88CaQjEZ/VJcgE0t4NqOXN5v0y0q9f5
ePQo9//BDdrNl7lV2G/SOEEXjIYybPTCYvcK9WNcaiYSUFUAsLjptnogvoE6hVCz
pvPSaB+pqmq9tvsoNN8Z71MM/eG0r+zpZFLRLzWyXKSIetwuzgKai0rO7MgjIbb/
Nyzg7KCIpUh13VRQ6unjGDpBd17tmlzgNbiM+7gKhLlal3V8Ez9uJh4BkzQ/7Yax
1GPJQL6xYpsry2fO8fiWeDcY4x4o9aiClZnTqQcc3K6WU2JYcJIfbfJXjP94cM/j
j6u73Fw10uK4SQX9tLSmovXPpACa3ljNMukJ9bfGR+/4GO8SFQYc6D9zqXkmA+2Q
7QFb2FJfdVQ8NsPcoJLW59xgY5A5QSki7lz3gImVR4EywOoGVkOJ7ydVe5qS64IO
kU8j3Jh4c4a9KDcRaKWwkqfFZ+PDWAPCREBSbOyJBy4NKmTHGDW0/s/n8QOTeV/M
WvTFGJAbTcVH+8irdVKxQW5kB8ZsfezsHKsuHy6eEJGtQyCSfSJyGt+MBxotz/e+
iVY8iwHRRadUvSmXQ6t7X9Ef7NKu4u/EVmBLMLsHJNMfXfWVLPeYfu7c0Zqd6Us7
+WDLjyEZJkB/zsmPr1NxC3uNfVChU+r0/RprtNaJeNjUsJ8vVBsMXCfB6lFyYYhg
2U7wPUaUMQh314oyVW4J7HqJhwOpiyBf2I0h9ATZH4+uZU0wssa8p2as6vP/9WKv
dwlYwpgyQG29pbTXlxjjFufQIxzk7sWx1Q0WO/f188zXsuYn7SZxTg1FlD9lhRgp
RsbwWDAInKm3QY5ZUisv8cL2q03F6bJrbIr5W18dBoqFyyH6MkhqCaWdHAQfGdLh
vjCtZtRhvxTTVX7UQ2eUDZrKEwMh6ylgIGleQXODLIumxfqkh1gjiP2pbpp6JbwC
gOZCzrbojlI/FkGCW96e7LPlR6htOB4Fzo7wyuBaTp4Pa+9Q3ff8MRGUeI66wB3A
Nih5roSNZTQr2IPwU5k1fWXuDxDmWTOvMmfUeb2h0VUamg7hE8wq9CvoJ/Yrorgb
Rt+BXQTyRmfFJMWr9Ht9WnaqHy+LHSXkzB9QsD60v5dsJZ1UP2TWTPxP84NH/x6Q
6qr1SW60JhJax4pxcCk9sH4KU8pNmD+jYLOrmdN2x5Mtf1BE/WIlrIloKkaA8TzM
CVCqEIyDjpL+lR1ikWFqsQa8Wng5+7/DsmQdTSxjsXfnKDVq67qjIe8D+goDhfYi
ONtTt2bMy6qtvc+/yvayPr9z1y9BBh4XQbrC83Vm1rKuJt2ndFTkiQQRpqI6KgGG
2XnSICo1NN/ZMkJRecq5QZv3U9RKTuiZM3eY+YgfqzkVbvCcZ97smqMF0sKPnLIU
ujMdArzKRd7sNWPEGOwD+M4CfvXeVpd5FjFJMKWOwnoeGu4QTUfmx1NMTCUaO5lc
OtiMsOb74sD4sxFby6JI1Ywa/PwPEw/RI5wORQzMIcNLplnW1YAtjhHNIngditjS
2AdNs16bXuPEhNoU6HHcm93ODeEc6nddcVcG+dB/My5LrW9ZNrYHri6Rosx8xpFf
7LF13XkXIfs2rff7IrSqxA6LTj96jP7wt24q3OA6aVJa/Wo0mbyZYH+qWhaRZl2i
fcMjGNLCp3tAak2fpzD1ReE4b9pqltbAwHzOYlxgLCpFZhM6+t3eQqpA/XQhwclT
7QPUPPtFlmU3z1VBSYgp3lZmOlKE9RiYTDPUIYtG/KWjS4aAcsZvXdaC4ayfiZcH
rt+nWanTKxUNy481yshlqNlKQz8Q+GRy229v0wZ0layHgiCrXkgLod6WLOvj47Ri
gnwSer5PA2hh9kaLRzNvrEje7RQE9w174Ak/QS2hmddw/joISkg/G1zvk58K9izB
EbFOJpfFwWbTYv9dFYsGbODsmFKGsrNht1DBKt+GgyESegQJKe1Qdq/Xqf1jkS5C
wf0R9vASEy1KP4+0apw0I8ASpBycGIbFGAV4SxjdfmISmV67UtJ8khAbUzmEbPbi
YhHu2x/92+yOG1b3ZHbJ+ojEcSmDjPaeczmnkDtmdgaaxfbt8ZVgZujOdyRW4mCy
TYzaKpT/oOwQoBYafpNZEDuF5n8ffq8OO/tP46vCCwTYmuutnihIS7UtjcPJFbzK
TOObqO6dwVVah37fpTFxN3r9x5RJSLmXixyLso711/izt35VNhp9mTeYvUC3DU23
ulSOCauh6gMutQvWMYaZoWbbz+sQZt/PcvfmJzqZ41G2A1LEIHR81XZdinjzB/K7
PZpTmrsMdhZt9eSXEybPiGUvvbjDbaaRTLoELB6oUvRMW/CWO0bbHJA7XnSIw6MT
j333sU0rQ+FMFvb7b8urawnpzMKTm4Yl6XZGtkh/0wLywTSBnBqNqxAjrHlJCjwd
gFwiwT0pRy+dDT5e0nKleWUHkD/mcyZNPbJtQYZ90h6+wd7/XrcBYqjauGMfm/J8
9ib9896ti6Fi2Hq2HwjlnJOpME6pvzqB4XECPGey/3I0ax4JYDyy9JRiXCNL6d01
RVmX2/iUE44sGR13IG9mQ1dS6OGhyRNjdH++IEuqUUFt6GzxgWmKVMu9ZCOxbFng
O38K02ZQRW1z4xZDYsP8PYG5mEhcSvOSZjuK0pAygV5h+F1B2NfbdUiJiXi9HMtw
NAfkdGwPisg777qsjnreeUBe1xR5cRQWsIJxfZ5kaby2+Jhyd4r33tHbWVq2KgKx
wd8a9Lj0fNZl+axfvzFQa4MXQz8wfG0ZIpS9nVv4hYeFIHu9XPdWfaUWSy+f8zFd
ADJbNZAmcZ4Wpo0VgjNGjXu3/25ZzSwSxQ7ajATEmlBk6OPTspA0XOb7lNEAEUqP
gsaUzJVeO2ZjAh7GapgqGqy1KhuTqTnU1ccHVqs0WLsckFyv0mfk3q0eGTZlZu6Y
AsxL9zbZYpW7K9vEyPEUjxqKVMzYnMaqevFO+LUZR7zfa0jr9AjNO6S2ysp7eihB
rfEvuMA75N/bm4Yh4JotXQYIWZwVrV3f+tTWAVWYiDWu8RpV9u83hNZs2kwFKQpu
oDAYWXwwVKRDEN6TxJZCK5jyj4ipEHwvwm9UgZIb5JZYuoLFGjfzxKbcdqSmB6dF
Wu6rSljgpttAcjad4+uWlzJPSHKZScJ+Fm3nCCIOEBoetzcyt4mJ8XI+B6eZXY+1
wD6P/ZGcmLWsUXaLUh5UCJjFoRu8H7WdJrGSHJxiiT3nK/pgQdC3N4hpzpytBOHV
1J4eNkfLi7FC8vPWcRP1c5mKcWd5CDBZkJ75pm+K0nCvODqSLeGlKyO19TZ3MlGJ
pMif6i2PxUmsZcFA8Mmu5ObFnJoEvL9yHGWYhvWYkXwSJaYbMlsN6CUfBnWOZv8e
QDhYvtKiAi84sdvVDGgfPS/07I4Pf8NC72+mcuTuGVEXbNMQtd0ZI8ulx6tEE0Gg
/g7FuHaxHVRAmPwoJijefleqJhHgAFS8HSktxoeeaNfVk2nLfnBHspiftaQH4Rni
uYnkhi48j1voWMzhw5wLL742aORqMZoQ7UZy5OuPcpXTgYJJX3djhQo6+PwGZTlZ
4vk/PpjFBlB3S2Rpob3L5eDZevs2j36J82WJZRwQFcrFuHliFmJqTFRexAq8Kr7z
I+sNxHqprpCPZKkz/9G0p4UILljFvGTObaY5Im7+CNo241DxKnmBg9Bk8XMwPfxM
tw/iryozrG0YvzqJTohvSZf6wyR4fJH7QAPrmwrrpXwAndbrJKhwRvO79yuE4El8
vnx9zOEQ6KatWlrCy/hHwyB0CKNrajD5vZ827YqSp5C6DvHB31xZS73hqDSeMWrn
/GwkIpgKizqIq83PUfgVggplav9n6crVELnJ3CvEryxwIzW+sYrLHrPv4pwGyq3a
4HR8Wa/cJ1TE4GYZmy8pIOLJhs+bTqQ/uYMKbUxn8UcKd20TkEGRX/BhNIL+hGJ/
b70hGu0Myjlf6jNIJyiHkVBqtFPB2f/fINRWzXNIUtr/JfZ22NN+kjSefndxd4RF
NTvonUHbqcEUeTPdTMzro4adJEbxcUlAhnXdM+vkEWH93NsRPfk5cpTa+u8AACxy
U8huCcz3pwgJ8axYTxm4EjPeLHVluZ7ZLgljQvuT2CmwDuBQ0fP//X825yUojw3h
6A0UDJJ0iu1k61ZOJ1RDr/rri9/4HgZz/VtJbsEo6bP7um1dmhRnHX3T+jgVHDXX
uph30aM6BWNYNyPC4mrA1VyAkFFRsSDL1hNESqSNZma0mdFY5ty2wo1eCGpMzI57
I5uI4dDQMzkw/MalfJ88yDOJhWzuJhnvFMF8nNdxS/gle8JXoYq9rDAJThjKY6sj
CAihZmmTkMwHvTJ2k5KVeA8xONszdnUISrGRfZHOhZ8bjlGnqW+mkwUo0Kn5siWr
MFvE3WJgub8bvt9UIp4ZqE9NROBMjD4D0nlP40RbgFiqMtKsdEyLhHLADLIjBx8o
QZwo1ZMF1u2VBf7G1VtQ1VVfUaLTuk7gyCVzC3qWhwc1Kb1O3HIU2pvNs4OPjBtl
2o1sEx6rUv9UGNd5XxTnnmKKAmNH9q9TAKXjkofkrm8KHqzwvRkIN6SkVwCg7kFD
7Y3oworcoU6fEqkwrI6N5zoPdNbyrcfDhozuKiuID5vJRIsH+ceiZ9yWD4FmZWI/
8VPLeFgirhbIY0g7a1IY6RSj6XLjXXZCT54PZKny2q2JCqkRaFJEaQTh8L4ju1nk
9d4bphKqrtgk2VYoaqRAXjOBySkq+Ixl5a1IOO7oo5UlHZZ0p22hWZz2qN0gVDRV
AKoeoor4GijlGGnCoKs9N8uE4RqsDxfXE+fots1QKsEr6YetBbZKuwkR9TH9xQuH
RJ4g+1fnKQWqL2xsAXJWG9KRRgx6vk0WbPRlg/FSHEWt3fB9yiN7tl11aPiLQUrr
UCI7Kv7Iri06fb5x0Th6GkefzqXOFTHfwNBE4Jp/b/AVWK0rGbpcnzNYjwWtHacR
PBRnbE8ThbNb0UBoBb7XoZqf31uc+0PwPfluK+A4mjdO8F4kJHZo7a4gW2Mjq+zU
MYy/eprM4m5fAxfC2ur4F01xfXQU3VtYQ7AbDv2b4rOiNGn5Lxb/Bi/xQcTIBa6U
iAzL6qEwapiZVuMpWCfKyY8KftsWS+ZGSP7vpunFYrga0Y/cu3VXtQLjMNV7BRG7
wDW3rzJazwV/G+O6eMIAhBEJ/trIoUE1nX6aLpV/0dVS6FC48ROdh+NopcCGnWBz
K6+84hXx6XDjToRcLW7oeMsxNEljRnmtN8Yv8NpJxoA99nQm/MeA/Rm1mtxvDYel
c90rYlXTlLwRTW/k7st3DxiTvTsT9y6RZyjRuYR4E81IAq696ESn0eeZfsWJ66fT
NCxy+ZQB47eHzrrf5YlcubYuKFFGn15nDl4XvfQQ+QL+UPUBK/F6D557zUgDSEeu
nyNBD+cgQD1aOGq39wigG+CuhlLjad4QXvmDihwmcrSm6M0HfgAzlXi+fIHvg0Js
CilIBrGeScKn9QsJT2or4oqys8hAX9CFgDn6+VZTSgwq60/FYXUYB8zsjFAERXY1
pnis3Kz0Q/4RsZGEbieGpB+wnzN9n5wYI05YKzlG1X4/fx+WlZ5a0yH7XBQ5BQsE
xOQk4z1QnjuDe0JWn8a/5w7luv61TAOZxte5ZZw762wMQay2wmGoGSTSwSE/PoFD
yD40PSwNeOer4YN30FHkwGC94dIPU6Mo0AndBvmtIxS4cdRYssliZVq78tbybxr3
xpbq6JVCBToFzFCPA0M2l8UkC2e9q5jnV2kofkcSh/S4/ze9XDnV9FopRpoOyK+/
hvOea47fAkHpPHbFrtsytpDW4FmgzfobzGfbArlm1eM+9XmrR87t0vM9/wQRYTSa
DICbrPPFVnUZWbJI0tt9Mq/pVhartKxt7oyxm2BpbIc6HkEGrL0FQgAjDgIHl9Kp
3GbkThpi9nt5/xg9NsLm6Mz2mdZbFIok3NHDPFBRggQ8ChNU7qeIEXXvmqy8qF2i
pMv/e0RRyIAIcLPHiHnZScd+yqwD+UyYzGqCu1w1zDm8tjJnGErd/F8SpUd+xLsE
Up4Ji4Ikib0WLQxbRaISjGRD5aIiwWDbJHNxUg6P4FUheG5Y32S/HRYC5Z7YeivP
aDSSSGhlwGTZ4KfYxdphIX9O0htMDUFt1+ZkJfmkZfW1ZuOwYFzKx8UlclcoWFmj
UhwGtE3VGG+CLWzY/MYdYXZrnM1LFPsw2TK5kSMdqWe7yXa5Yt7heh/omMyHgtph
DrKlMXkJSGdT9TuXb+/0zVQfslduwJwzPWunEwTZflJ+EboAp2KpEANqkXSZNZJy
VBe53aqzu4sFDSnuZywZasFIXUYlbfIAkw5BsFLesVei/vOVozRUO46AMaKhDn+v
vfGWzDvjCo+KoWdcLKy9tVaFsspsXCY1eHlT5rtvbeij1wpEm8lslpRUtxee5Xf6
YMcWMR6cPJWf7ugNKtJWfI3jBCXfW0M4caexFLMGAwvq+D6F/nONocV7WABp0VVs
1BRlJLhkHgGTzWjK8EWjIWJOaDnYyh9jBPPf1NlbtyPSoHFV1lRzqFdKQtoFvCq0
kah2MA4Nrw0QFrI3XzHFZ6PrNbNgRx6/xtXozJYv+YmIYUAZ+zJZgtpBIkRqjwLU
aMOpGEbe6Y3J3Ux706fJvqc7D39kYKfN1p964+21zZKFx6fJIqCTM3o7VEYCG1Fa
vN+QgkVBcFMTZTEF8uZN485bjUJRBQJ1UwalVKBZNRPFdv31Legw7/49QRPcU7lI
ygluL0Qo3fC4sT9g4D/HmSJEDVDihH6KF4JZwAATYuXY2DL3w0nSws8B1Soe6Iym
76bps2oE+k6OvSunpIscyPiajU5AwWwjHVYHWE1Fts+jAs14dhpW85qU5RZlR8lz
mdXov0FruIQrqhkmVxF8ErCpKiRhrPwT/+YUyxPjvSlPFpbUVVpKjo3Hl5Q3Rn+O
xTvrNCqWKuDMv/YuKoEhjThW4rkdLpykxfrq+7rc5QjfkzFRgExHDLOyPv2NpFvz
AzKAyqjJJGZqQFNnrfC/oIoSxfFBNMT4Yc+VXtc/CgTyCLrrSxXB5JAtJXxtr833
8Q2CpiaxwyNHvKpYAD7vbNVy6nuQ5PL3+JNV/MHTO0bHRd2w6ArB7rsLrWGyjjjB
Tu0WT9EFgVuwBl9llKJUU+cOO0xOHy1cxneGp6wtaXtHv+GGTs6r/e0XTJ9FA9nH
2GuGDdOy6cxE8ok7sB7CA+5oulZQkbkLoV4uzbGrtXpX0QR2TfBF3WdwYffTS9E+
TVjS5bpgW+xqm2ONmD8tmwqmdgj2mLNHLaCJLIdesLmLB/Vbgd12QH/Ncse3Y5pq
jK160/YQR1EG8GpgA+36IOjv8TP8NyAK22VLq8OOxblnv1RbROkVg2oPMyqcp9L0
Vj1ojSIWX3bLs1ReM5PUcXMAgSqFLGUsEqLHeJpoNaJ7tBEtSCoS3TpItchWKAIo
Umb/26Lww7GEzhtM5zM7/vy/grjBucCVqXAn2EMKkMWqXticB3c7wNvTnbR9FTdL
9bwdVE1TcDnmcPilYNKN7ERCQ40EaX+7LmC+7pr9ES+DlRgK04UpbCHQNi1reYpt
Z+z3sIcf2edIkw1fg6aKAi1BWEvke7/esyzvDYS4FrklXzd9HcS4Y6zd1bw75R0F
WTy2rCOwN9cexsOvWxegqjymvdPR9sElYsUVZM0IgLP90wlwngdHLjsjOooYIxHU
SA/PoYeZ93j5BvZ9nAe26HOqKTcGs4gubSNx9Aoa8tCMirDCH/BBvIf5Ublu6E3p
/qPt0AIVXBeGN7Sddv38pzm2dtJ8JLTSIHk3QCSsUABxJ4ucscX1TfSe97fi2VqV
3v4oqhTxzOkHkqqMZjJpPv5Z9vWurm6B6Nx2Vmne8St73WSkcEVr0xyXQAfLM/tV
TUz1RgYLm61LQdXjakLRAnCpW7CZw5TzV7Q1VJXbnjF320SlAeH5sMp01WTXONOZ
tseZDYqB6pWqT2TX9EfFclouL5hTXesE9gV8tabnrDzMhDvHbMW1Zw4/4j18rYIi
WL+RiAFCNe8YP1JfWokIIf5Wi33Gb6pDFFsY0XTclM6hfUp6naSo0SmTS2Ms6ENv
Kxs1oAuN3y1CKVHUPKfceoG8mEAgzBQ/A8xOuTGfnXEECfL+6ao6HlDSNfuDklOx
rdB6Rt724gU3xb7U6oEWGW9FoxV3QBYlXboTz8FB1RJnJNXJkAQ9iyJYFUOvHK/J
NK05Sj0207wr5fMT/wSccgUnWDTFl4toYJ7VCIlr7S1PS/xVC8dnxrCT5qNk723R
5i9DIhPPIMf0ruO1NY8gwHzuhRph4gnG/hVJwF09o4k3oppaQY2dCeBx0Zbu0wJP
Jte/RYGKI4zqjMfuqd3KaQJwLQIT6Pzq17HBfgCCUNG02wCNNazOK47n12MDT/Ki
bjP4Z/9PJ5NzjzD1kuGdl/hYD15o+uz9ryGILgpWnP37e+yyMtpoifAvbar82Koc
cEzwwRO6oq9XzqEROJpWIcb9liMEsiX2/BtOXJpniCk=
`pragma protect end_protected
