// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IgfHoA4DxYodirmv3Jem4xL9EzXjkKm99aroXFara6NIAMNWNoYw7+OzonddIqkG
Nvyb1opOuLK6EZLLX4TeEns+QLYRZM5VMsY171F9v6Q7ukOTWkdeuWZTL/u4r3SK
9SsJNGX8KLpl8eU+wLEq880uaWLZ9hhAJVo4TdB8spE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
Tl5cxK9jE3htr0qY28gUD+6Bg7PLKNHgY9uTuHJVhLyaWlpCo5Wb95Jh8456OSdz
kCUmqxJgQM2Wb1hgqSV12VuRApfBwjV7YLpAKoN/uFaCIjUlsfrA+Dsq/vUrGyiv
dSErgheXSBO91CfFzPzkxvETa+Ii1nPn5yPgi/ZtryX8Ba9EqPKqgrJbHYfX1SVl
lCPVe3oKeOLnNKStayO2ruc90PNHvaHwIKvnXVwvFkhKRRwNdKqkBwCEwkhk4qNL
0jY6M7/V4T/m8wyjSN3EKfTocarNED6Ep8i45iZ/lcA7jzCT4GDNAOrhTHMFima5
k7xYECdA/b2/e6p623Id88hQEUGjbRPFARtsmn+5/zxmdHnSNbSJ8q6CU3wXz/hG
EABc4bI2SBPWGC4RUvWU6hgWMXinSHILvxM9RtbCeMgGcrYc04w36X0FTtpdiTI7
Ja7qWhLVVLNZPcLNvvbtvwvl9XLDf1wDc9jTkG6p5wFUzynv/3dY2dk53rFH8Ask
GE9knuWUTAPHlZWFRSs1HIIqvE76nb87ZOfcqxf4JXRcnAOlMlclzg1NX6AIeDf3
i9lp0JAgo+OZqrUw69GZsq++W2cJZwK8ZB3I4qFtDeUQHwS+kLMuzb2Fu6BIE/IG
NVQfslxvxHj+GseUArJ3SrljPCBEKyjVoMPtVEwHioAIi+A1opFNnGXN46OyTpOm
WKkr5466mAcYpsafZrEfMgs1WrCnAPE/4QMW6gpYgTFbFbIu+G5gk7yCDaKXAlpR
G6YBHYVagChL8NoBQHonOzBDM1itfl4dPLcbSMPNPLK4CWB68fAcnRUB3fWaR0NY
C8RkM0RlaDCcgtwoe1lPqwGLEsDW+o7AuTI3jf4uys5EF0EHl+HVvu+lJna2sgIf
0Du/ehfrw5zqqRoj9DgDfT8YkjFfVSlw2kOZYuftOK2MkDkbjxqz3AhWSICY7YUX
qYbM/fGu+mbEEUuaFRvQwoY9P+euaEpbfQcEuEvjJtU+cXowYgKrjgNo83hWvFy8
csiFIPCfyBm9fsc51c1H7rT/LiCIhSc+8zDJFrgjD6fTioKdpBUjoRL9OVSdir2c
wlv2EEB7gUhDMChrOohVscB32GLtdKXO7ZtE0RzSv9rK5Fkcr1VsX3NnwroPbV5d
7WWrbnzwhz8T1pW7IjiRBdl1zFKJfvv+9pZnxmUyRBgBiX4Q98SqXrBebHUPM7gu
I4zfkhgMuvU5OXQ+mwEzGNc1gGbDqxiOE+dQqy6s9qeTiIIaImkIQnOD2Vo2Kb8+
SEBrBIWZ3ALkb/TQNbsBJRwQ5TYPrjdbIX5K2bt8UT6A7cTj1S2S9BrUJsiCvV8c
nCuB4vbJJMVyI2AqHgUpROBH5DIalq2ih26MAE7H8ttjkpNb76chyUZMe1/Q6cJZ
tRECljEHSUVDC16uoNtU0LWmZm8mqx7rVuEYCfKA7FIGOK/Wq+gCYnA+peHzcEBy
+JLN0qx+14lVOvP+TGQu+1poM/H1D9qSvFq5SKdM7P9BxXScRuDPp4Y52pPSu0Vm
po8Ic41iEjHiGHkjDs0C36S4AXuPrl8Fj1Yf42Mt0TVUhN10eQeVkxED3e+84AQ3
2cQvGEGAci0Ou5VZWYmhibYAVCMEvMTmYW4rEuItDjuyREn9H+wseFLMo7tymrKw
Oxn7HGhQWGPheq26evAwyGKRn3+BNh28cGuR63sVBhyyXL18g2YDg4BwNpJbVNO6
G5clz0PMzUK7UVT34aNd/Q9OpbXRAhq95CvPNHbTtTjeCZzpt5IoDsQJHRpSItOq
VK4NwcX1u1tZ2zXZJw9rV/qMKx5unpA3dwnHGBaxmKTlukl0VOVu05KDCzd+N/4f
bXXX2Fo5KA5b+7t5Ry2+qK6zpeVQiztp7hosiZZbQu2nHUeb1mActjhE/pNcbi9m
Gsxti/k/SB+wzb8gEEpDiv7H6ITTRo/lFwfQuvL6DUDhteVmRdo0cKvGVRqxi7AJ
YkBhI6CcC588DO+us/5oJgG5pj6rmQAuBrfcEDdDIsn3CaWnUS0HmyjZD2FgOrNC
e4yh/9/asnOc6sXG5E0gnw6SLxI+dvxS4FzDzPyLD3g5JErow3Vdc97SRMF3iPHr
skrI9zQpXit/CAINkMVBw+zCM74ERjGnr+W2+3L8I+GDc9o5578rNb7ibQDVP66h
nzGN4mRwKIJb7N422Dg4zcUjPpW2Y337ZNyDImt/Rz/ENSgKgtaLMT2NOceuGsA4
wv7WErXrJYzCOqOGy9fljDMgX5r1rjyP8C+02WXBR3hgpShzJUwnRJVCQMhAND3H
sfbkFFf3nq48pN4BEjRRxNEGDikkoYP8DjrU3O6lwdnTSuWgF8y6Hz6A3GvOLZql
/XaBb08kVb61iCaRTyADk2vm/haD62G1mBbMyTBMLfJQSrSbYhV+hosPCxh6AyPK
hiRTb/hkrVu9EIc6wWYQyXLd038U+OO6uRWdsLLVpALe6pip7e4WZPndMfh2rrCB
RZYhsYp+pnhFM3nfF3YfNXCBZTeljfmwql4He9NOEV9bLEQ5MlwcD1sO1e8EuF6S
ttj5vqVyeTeBGaRl0zF6UT8yu4iBNdWDz7vsNNChvFlIZ/RnauEglavJAnqeRCWc
JW55a2vv+Kfsua7HUl2eG68bETggViOKIJvflxoZwubyJzFy+mZ8eASRepBx59y6
5x7mOkWfkUbEmZNIpak4TIIh8RwZdVdt78nED0L1TfcSLCkBz3TJle0OSoeMYkBr
pJTAzxBFWCPEDGXBZvY7LJG/lO1bCSIHJeG7SBvhA6fArB5N0Yh2Zd4xPqK+4xGD
yzvkETGTowuqhyPlHYJ6tQ3uWk5BMYc+3wxN61JI+tS7/Tt3MwI5nqMOmI9G2gKP
BHRSmXOrQzd1cc5EvTSoVKCAgxdJaYCUX6YHWDbhRT473k3Tt0X5lvhPMGZVCGKs
fo7m9WODHOolI2qWilHXsR7jHqVbudysifKGMaI2ScAy+UNgzb7Dq2loLtP55Ux9
9rfi5oQ7pIRUcW/d8jrF5T3bSpNgi+AT6SH5xGMyP/KH3GNuj434D+F3znF2Lk0f
vWGDTIktMu5vv6jzzvBKQoF1hKKcVJG6jrzCkrIraxvEuAesfGwm4jZoa9NAfxsY
X0vdhA8lz4iRhAPzOA0K0LrFY9SWG8PUhVLmA9V7E9h0c5kPy2ohLnk23oTuQW7/
D98QA5O1HhT5jxFZ1OWFzKDNBjkHElgfCXgyy+2QMVWODsOTmx88cg72nvPsuddN
0hEY21Nic+PXxRhLMV1rEBroZFj4kjHQT62v5Sc4bEywAFUmLfBdMp/Y4zsKT0eA
vu0trG4ZC55GfbSHZNozav/PzRuTU2OVYAD2w9SrO/AI7waMM9jl0QCe74TUrU17
hGSxId037jBfBAW7pKRvWoVQIYfg+6lAWXuwC2sFGVqRRIk3UNn3KaiwlK6Fszfy
wprADNMX6d46+Lgy4CHvyHwohqpemgfnVH7Jk1vdAd1Kacjic33AtYgMyoJsGlhm
17w2r7qqXJ7dGgq6wGMOUMytb122LfocPzdyzXpxQ71ByJktGW5xUvuO5HDWigms
QFIvT4qeMH7c9D8bBuV4ii3VBQa9Bq2d1yGlCKO80XhbQSedSieFcbh0G6HC1A0M
PhV9wLbBKodA2AmEUhX9kLlSVDbNUC303QTjqnpZlRQVo2acu+l7w7IDRaa5ZjQd
+bpcFojFLAoSDJH46PeUr8wNq6U7YJWTDIZXvLi7W87n8hPo/ybC17HNIo4TuHOl
LowYNY2tV7E7RwIhnSq3JaUQzAJ2X8MZnwDv36xriFvKzJqKpQoaFdMEkv5pRElG
vhaN4T1yv7feRsBRqCNp2kPryy+Wlv98Ol7eYQYoLoT7JQVQ/9Cct3NHfYBn6o8l
nUnBDMI2j9cNtyXS3f6crScd6W5W2Ty6StFdkMn6cjQAuEQOKJeVbwjSZ1f0+ZXr
MPJK+iy4qJfD4osJEJIPLzg59OH+AD3GsWdZrrmff0/4vSpjmqskgyBWsac/xgLz
+B86cbAysKzZsoWYNwCz3h+/2J3bS+gh7fmNOfO2+WSvrStoICm+SycyRefrCLWH
ZTnx4JbOljq3z7Vp2Wd1DHq0gC3iJjG3MznI/Y1fHf7lwpkk8u7iLnc0CFXOqXc8
QWQ6pClmPim5XM4ONN5Yh82IBxfZsv2kaFIRvcadjNI8ytp4C7AnMlMW+OQPPAc9
kJP4J2XJxQQNW0f8HXicKN7x0+B9Sa0PLRIyrTOJxyAHLSnvOQ4J9pzKGQWJRHuM
jGIUaddfsieYItVVgvSDVBChe8NYTO7w4+QX7p4YLgUgpDIgQhXFCnkJxjVYkqLz
VxN2N6Fj/0mS9Otlsj9kdrxowyI2jhluBUT9iQmMBhxGtyE8msMIgHD6c8Bc55WC
AFmidML1sUQWsTS5L0s3lNOCh76f/laJ9MPyqo/70DuKDg2wN0GbPOMunJRNbtt3
SPDjA4C/M4Wz2TOZqqoh5PwS+CAY0UCgXIr4mj70yNp5dKeJ3ZCO3N0cQiMp3mry
8ILcw4SJJK4mIcnAdYtjSm3LoOR0s8/zbvgd4010fFECFjCNO8SBK3/8r0B5qE3K
MU1em4h8iztQ2Japury0pnoV2fj9CVcZebLAoBN1towXrnpDNr6CJdr5pyrD4hlw
w905Fc7mTT3HRoOMlFf1FqbXZ303ybW5a5X14+qedxlRGh4Lrwt9NU9fMJWS86Xr
rxDmuWng+MA9CWpps3JKlbmBD8fYCXZtBSov3MoGdZeH+a9KPxt0A9AdDgp0x2FE
LwvnXSKMFOuFuGY0kdc2JTMkqtRnwe7b+JPIMrLwNu7A/sMKGOfxbT5EBBS7emwu
w+h+kprVqKU6oCO+j3CEo9VKFyjFXB2IO30nVvOnQqr6aOaukRuXupL51TjwOSya
AmlzchGqWoqtO2EKwSBhCauz0lZiBkOazDQu0gdj1r2q8cvy6sK6sSxChqxYeJ2b
i+bz0j2JIxmKg8VaeoTjcVWrVflczsg2S7evGsSHK+YB0hC36h58TU4dpjVftqRc
5QUIW3OND+9WGQFMBxIHEc37cZ0HfuIH+OEvLsitGwd5hwHjvROIHHRxmAzXwkWj
YAuD+MCY6a3ieO3P0AZ1rZBnGhqFoHOY98rlFOkNV4js0Tqvrrr8FqDSJ+rudW7d
iKPNlGui0UcxdtUX5E44CYj46FclITnYDXfHOjmaa0aKXSbzrFEmPZc9iQU6S5q2
d75AFXbSKR3irzEpRRptjVR27mwkiZuMwGt1Dl7aA+oo+iiP7mXcXdWDkH+fUxIU
7GNMvukPxGDOVW1kdP5/iYlvVWzuFmQuR1qGAmYt+C+iH1V5m/9ooFpT347NHGqy
me9NOgckRFPDuZ8FoOmgkIJhFuXRVjkK9Lqln6hNeC/47TSmDqlXZF9OLDKzllgH
iohNGZ9qpar1WAhZWRPZjc4yFN2+xfEm5HsXrFsn6GwBh153nGwNq6tL5NhTA08L
hbyEzKELNsXfMAThPeXC93TM16qJQkHkOf/Ll+x7cQyww2oRlE/1lF9cP/4lU583
8PmtC7S+WIG+fU9pYdwRys4x5fAV6h76Q1oOaCAmaGc09gIfisolMa/BHOl9naeO
B12iAFVdULN6fUtk3ex8iS0ZVCFy+tpPgEp2lIQ7gk/d4HVrC4dBe68IFZNgF9yZ
VgvYzKd07MYlqvZSZ7oRVv6Nt3J24MxPjJF/7wz8oHl0uqgFFRD897M52g6CMImH
+EkFaq8nH4kccNuEyXAbvcG1NAVEsFqZ/F15v1pt7lZGcb2btkcsDrNzdVeGiGY4
XhdK82LtPetmoB31GWWa2ZTo39djfZC7sSRXYOmlmjq10lE7pmb928Qg8tb95nVm
FXTaJ5R/eBoa6CMvluanQC1uUPl13e13B4SGf5L6JPxFsl3JeU24ItPUIYYUuQrx
HDXeKbZ1G94q+Xr0DtVrq8gQxGG8fvS61rz/GphThcaVMPQ+6gpA4+fF4iFCq7Ae
5f6S7dZ+UdLG6P2L6PDEFH74R/jdDRXe54k8WGplXQsVWBtiqFrc55vVpMyb5Kl6
jZquQu6XnNTpdn4NfwcXLiV7fWuVA7oa08t3MZEGsOj9IAe8XowP+u/6SWJVcd93
Gm/MDm7dtZ5KoACm3mXdgP4WLWu9yEksZgvE+cnjYxMRKgtWq3bmjbGL9ARvaBI2
W5hn4VjkjVrylGq+3npwBR1ddXJ6PPNCik2pxRqCTRgFqhec11S9nMzBIt0PWpMo
H2nG+RbgqQ104sktWksxT0kbH9fymipbpd8hgu7qVfCE1U4tCGZKud13qHvcCtIy
vATyt4NnhmNQKvzG8/tQgkYrAtSfBExxYqTiZx/Rtn6sNTvoCWFQXtK9jq1NdxLl
2O4n+WPRjTXkhi6oIsMhw100B+MKpcAfh76vIYxtwosW2xFwn2rTlg9qW48OarvT
8RW3XoFy64l0Afl5L0JhR5IlPM6Iu4AbOMQMfmWvk4cJgHj1ZMaTXXPrumvdycPo
qEMxQ9H/XVzSTjUsOrPQlBdWBkiteu/A0sBcvI1rExW51EWNmAlmPA0jeoMAUMBZ
TJXIVJymUYumfsPQyYVHL6owsLJCUepFQ6pPJpeq1MRz4DIw8UD0DKvb6NSnhnma
MDf2WdSV17owN9Mg4/QsQHykTRrQLButSTMEo5yTWamxk0NPhAHdeHU7OFsxwLRU
vOQcxj5m1ONkt0ges5gkda062cp8MKvhHKu2oEMb5cWM3K9hESnBTuOMTQsKDH6S
pOQTry9qsvZlhaFn2BHaMdNGPmZN9/UzO00kug0aMsXpTtFqCShp5BKpPzkOXP7V
i3G4+B0COmDDALwg831mVtlLqlOT1cKZL+AcbY/01mOMs4L+9He/G676N6YoyiM1
1sCUIcWjLBlDyuFrtRrQ1vJx08VZPIMhhmvSNYLKeRjuRlUhqDhuIluWBLSb1ZY9
hfQH0Vp/cIN/z9pVRiF47wkalz23VYQMK78AwndmQq2pWrDlRLWZ9qLpMjdEgZ+x
kR4E/3GNxxJk1VQql1eH3w2fRvbdbtVo8IQIsu0mIkhSFIByPPZhgYKjdE13z9wm
ufssfdaUi8uQ5BOP+VaOfdB9bhY0uytUSibCcI1YzDX8Rya0TiAcOnOHMbWGF+hw
RYSfEYzsD5+3a9OcHM5n5ZPr6AS7hqTuD4cQSFH46AiolPiivw3OO+2MR7+7Zwqi
YKAvXd+eU55Fub0ZSHgbvgF/B8NrWAQsu/+Ie4onOS9rhnDSYE2sbOmmoC5fE8ry
MYpGCyF1HhHM2Q8nzLpJg2CnRIDc6sxrx78PkZFbjN7agfTk2Ekw+ulTzlwHLm42
OBLjBe59mDigXg9WxeEDzneowryP67rUYatEw86fhyhvo0knnsELhIksfdZtMvlD
/bfE8goKv7qWAgk1jvMxnIezCYU3ZHdQkZJt1bJT+89RUoTLyIFu3AuMtXUZPlEU
vSdT33Yeo9SRBuHH/sU3zxLfp8B8dggpa05pWkZzqpONoE0uxoOu2M1atGo+sSaE
C3mBgyJasLOojK3FKl0EzFE6O5fw0zwQsQWX72A4r4GuhUzmIqk8mEQ4XoAfIFQK
EzEygYx8w0kE3DevEAESaBlYSp+dncv4HiAcI2IV2yuRafbA1kHrOPgPkfm42KrH
v4nsY13T2QBuhurPHZfS/nIYPguTiuPo9Q64hJFL57mbePV8aW6XmEIllbLendLv
lrr0ClbSHbjb/I4dUVs6oE5F2ya4uZ7i1Vv1mSqEQ9goG+idpY3Vdp1db6kENXGa
QqtUA2Vk32Kqm/rFoJILCYePkykwVZdxAGQAmF6UEZiC8+NN6RcFu/nwTeS/Gfxd
IRHOgp5xxWjtsTDivkkaIc0YcwvXPocpsTJRgJHd1rQ3b0ri3Vmc6LQKOca103kU
fikhgeOCdffyOWMshUSi/HepaCNi8LNEngN+liW8eRmsU9KM6jvRVgMKEX34/TSV
8lryQf2c+g7sRviQnyrYwzNhKPrpKm2o32W4OrFaBt1DwV4YjRbtgovd2vSePpxb
reOkEQfyHatBtbWnVRHf62tdYbGeczaitrzH0O1D8SWYzYj9bLtrnEvFx/SAVNS9
P6wNSy666mPDNG66XnYe/aQDv5E1QS403UBCkzS4Cx0NvTVCOjicFOoz4r6aLpL+
k384DhB5e0HJpj165427Fbb2xlrPqL3QvJjeqopWrAIHUdwLIt/RDG10fDjU2J7N
u+4VChtgqGgLmkX/YRWroTRKaLmIo+TORDsmT6uA0Al7Udm5YIzbHR1qHwLxvpDL
1h5AO9Mut7RRn6q9L1RadIPMCJnxFMAGzmpAZvn3tSU9OkB1T4ANWNQtfD1z4LgQ
j6M7AC7bE+WjVzlWnR+z+Aok7otv09+EneUsgPemXLpiWeAl1598vBoJF+AegLON
sfISuviLWZcw4FFLAMfnEV/pTP/gxc/jWIo7DFCEEAoGLMcmyPEbi5Bu9KRXyj2c
KJV1U68jueYIOo4VOqVF9PQAWr5ZRHI5+aaDQTWl8MnweO3rIIu0JE3cCNEqOQAz
bfYbUVcEeUxojm11qYaI7AeeS8KGScoen1v5S3jCU05qDs/qI6OT3G6ivgwm3iG1
Vd/wajePrylwojx/EtwAZwzuTzyPOTacUWPCdHKx6t+D3jDH+Qrt25Ac3RJVyXry
eqEQh4vV8wIo51ZZF6zxozddCdMM2weRsfUKm7TpJaYLAjsvRhGCKJln74FgYLz3
gWGFrH3M1C3B7+2l+QIeHoxtPSXvZL2FrqOWe4g98zxdaQFxJKwdatoX1FRmOx9X
LjgxG5esnedwIU0gNtDhcks2VWiO7PtzW21iu1eawvbf1NAHa+zCPjMI5MYxs1n5
LSV3UpaO7+i3K5dcJudKrUTmFKkw7T7WCDGxIi5Oe8bZaa2YTOlF89cTwOguDfSz
K/bBb5s/LEREAawVTO4S84/1MJKQr0gWtfvj8IySSGAreqnXTYgq8YIR/JVn9Mz+
xw4TgJXiCiPvEcZSKIacwMsONkJUuIShfKY82YGa64DtH7yuH3A1a0VO7iLVcKp1
TcKcvvQtaR6QH0gIVkuIdwRpcX2i4YA/Y2yzU+ckiwPsO24S3cqsvZV/4UhYHp0R
o9UYD4aCcUCiyA041xTKootP+8f2P3lv/jr780BanvLkAepuUmzaCu8ZAsj7q4c/
5UvELLaSvZ1CBKGOjbuXWZgVqSNyQRh0Zhc4I+BjIffeqUv2ILDy4cnE76nQsQOq
K1rY3h1hxYOcUltxFzj7SdLftzuzAcxvz+0v4yKDnwbE3TUpsqmI0MnfEYcQtMv7
DcSZG3YCRrUj1WGgBKZ8FsE3YPLjbo2XhrkqkPqogWBJ23Zr90i24tqx/gRt+J48
ySrU2+kQlcROHhbJnhtHxoyGejRobkbZzaitt4Tlns+ppbFjykR1dqMoq8Ix+5Zi
eNaSkHqlwXTs4bAP5DHpbQgxqXe91zTmPSw4NhTbhheTyCPwXKjrxqYZOIgxqKgM
KMMuJlMRaZmEK9a6EyrZsmtRqZpxaj4rRhcDIZHCsETYnKOK4WixWRjtEf5mMOqf
UKN6gp8l8R0bMdhE4EpYXKnsSq8AtWnH8ufVN9ZZn1c56xMU7W+pu8yD7a8T8M9k
yeMPuppNPvcBx8R46UnkJ3WJJsGVusVr6+OkNEOLHTmT42dyNSYpMENghTq1SGuF
qIm/RCqCvL/LKukWkYjRTQBhMiCMn5jf3D1eoq4ThOKFKyMI5oMJwT1zLdq/Gk0L
73uH+uy8El1bvc9tyyGi+SOsBz8JW/8sLSTvjaduslOIKKy48NPCGQFY1u22Fj0B
mgkIryP8IvEng3D9Q84mn0VcehIAHIUDOiNmd4dWup9lRYF3H5AHeFSEy7cvUhli
xbyFpzJLUC0PaTNyGi0sryk/3/Pr8MhCJ1wOrJUntmAcKAZoyz7AMjmnNzs1ouEq
8WF/0FbE/Q54KNgaT2fgJMPdXvLpGqeoK/5CNXDK9HTK/TI2C/rE4uFLpchJgINu
qTxIgNKJHTFtoQDe1Yggc5R+jXnaaFg+ExcO3LXEYo9Dr2hZXKTUR7nZbbKQRtZN
h04aBqbEZwvxkR2BZ6wrQJ3/4GKMeAWW7pn8XeNyDdQAp7sIGHPPHc1YZrygyeH8
5aFPNI2PguvrAUro92IOwHoYNTZCtERUzF5DIkRFqg1drDj3VbWCcfGCJ+ND3CHx
HATF2Jl72+JNyVhOFqEeCe/9eZpk295qYmpYy2crqWsEj33b4mB1WPjRcIhvP4CF
cFsspkFrZVQWJ/6kEmJgkwcRTl+sDERnBZOJT7y6qUqmbExileHEca3PRYPUex/X
jrDquQk+Rzr2EIPD/ruO/OBusp+ZlxNaLq/FkvkBZQ5bzUhsc/9qaltXhqo0WhWW
Le4T2dyAs1XiY41QktQvAjbGDZhqNLPeHV6xGAzg24M2184+H8wp7T65i5TUp9Ez
D5Ixa7sDxC3tUk8dt70EecEcXZwjxpGdNxf+MIOtgrt+vvKoBdSJBuo48dJ5h4wZ
Rdqld04XqHVipgUijlRvHpoTHt9+Gcbr942gS2rmpRr4u6qLX2t6IN9Y5rwSn+XF
kCzGjsWtgg0nCNRRA7+JTgdg+E6fkf33g3gpatT2gHpDKtuiJol8FVEFNACRLrdx
XsSLzY2sO3kLuZGpCBAc/Nh+Z52nJ1hdlCjS4f4shsaKKK9N0Wftogg/2WzZa877
hIr+X+M9Ax6HjEqzGBlkS4m6QYkAwvLJAtZXD6mBCr+AZUrbhyCtLZ3nshHLV78W
3bZX0WhZA7y14CjaMEY+w0fw0hXArfhxs6capD53jStgF3gzzgQ4OeOHxdfIMRf7
75qTFLlHjCCUl421Bu9N4zNRSE18K/9xFp3Uja4o7P0wwWFaJUwGP4eth9bI12PS
XyQzW7l8a/niLRSEkHVP+u8EnaxCPAivmIhI3mmxpJX8a2kHXsI/X+smFK7Dmgpk
nSxq2vXuZsGqzYx0gx/faA==
`pragma protect end_protected
