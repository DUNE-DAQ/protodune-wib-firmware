// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
enS7nXHCR4ShgGPfR0vF3bcS7mbqUB2S1ghTjeGOug8S5dfX0jdB68mkwXvk1SuJ
rlfoftn0dKQPkhkBiUNLNT7G2LrtFzfxY7XKPXqoPx+bxs+oFlGjHSQz1y7FpnC9
356h/J5fpme2kS4/q+jOhWdofrpvrCSf4uTYohlLAug=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
qJgLcqf/R/NmVBLE9OgJHIDWb3tXrj6Dz1ig43+kvu/S4n+PcsvOl2Q7/nl2lQx5
zQdpJ1wXqEoupVrsgZ7z0U4//9xKYyHYEJM/SHb4eHUXDMpEgv6P9zd0M2ImpXHD
CIeKhfmCOaethTK2wHjY+e9YnVXATUMwRjR19DjYvzoTinydoRKa1TRa1Rzb+upo
y+ET4mGEqyP+HY1MJ+vRgRlwUa0x6CHK6nqXlzdToUwU9wrtUFU4SEMPYmld71A3
/GcI8t6Sq+9x+W+5jvc8hrBIj600uNzsDRgYb0BG4wup6FgKTDZIDK51n82BNX/X
z9TtmoEw52HxnHc+rLL8M9xDn75emfMF2b7k+JiqJ4U87CsEYsVcbbhL/zLLDI8t
sMB5sAzi7zi57iYkaVmKCTA+CqVu77HYoDqVoLonV9cKNaMDidfRL6oK6//eDIQh
rKpWvi5mPNhRE2aEAXTng2YzOCc5/FjiBkvxqMif/hVwyicOLRgsiGyLbhVrFabY
vOO50SgmZLloSEb88uA8I2iFoD6KZnRJXOdmH3Q8vds6v4zLZV58VvbIv9yUYytY
jfbHOkMK+f5Qypxfykdj1jZHL5qYkdYWQWsoeKawKe5BoLBzaA7KeFeTL53GrXWk
6pdjpY9Rd/SZjb0dRN1kVae59uGWOFwcc2Y55czYVdv/NW/nFa2Zat7bs8srBRfm
6oGfOIRS+qD/7FcuxXq3Colrlrb0Z1Cf/cj/JykZHlGl1WMY9kZVXF7G3vHUqYeN
poRrqretDhZ/rskYGP3AutGHRRceKFpvBb/Gls5+MhmYMAgWVsl4b86nmCOVkduf
1tngsU5cpR9A4nQNDTmLgGBcfcdgixhtA8m2U2vhdEG6JFIgjmLxCyXohOLShpVY
56mfch7552z0K/lTXxVoKHgwtcoTrMnFcioZSKz2MNlC5MSCnzrNmZZ1u/folwdO
+xRCA/d6Nig1krYaMo8Wa5tWvxNlJR1MCQ3EMk1qmp24EBnUsE/WyQJFCnO2S04H
PL0vTbSz+tHKzeBjMbNOK1ExeBcz6G9R/Md3lgfKhAVzrrUeHektuX9BB8IXogId
WiuwlzoKt8iBHxzK6nsj9CO8Ym09+enDHcGrFzm/aDodJ+TwT67b+CPZotL1rRIX
WX2rBcEYyrY9RNjVc89C4YcDHUKsq6dAMoq9qotBPm760ZzCU+8jwycEQVX9ZFKv
urGhC69JbEOta/lT39NxTBzUl2qakHt6gcSgh+5WeXD6D/k32mIwV7ZcpYoJcXlN
4yj9qjqgyIYw+Dab82L6wWxZbSpFFg6rVb4l9y4BgFCEhB96mdYihoLJpqbWK2g5
pnOYqEwHac7Kvby1avaoiyg8PgjilPH1wJICt13PQukBvXWcNZaFl2r6P83XXGA4
rVEnuWjEVYNzXPMQkokUFuvpjhZTC6cuVVdWQdTiudQi06jopL3o/KAfgiy+tDTh
I/WCFo+JOQZpqWGN3JTkToLPfX0bEB5EWAlqTl3eqhtgAW7UvPQsKH3LQOmUMock
EKq5s8NBeP/Ze+bnyD1FWIP5lfSAkFl5//T3LkI5TNzMade9MUqTp4aIl1JxvBKU
bsLGfU/tlJ/EdB9NvWqIm+5gSNXkeDTBaPxB+Y77bgmC7kcnHFTnRC8ruDpmAY0m
WWSpK9JBH/NFONjIlg3NdS6Fpsc5gyBRSwu+W4mjif+r2N2WS+YtEyfQV6833oVE
4QSL27NQgSPTXtjPfRrUT/gSPazOt54q2AdEKRgQ4VxlNMUiSEfvMhclQfLY1l81
axOl4khFc/8MALRBNPvk8aWvl4exZ3iZZo91CEwKdr5DG4dBiAr8nUcd/TdH4ndi
rOczAao9Re7dqGsYRLfzv0QxIVIVEZdHGnxToQsG3hl/y1lLN8VnZQDr/L0Id5+r
H90UdqGAFsgGjkwtO//Hh1zfFCMZktqOpkkbI88MsW00NMmGt5jUpvXp27zdHl6I
psfpm1pg02Pico9XkGAy0lbP8ZK6bPeTYA2luLtZwy/dE4GOuRj8MXTQMbXEyC+t
wUxXjmX7EIkN2qWUDv4DXObUCn8uVCDHyi82LQCFZaJ0nLfftal1lBZ0r5jtUDnn
XYfWtCmHIR8xp3qvKbciHX9JnZcnOX/u+gbPSmCt5MpAWNkkh+eEiOkPCSrHJ5a0
ZeWaiapKfW4TgX4b3CkR3HCDMaetXHWMFwZKH8OmIp/EsP+VOGr9qhzZ1bWahAEc
X9b3tX918QLMhWsvGrJ4bGdWn5pz46oEvYt7tR1TCBJFZ+uz2yMKg3CZ4IXOJ+2H
7hfRrVAGM/0s+k6wSrdTpNwX57b4RMe7pzKtvb1EuNpjfxH02vjdIXEByuc9Uc+U
6PfGiaizwD/QMl/+RjNS9nC9PraGdX8iUhViT253KW8LV3H+lvChT2KPZd56nMfo
/VH/ArGzXoGbBU+nW086aKh/iDpZqD77EbovjSG55qopvgLw1wg1/ZoiWHii39ym
RfJKYzfCBCkNLcFUUh9DUEk2q6qsMXiD0shOatseO7TnvNBVQS+90f7L7SQ2z1QD
FlRBeebp/z6APHbfENPOYc/G2QBdlNJjeMcyNdMFCBe8jwKJ7hr/69Zf6TwqcX9x
YXhmgvtT2KGEFXox2QjYq80eHDdCKIZemjp5w/Q4ogwFgnnM4Tzlzp8W9KzoM3lE
3bz5FATWTbLts+gRe2EXHFfwzDEE0Rl5QGtN5QE5IBXMiI1mzIQfwcY1slzRAN/w
KiRG8aBu0WTw0w8NhKcR2WHaeIoO23RVzpFoF+2qbMZXrQOP9aXmQ1HR4xdtDwsZ
BJN1kvs6GOqELcT4xBf44vvl1dN0cYWhmA7MkeNTAuNt85an1fFr28uIRcnKXcgT
dTzYhDW5aIuYo3Z9fBWXkqrshZQ3HRyXNwiotXXhyunP+UUzuE7znAnYugwn0Rrn
sA+ppY848z13uvoJAcTFiKgXbMTqrAt2pStFjC/KP1bINvfAkae2bVMPhzT1K9xL
dUJ51pk6Gx8+l5qEKkVmfGSsNyPwi9qDdqQHRGdmAOc0rLlW+KPieGHAtti8/3II
cqtF3xK5gliHq1IQgvjY2uhawnz1PuP535/KvIfIixSmZBiHOEnv0Kqv4MHtAyD+
znbnJoaqnFnU+iNkIcJTNTAUvUEsvEBvZSLWbE/g7vWUAeJRQMqCEKZVpdAUi7K1
S2gxkaoOb6HK2ZZEacN4Hx5FA+HEuWFcJu8ItQ0Y1JRXnWC3KwCc/VblwQwlxxY5
HTbyvkFqeQ1hNi4bTOw2zKHwCh6I6egAS4ptbAyDExJ5ISvLyQhCyz3BmeNd4EgQ
eyAdyKKF35ZdqPh1OM9pMN+HFT5nAMIeA9+p2As/uOYyYWxI5ALPHHGhbhbU0h5W
l9fhgiYmHMPDkWG0ObEqcjXf6qe3C9K9wOpWHV9dEklEPAGcYouRvwh99173WIOB
3pRGdUK3JZqR1DzptvfHuXVNNvQWTD5I3VcE/2RTtPdv+144PLRmCZ5Mt0UlbjrZ
7HbI620aTz3vAp72n8TRX0WX4U2HO6kEfk6Zvja0afdtmKp87ox53JLYpP7gjNSv
mEtHhYsoxttv+91Zo577q7I6etH8fw1in9SEBIPUJ7hCO+21/TkQGOGk/0kDaYD1
l8OBO/fXvKLk19CJr7eezXTFjW7Fmea7Qnz8znB0G0iLzMVS8TWsYICF6wAlPMhk
QCLj8THJsCkMHLdv0X80+MXvTRMMc/V2mfInlTXDpWKGB+DxBJZ5JHHBkOAPWqQ5
S7VhKnlUiH744EfdxG2STm+IkoP9htFnJqnZYqBPUbWTeMupb/k1noctNedGWkvR
9VXRb9vaGxlIPRSlPOJSDca8FJT30yJ13XgSOOF+QOMpeWKBVCtCMjXWJYbSor4x
8Wn4YN83mPDdafBEmRSf8vU+I7otTQqDVChWUN7UP69A5I+gIs1ElfrwA8C4qNmt
9xmizqdwXXt8H6jsV5AxUYZ6ZvPaJblrGqCTzjcGhOOaIFfsuTJX5fz1yAGiCuxb
2AhHUx5lK1BLZiQdZgefTC/2DHhxs7YjkNUyOYuaN4kkDMFD8DLrL6QOvT9kiPBR
AybvM7A5nanZbrp+vwFHK6mDZFdyjniH3FtLM88QDaB3i44DDwAt3+DNdWLJ4ZIp
iZZ7uvrIsPUbbPiDM9S+rMwBwt0+jZfLfrYdWbf7JEPSRcjFtZw5/aubVEDh6qBW
ZoW8krBiqZjx6t5uBn5Wb9rg8cUjKnlH6g2HVDw+fxo4ha09lTcQjoB368jm4/fm
WhtVHL/v2F9LMrvNYin0KWi2JGYxXpnGHyX5cyKdbDAcrlp9M9XG9hDSoKVV3Wlj
Sx8IA6g9q2QOR1cEtIyeqqjh5N789uefIVpsWmn3QxyhgcCauG0nKf9f5oR65KwH
BdIczTQSX/Muw6BFeQUF1MXuP/E0Un6u7dpW/+UTo5wCp+g3b7f/4DbEREd3EiwC
FU8DSG9f6EtZbxTiDHhWPQMe+YLuvrmeD+YVam59xL7vcsNHF5Tzzaj9MFksuxhV
5ANFAP6dIDdYrExhsERYWm4mO4wINNT0jKDW0ADzrjNn8rLhg4TaqQYctBcL2ncJ
mqhPFXicmbziIOqvl099dEGf7TqJzztkKLdDqKn0bt8dgA9YxwKeJp/bMt5CV38m
8IrN/GksIJtlQj+9KR670+59/St8Y5Sh9EZThiiEmLtf72ak+m9JuO+nn78sj+mP
QRmd2SY4k0kBhQG5HFulQpTgnyP3SGV/zvy6xza1My0p6ADGhUTYjKIxoW0zFxG0
CjEDYDoy+ERu2dVaV7qmiGisUUb2w5sJPBqh7WwvkmlFo1eJ5E/htUKpSQugZSml
Ajwf+dYzAeARru7gQX1zU+DBNf0UjcZT7ReQ7elMzQqbtlU7Z25xxhKeqAGf8Rb8
ZVuSKEgEdF/68qFkfPP+bVnoPFPCdwKexnswBmZM6+zUGViSBWrqVCpFc/scYZ3i
jU5ioNczmDnD8e9xkNLrCrKdZ71cNksmY2PA2kD9jWk5vWIAvVF56hgkOleb98A/
KOov1FFhNW3+nQgTJ51nMgdB0K3A/D4cmxfe3z55Cdt7x+iQJUlN5b4dnb/A7kKy
ku6W7bBsfeb0reCDgmYyVEKhfjIZW4jnD/7CjZ+eLWkMO7Sk2J6XOk/jz9XIDpqn
wbcnwVGb18M7UYBwKfgF1U3pZE1RV59R9hzJuAt4oxRXxsutTalGK+Sd92jI0Tei
lKyuxaghLhqkZCN4U2Ak0OGYswXodH2GWcxtlTMfSVTg1qlyH/3JnufM6QD2T81N
1P+arXjS1BVK/SWF3dWluiy6USitzIsMT1lfJZ0TKdi4xMdbimOc+w7glVecsx53
+shnql0Bj0QSPpAhrOTz0O/yAZjmUEh1/LIxzUn6AuI5K1IUahY/9guxsgftrZAR
GPfv2kdTwO3rtw8k/2xNufuXeUxZVjcJ6tOmA1a/zh4NVFJ1gUvAhH9PnuyOKl1G
nrKtTfvCY3+NlMoahkOilhaeEmr/8lcoRoLYn8i6vVcF593Tu7rlxrxNoHFZDR60
xP9y61ZPmzvT+HHLMy0PjVoZp2wFxIa356wytEN0XeBJ6sAyBWH/ghbJhCo5kM7r
OM5918bQwd6LZhoWDw8mjfTt9KsFuO2LytnZIZrjrJfB0S0RaL4vDoY+v2O2zoIo
/Q7wVRNnxp6wW6EJDfX8Fqx7ZG1f54jB/ik/gpobqOFpuZs/BD64JrheqpB4l49U
EUn1V6wbgt/4KZ6AFLmYRS+2nMfqKaaz9328eXWz6cdN0pbU0LinWYkNxquG7VNZ
eBnpv8l4yV36xipGCVBoEUthNhZMTbVuIIQdRWco2I/2eLzsKBIlz2xneXwrl5ov
V+tif3p0E2sauNG7Nq81teUhL+9NKs7Fg7vNIwnxvzq6ZFL57uoWdwWKIT6FNnt6
YrsXRaKavwgxHR4EO5EfwD1QCTr0XWBJECiIDmIIyGcnnNqp9hELVw4nYPELWDqx
majuXU4TxtC6xVIFQqN6MZJQTUTHqaw6ahP7RrtSaLS4IqA5F3PG9/dOk8z0pJ2y
avbRXzRzFkxZ+vAQtKOt38TSEG6uLNUKhBECVcr+gQr5ZpjVps6sixexECe7uASE
SGhNr2rDfHJFy3E0gzMlXvU7Y+A69g6PXnBgzbh2QjXSnGLDpNwPrwlWJjQCgVIM
R06IhGYjVWdzJzbjl2MQdQK+ulXgyXrFPRfW3/mdNVpQlcP1m+Tq22IGfAouJowM
2hVIFqg/vSGgnusaAKzA0ef9rInWJ6UGxwD/6kvHM856EEfzmxPOVIU/PQIdjOxg
5hZG5jqk6H0x/2PhMW0TYtwgPhxwww+LmcRTiyUZMhyGDnyNPwzMdAiQf2R4D/+0
lp15m8SkTDaLqTvhyYHzK+GN3vSTRYDfzoR1JfsnFArqKCIX0HqxkSnYXqoPTuHA
5c0yKbl0dOmVAPodODLjzWPuUm0HGNc0LPaInB5nBjvZJHW3hfF9mgHzNVJLqJwD
jdNjtbetQAQ+pRRbWKH5QI3KNzLcDzQFRDqSjJqexjExFODQGuQpBZbpT66FtDrh
G4K6P5WKW29zr0QsRgNy9nid4QlzOi90QWML53igbcwLDzBD7LynVrsMjLyLQpEa
Dkx++c7QOHkuhA58tbyVwHELh0iqe/Sj/jprO2MygZw+/hO2Dj8E+XsMdgeosX0a
xUUEwZ62LPtH48U0X9LDjX/I3jL90IVVEJEBtZzq/KFCLcD1EuVPbfJ/hOJqyx3a
z6jDqotphbUmpWH8bxGjpjKwOB66YQVxjZK3agwQPFxNaiTz4OQimY1X4jdtxJYw
XJgQYi+KJgkszxDNjjpy3ORFRaItBmd1cjAk8QN5yzbJ+qtUi3YUpHWdD1uNerCx
NwcBbhR9AJQlmMda5gIXi5Xb6GHmJUnFTaw79WJeSB0VZ4vyqgX0El+bZ+IvwAgr
1AvCxRgF9GIguZIpw/SupykZDEEX6VqRDWmky/12Q0xhie4JReg0D/Af4mIgqXFc
MWDv1oBeyA7uXzlmlOLiQh+07onrqa63Y28UkllK+x1CvgpTtEWiMyT9guE8iPDf
ZUXmTp8Kxd0bC+gTPRgvJQskIrJ5zdky3kMIYh4JWGo+APAYuPrmjv+xA2a+umVV
4mZkbL1ee5YOKlBS3axOzLMAAt6rVYvfrH0NbtN8v0vuZW4EbrXYmD2eGETpFVBO
/iUr12R3juzfUKn9ATEeWnQVfnFiQWcIgWRSPxrSY+9eTCdlIKuqzfCgQBeiSjfI
VXjpAiErK+ZT6X977rgg/mJPY9568xa89m75A5Zcc8HxTkW2S8lR2f3MaG6Bvzbv
PNxfjjsW8h7wEYgdN2qQX/HHG0q9cyAtQ5yXP0miC2mmX2ImMONz7TAOd5aAXfHI
bX/TCK2ISsDDeHsYVlUeswvIFhMijyT+YKDDtAP48zCFUn/0RE6re623C8xV9wVr
TROpDitwTyNl/8QXwbuHTXWYsvKJEaxwELiR6O8HHZJgJdNhYLfEOmMg7OhyFLsr
1bWccWk8UVr+RIFUaa1c58pJ8hzJjkWwDxmN7c2Hie1AVK4j1qn5ogLRokpGugfB
J8m0yksxPCy3suHmIiNqMVh9s/6Iywmxqihx+sB/p1ZTuS5GxPwNd8vTI+bY9Z+j
lrP640LmYkbmWFWJjG9py6qpLd7e6db362uMVKsfh4OXxjXJR+tQnNdlDtitT5o3
R54rhHovqLO2dftM5nbjf5XdFuYfYkcTKTfeSga3EoJmB8ubagZOvJtAyx0XLgwE
ZSO27oDXIb92MhIqEu2KjyGD9ZHuu38IPINs0PggmN5vx6p3i0JLjylOhwgZGxbW
JHpcdZzPZnneBKVSnNUVfdHnwwD+XnfzK20/0XeEgRHd1QRx4ioJM9tyTaHPwF8R
5IOVH6y0edIIZXEXLgIf+Ibe5A1df/0/k19tAAiCiCX7HG+g1www9zxjzXBu3U5w
4Vg7UGUm7IdyasJi37O/imB2BnJc6Q7A7QHS8xiYMYEDWE3wYZ9FExQ8w7OQJd7p
0uFdLIlEwhm+P5SgiLPUQuBOMIE7wbsHbuJq/Q5B9f7sI69cT5sJOu6fVQImAKlr
LM3iVgDjRCqJhnZwhiqUb6v+UXIOSr83T8eV7lfNF6SWcrQtTmlFlgkVBcT+/giP
lWFwHVkBiZfO99vdpZGAykQbO6xsffuKQuYs4UzhiBqcocOIuiKCUtUhQgP9HrF/
XXMQT+QU7NFcC/vFfWPwdOZk9Ev78QStskh7YgqU0kSRHUwMU4JaUdEvjQSfVXLA
BrqnSxM1DFPrVHG5EoTtfQKu5gxEmubIWpAoaTOgKYrZHlNxKbzGfWfDLgu7qXIY
RQ6kDg4Vibq6L0jAE4AbyjGSDmnn05xjxh92VgKJn5rJ5yO6kYEgJ9hrVHLG7MTj
CLjJcWV67bglaP8NFkBbYkjsuj3F1afmWfQFB635cuH6hHBwvzlgJmfy7M5L7S/0
pQKTaUVva7CRfNploRuWCQ5XUqWMCKIZ//i3JKowCgiW/7EbECXVTB3e0RXxdTJ5
0tSADkuvh+9oR5laHhahAxudZonoY1HaVJtLXHtv6BHxMh0r5nEFPm1xgD2F/2ij
8CqkRa9cs6n8GXHz5VpkMK1lv+5cmtjEDcHgEq30i7X2sdGzXAOIhS1p5HwrtSvO
a+IpSwm4gTzO/cmogerwArUwrK5WJ4bhg/YNx+PpVg74dWPsiZx9S8cstmX21FdK
gNLnquklI+MbePQeLGI1NbWKBs21hmCw4f9BtnZXcUMSODsGLtjtsyJ3xclcTYjY
rE/RvrAY2tBpi08AhPMT0EMPsuIZqPDt6IOX28IdJ1nwvXJItrJ9qeKHpQu02mz5
DvkCkth5YG/x33+LU4zJ3tk8RGFvs11SEkHLbNJdg8lv1XcPp9c5Wz+sJFoePfln
3DOJhpuncMlWejE9ZbeZ+0QUhFQ4vqAbu6kBDvDAmR8LQ1kMWp8mMHkc/onJECWL
EgfF/rg8UC7AFokUPMPLJNDzY+Qn93k6DuxeTYDOVMKUtIeFR3vDLmKpRZNgKw5D
Ff9NN8pH7BM8KiA/avxrOKBK2bElQhHNzNnUolO3Mi3CK0i2CX/0oRNSVUBeURqz
5j+32bU5WXouhA87ws6jCBYoggZN/npONIZNHJmpsuN4WsxhZtzavobo/y+a9Ycb
tDM2oAMSC256ZMqrAV+4is9WPu2gXvvlgBmrAWkITnTAEgwGvgqeu4k8O0b0kpyu
SS2MC5enx5XgWd0r5rT2t5kaLwpP4WvtNl8MVWhG0rTOjkhv1BVez3xALEkgQd7d
FaVLTW7EB7YMPI8KrGl1+G0XhHY8rULQ/1KB0V+2J/NfgnPUqqHg7mbNmlDopqAz
OmzrfVnphYmUH1PaJ+nsQa33M7WFzjDGYIuwwGPQaUibmW5g2ZsX6jJnBXwc0Esu
3fOF9/t9MD35+V+yFFERUFUIdjNZdrES/Al77KkS0LdOUrzIRWJIKfo/8uH1sdw6
9WZh6MnOdM5L1FxWWK2Pwx4G0G5mZB6m8WAi6YP4GLEp+dKlf5BGgIfXPR3Vd1J4
qr7OYOJV/Abw7WKezQb/p8dttzwVQLgdhhuJXGe/LPoII6CaBds18e0tLql/oLzY
MlExai3qng0DjHIrO7P5ulZAoIFcl/GZeN7jxdtnwEe6Wz8q3X5AUUotkcjWsb+w
MPAJtTFGvl8lkAcBtkUwRgvmfIHW/DqXrDZVM5rDAqIkyPCe5/thW8CXDaQUw9IE
IwG53kJQ8uuBpzoEN4/GznFJM0te1I2/6DHk43T+BFn0XiZYT9zvg6LKuW0yWbyg
b2r+zaKLgDMj3Dopl8j+734mXBuVUE10fcw1YZ7PrTBE8zfZO0Ar0K68XysodNVR
rWrqr+gIAvZlWaFzjxrpjBKG+2MNbtapATO/HfOOvjndst/OibF3HQLdDg6EoNSa
tysX6975s2WhKu4sLlcCj4bBQKKK90PJ+IMrGG4FKPk+ugfdzibxtmF9aLtWzdxy
CXFDdTEt3RZPr6v4U50AoHBjElI3s2Rhx6lbxWt6m1tvm7644ZKUzjPkR1AdxptI
St0syVsGnRyq7irGwJz1k5CWBaD39Qqa39ebb/mMPdnRvMEVWQP+PgplsJn5867m
bS1dkv/gAVp0dQLUIAWdBXRnvyWKC4Su+ru7XDHPoVXz5/P8v1ctHjAnaSzEq4Gi
P9nTMUUDJvLX3CI6AX5Ek3EEjQ6i7XxTqS9kjO+FQ+8RctTbINR7AUAC8LBYqZmi
yV/cJHLFq37sCUJAMgvhmpT6uhU4hCnnZUcbLsRrb3sbbOW91Ru4EXQESoNIpx9L
qbVaIeS5FDZ60cE+LwYoRZAlG7EzlZeqmRP8xuL5ZZeoJtB1B4vmfvEsWUpHij2h
qOLYAVtyTG4seBlTV3XnCTVCi5ig2SrElxZoiva/PgslzeOF4TsPNkskzxu5vylb
1PHaX1qgW40VvZfaL3gzS80hMk83DEdUvPsjwBYd0stQwilbqvtKfft/TRNQQFOu
V264229+1LhWLRZHcvQA5LX/5lzhzS3QuCLL7iKB50IR0tPU5ATIM57W77JGcWqm
uMdFg0nN7yqCKcGXmRqeD7+MQuHpLPwysKYd5df91udrBsH1v6GsSioE1kCZykJT
FtRdOLx51TzX6DIduin+NeWIEFOGD8z3uGpVrk874quwLYzzABceUQzIySp4iOhK
gDfqCr9oWTDBpDeya6SW+KsSX+a2xs8KWESVtKmcFCpvjVbKMVX0janpcaaCxPAT
ggJuQghqypyyZSzgQ/hEWzRTiv04lt1u7EO6Qc588Gg/EIDztn9MV/6EuxdtxNg0
PKIREBbrQq5Lkxq8lSD27p8/L7/Cppd/gr2E6+4QZERD8E9UX9f4OvXgS3O+H9wC
tuqs+1Ozw42YNkdlOoyhcaDVQ+qO9/uiqePx2zDn2eWfRbn6xgrzedb7CgCp16uQ
/YzYeNanbrFjekAkCK17dPeGczOjuq9k/GOoVDjQuDgQI0zhBW9kajOiToIgqQSJ
iXf58bKbFPMLJnRF4UsCbATmrOD73v5xRFU+3z8iTE/uYnlvE9o6P+h/1AWG0Sky
cJY5iEyrdA9EYJN2GGm7vLwi6mqfuCVC3KsZaIlXfssQeeqrzRJ22EhpRFL01Oi3
51uw9JjEHHcgY7vagQccMfoVfzlGQP7UJfX0omyru4M7nAcmEwk/Avrl32EWPVDz
bfBfuhzUNCSuK0Z/T8UQWpZm24vSahYJJjROOy0VpEVjA/xncTsqXUoJ8i25Ky86
FMtnT0htjQhMsN+/jVzgxqyf0pqO28WE2hmCE4Dr7O5/+OwMcS+On+t2FxSDrs4v
5zsBsGuq+sESqsz7rFtm1GeT8aK02iy8sf6oKHbdmLKsDeWqqv2M/MnvXdnSD7QM
GKQCmKmOuUUIhPL5x1ONIFIePNc9foOf9IJ4UaDahRcsXX9u/PDVJSaHK1F7g2Pa
ZYsE6/dhUhqC3f/xTMeZOi5F4jBd1JyU8zvEHM0M5OaE67ctQCaXoELqvHX7wYdj
EKJalCvLxD22PrkzlbeClwous9Vxg3YpU3TtcmwxAEGRT0Fj6DEue30Th4BDzW61
/xGcPrn+Zd0uFqmRdw3jrcfcHnqU4PHErwEewI7j+emmuLLeSObUoq+9U5is1gUV
B4eRS+WfXOLmMQr2/8SZ4NLs89OebkgRlmrGFgr5JUbgMgFOcRWhE07BUfN6jXuN
1KIgtYVTBJ8L2QVzwhCoP5HrmS0n+GX1I558rvzY46Bsk6a7jH2Lwf9cmzPWgz/F
UNZLaih8VeUIhifEyrOFc/iZqpf5UdnPIYD2eJV+m9lrjw+xHAfaSM6kHBWug5Vq
bsno/8yKMTQobPQ6AF+OrYK30Mgktppab6ELzVAgOg3Hb5dWC0MLfPVe+5iVxMG7
d/XTXCADW9j+qpQA52AfcRejo4c3TgReRtBvPuQxgXsmJA+yc4DcLtaEkNoNCoKI
BNPwxUUSllgB1LN2XPuCfjv6tsTxpskcEaakRe+uT5af4YzGVXaRGbWLSMwFpMMz
GMtzIOrMY+mb7iOWjk1i6wGhlLUVeMwMDG9LKzwNc/pO7V5JbQb76vaZ2vkjviUa
v8nofPJ8ZFaPbGsJpWPA14akibZlKpiJfivcQg5KfVbLeBiNBjcGIC5LOoKKgjLh
8MfXBqqA6Wt+tokfxZlHXx50gKVM+ee2/KD1ifLIVPYQVptrADuZgto531fX1wKS
PoEwY5YnRPE0+/4ULVCaAr9ltCplEW92giaycEQGX7+zncUlSEquaCZlTbfVYOJJ
ardLHwl0ZUyBY0JLtKkhujp+6WaYbabGxanB13xR8fglls028Nwv6hVudiMohRBS
uJFgg3+VfrUNAriHAh4B0/WvqewSD5B6U2EsxBMXWTlymvIdEpPNDOTYwpAj4XKF
CoSgA7DacEZW0oFrxzENgaBPSaTtm7CCbFAjcMj/y/PR/beqthVaJS8lvz1pcU/l
qHPv0+3MdbPq68mryFs/NW2ov2tV8TYLp+wcTGedHh3pbR07LjvOYHPmG0YRy9RD
ZIaD9GVj4D7gqK7g5ToML297Znx0z/Q1QJjBYLbllJfw0F9jY5gW8VFUmsABmvPg
88tIfMJX0W155ecKcwiVFM5Ft3uJqukrMfe5p0qcqsbe/ort7cdUzkzUD9Y9QHdd
DqbOMFMNuTUFQV6wO6kxdwx1pZ8rPaCCWkCuiwyH7dVpFMjHizE0+P0USePSfOz+
mr07KxEVKubcTJF3nEDKMfY/afovDvrN1s083mqSGXeVeFfwFeBjbIMfhkkHueM3
2wj74uJjhqmOKEx53V4WHfeHfcijhmd6IopZmsuwsO9nPZC166f98HrX58T5M99N
Wf3cyprq8PEFv9xoKMx3gitXCTZxDhIHF6bKbL6abgLyiaoc0HF6q+sdWxra1D5w
lrv6EGuwbWgas3PYZCmW7aYF3nuOYaVyK/AStzea46Q61BX1AJhaVrxgOI45Fsmp
ud2efnCBMZA53kkznVt2fwha/8pJjLqnfxjpeNemq10RNUrHzKpdKysabvkvdtuv
TdXNkYL/WqghTusc6hEiZIRr5xgJyXwV78ZCn5Ftb+cr5mv3QhdyEf3F9Lc5j3WR
w1+kIf/T5fuIoUlPdFQdCNKnRdz7idzyJWnxRwC8QgkzIEI8SL7J00KFtW1WWO8l
Qkk2q8/tPFV1lcV+wkJLEBJJKHaW69eCv0hoNcUKjUkYniL17K70+hqgbtyW69cG
fbGlRzjvLPqd7cWsNBHxf6GVJTIV4Ivc3WpAsBpOZX192ZRBZWwfkRqWMaEtcab9
HthKEwgdQRZl1YVPgWYcT7whcg/qmFHQb7ugchl0mhYG47VHSBveX0/1wsRD4u9x
962y0SdoBvPC442dXltAF9JnOsmwDZxb/JhLJbh1PquigiCd5MIvjrsNDa7H/NOf
/WPATQ4bSVIK0ExtqS/y5gxG8fhBIkbUAbvvTjMfzc7uoNLhhzQRuDnK3GpnI0Gz
HRr7IiwIdf8bDa9VbNuptZvZBt/IiOR6dPLZOLHL8P7utTIZwYEhCcrft7ePw5Q/
bbJJ036FNnW7chWJkRkS81ndAkjd0aRDXYcKSlDJZtEmUs6XXg43c70DAa3oqa/8
eOx3OnkcSDu0AFGY3oCzDfIxnIPSR0EHkWZaCdiAmOOs0OKbIqXKDlNTOOs6gNLa
mSP3Z2FI5vBXWMyPU/yZ5/L6eKeOs8pkSVwv13nLoUN/d2dIvRFbrSyVE0uApq2Y
Z44b28LumnvIrnES8II7g5IA8gSpek6ywfyMwa+vJ6Vgs0ENg3ZbhV5QJcl7Y9bp
xuh4OT3wl1dPIBQZNkzxx4HB89Ylbyp5idSJwAYojUdxGVxJQ9Ksg6UqiL8+I0gs
f043ToBo0pth1077nSQgdBWbPHe1dB7E7tecnAYSktdCrzJYTxBRRKUI6LxFjAvA
OztHK5IUpgUJcOd+iOBUzwqqv4XvXdNrn+LQmORcBr0sQpyh0z04H3XlCk1ce277
sB4/8RP7WdY6hpNRdZ7AVnDu96bVFtAdXMhz4tDY2alg8g8svzO2mb7GjeMP7sUG
OnEhmfCUchhMDKmQisjOTvkQskq8Mti3V4IRCGQC165xXy6s50aUqNeW84oK88v1
ok0WHyjMF/Aq9WMTQan/LsByQlcmSq/7ZO+trjZUq/kJpXmescmsmDHf0felf57q
4dPP5HLZjC6z4yd0KI+a6/whQmCoxuLJQIWcOrYYGI0XW4UFlJuLIceCtcdnHbYU
cUNjOKGK08GuqB9YYFcfZOL18omEOdJqhJv/2IaFkP+8sRuMUFLFs91zbhu7oLN4
HptQVkJmUwpEhrBldReABPocDDCLQEWigXY6ZQZMEvCWZoI6ODGNBHb6izkFhrrl
FnTAp+IrmjBWNIeVqVeEl6tU4p/TsbyBaJyTOVRRsS+BDEmMTs0ptpSPU2DvfvJ4
mtDxlv/z8hG10oy83aqgH59mwcl+WqYAjg6t1KLn95C3nDa2lXsVX6GCfSjKu24f
YKb3VJN5Qmnu/Iplo126snF3uqFv5kf31ZlRLXeiStg2kCcsnJl4vN0I+owo8TFL
zHKZLY/DPP7JCZsAnPmZsnXnoVhjfKdIiqAHhlWX7RUOyGC6bqoUIR6b3c3go0/C
4/L4mQNKGnmcehutjMR5/ajE37E3n9zWAXT3iDYgk01oYq3EnHtM5RNTsg0ogKLD
ng6aaCDDW2vgL5/AgCuw152CKOMpLAgyt10FIX8+mZFXjI1icayw9LctkXvtbLmO
T1Zwb+vFO4L4771/DQjOUA+oB7eSqf/yPCLt7jVxg2G0BnzyG4mfFrNpVnxHcKh9
LF2CNkBLLGtZZPUWW21+NvMuC8lbzX9Ya4eo7HqQnysdWJuRTCTY483GnD8pDwRQ
7oLadRrXpNgxOMdBviL6lOTC5Z+ri0ep3GBFi/eLrHIo2HG+X3RcKRmHnlSQzjtr
sn4tKWcgyUtNPz2xnN4XqqVoqWGJYgqD6+1Ioepvz97RqLu845+zLQbhBIFRQ8RI
MZ5C/k6+iqSDhGhs7w24OhstbNYKLOWHeQeV7t7lfPgvMGvcVzsCiOnk/pZj1t6J
RakWcNje/mRAOFoBDxPhu/QHLZr18eWdqB4ZTMKfTwVvgqykO7yNqSI3kIx4K/UM
S1L5cNo1NHpYr0VZqwk9Zr4jTgHsruCfVE7ZlA0WlIJgFl/MkUUGRVa1tFWn6Bpv
xLqOPJIYp1hwGrQayQqWpVrFyZ3wu5XJcNDgoawcEd6OfqvsPStfvN15fdtQXPED
wCeHbX/GS6u7m3dQhaAlXGXsTKglE5jIou22KBNLQBUgfhlz0+F/A1/zcydXvl73
k+cxBgCx5Du2PFoP29vrmN0yDUUNjUS3szIz42cw5zWg9mCgn9NrgNOPmhGcUDlu
Fz2ZOtJ6AK5SpGJqRNlGONDQ8eyrHTFXAYM4GUXhRxYjwOON0W7VHca9inT0K19x
TDcnyzJbtYRfdRmcvkSyswrDFFQV7vDL7f5KhhkhpwMPP+Nq6umTP9/jwFrwzafv
PEB/f1WhJAZD/sRaKxhxAEi+toZOQ9xJbUAibbb+DwcKWSbJULEh9dz4t8SwQT5g
L3lYWTY28pKaAIRlIiY8M+klTa2i3m7HWCd6opFSMs4Eer3YWJmTW2g0FbcLFgYP
9RdAdsyZRv/O9f39GVTxIaBD+zgenX6BsD4C7HTn7tCkN9pMEi/qy3n7m/jr6uPz
xteCNPaAaX5Zfx2x9cIne/76y/xtgs8sbtrtOB+eVbKxc031/io/CLaJ7ERnhWv8
+nJ9RGVMmje6+10p/L+B1Pypprgs2df5nADSP+g+DcLFT9HO0SE6q8J1p8mOu7t5
lRcV0F3y3PGgsbzefmHYfvJdr0LZ8gE7Kc/ssVCXdEMwH75HHfq8gpxO82bx+Yew
jP4k/E+woIYnESZjlhrCNiNwmN/uA514MPdKWl3zW05LbuByDPtELTvw22LuZ6fy
6LG6trnfp4sQMHiF6Gj9jOcToc5WLZfhvFWy9h7OuU0dmHO2n5pFh2x7ltDzKXAE
w3GSCh18tuzaRWbTtpieM2IFPFHV3DkdH5RJOAze7g+uBpwaTsZC6qalCZPMMyXb
ToDM0I/lFXhEEkoofu64OxMxkyF4jSR5y3UlV7lMFrrCDScL0/FHwmCEgQ9Lmpyg
JFdDJHTcVIPPu0oVmB4URqBTMzm9oGcl5lBHk+XmI2GQLlT4Y62QvUYmJiPYm+jh
PmznJjGZboef6F+bXDjgh57QWMB2W1x6mtfSCQVZNPEVHtwnN1KysWWHK6qSSyLY
5zg4OK56ys53QEuwSinkeaA0rSCTXemEy4XwWCKG7aGX5wWLZxqLOjacarx/poX3
4sI36mHJie5GxA5d8n2FRJzRYmgZ9ycY9ex6Pwjr+4m9Fjp697ORuJ+jZAiyUYWK
cANCYHQtd7ZqYwDE4cFQhE2JKAuyqGk/YjtrbY/PCbhKEmRU5GsJyJ+V2HN73ILm
7E2T0AR2g/zyDq/OlAmpvQprnyndSfsosIB3a60RbH7c0mQexHH4d0ezuCLUkoPu
lA1tuopXHM1Zdh2lKhJXOLOLajCbCy0bFo3mSEdTbCc8IXOl+6EH9XUy8dbJcL4P
nUHMkGFUCzx+mWJRzQApDbt4iJ1mx/a/LFEM4oUHhF68d7N9smWx9z0rVNxKpMO8
J49R2yAjVEeMv4m1cYZ4mdv6NXYwBnfkqVr0MWEAgLBDvW6wBrv/anXEF0oSEpxQ
zbuTRG03m0GuGCatmzKRpQQo1GnCpQ4qgmnXqlDRblgW3XOMqUbAswFhUP5ypoie
1GUF77XLu2JvlMhPm7nMyp5eSCSXMvslKyjSBHit8urKjinlO5FNtTGadRMSX9pV
hQJ2fj8Xaq4R2/D4095QBNiE1WZLdjYDDerL+7h0BKjBzdZwZKJKlVFiWVcv9WkW
Mqqlyg1fje6DqhxU6WDyP9bqf6/YFELR3tYeCviCgiKlnHRWaoOzWN6nPDhiMezP
jxj/O6uTyb4OEV3z8y5zpOVmRsCRarLZd+qpL/87H5P5pG9BSeKVBud4G6WD8+yW
urwERpiAGHJbEpdy58n3fqashXhMmLR1zQ4lsjARGopW637LYoIog0LPQ6DBDlma
FFFC6eT7MP2SAxZOPctOklcpB17XVGBh88yc17oTZFQBBejSOXv2mOouahKpgKQi
+x8C4sGKMLCIoV0U+a2MfTjl09uCKSbrewGbrGoKRBvVvLnMzDpxn06z3m59iBFG
iVctUYD/R1v4s/VLRAqt7HXMXb5Fr+fJc3YWhBdLSgQdJIW1tT6oOrBaP47+UFO4
T7rTLGapZlchpNrFIu4CviRUQm4Awaa1PbYLJWoQBeHyXG745JCCQeQd0B7x/iqT
91zsICs2OcHAKMyIVoWoV4T1qmVjlButWaAtw8IuMYD68k2zmuQ+v8bOWX7GZ5Kv
0RLhVYJgo2BXPbOvonyvSrq0pg55wBFdoHjplNxMKSzP+hluxC7T9kY4U8PlB7D6
Df0zVhqXWx+1qD2WN2hk6XvmDwkC+3fSe7oyeuIh4NsHkEi0eT4RC912tsPychAy
lC0nrkkRlKVWCb5mGHSc6MgCV6QiOn+gDcTYk54YSUoVLIvJsrndSLTD7y3qg6ks
La+G3PNyYGKN03ypvWbHsiNOGakfarP6EXh42iv8a9odmlPdzPTe+xAznM9EVIOI
2vswI69Hx5V1a9mP5UBJXajfIteDqxweF1+FXil6VG8BtjEdbLxFW+d0kQ7t3sch
YR+keKKkJUAEsAwbLD/60Ku1k4suonI9WfJPhnN+3YLXAFS6eJ5gCElHaUQDcBbc
mEGlDovG7CBgbb/OuuWqkJ1l7xF5D2sgASPOYzJiJ2kZYAbKEtBd9fuSW6mHJT99
MOVS23ZAgE8cpqY038fMKiubojj4NBe2go0+F3MZhxJQIgfQZOwojVXpCU5x16bG
niEMmYPulgEPdKBWJ8WAvm/2prRm+HlvpYhBTdHJQZ0MIKAGCyYhAXECBUMMRL/U
Dqtfue6XYBxx/s6sh27M1Cg+mbC+bqPcQmlzaDF1jtnNH2o2sR2aQsEpB/ykCE9M
W6PzCb4aaUT3jZ0W/76BMvvqR5Hv++kGzDIC7Aeff9gEPfSKV4aXYAe5natCSpYh
OT2zSrcN3LZaWUhf++UzjYstZnUE1PXBp2SUCwV38YQGl9804td1yhx5lNaLWYDW
L9cwzyRvVioAOpzi8DSRMGqz5o8/PxlM83n7VK5xYPgU4Uk+BNmwWQ2BxFy9nf/P
JIxgtELBsLFal6DLd+ZqIg48c5s48dQqjd0OySTwjvrFmrPuJvUNn/J7v1XfIbeQ
p1aAwynLJM1WUEoH/tflE9lnzmiUesOBVuzcuJYca8bnosUqBgcNgysqHbiI0blM
cnlpw69xECGp6B4R+hRb6CNq+RXsbxVmU5Vg7z/CZf6uj8j2cgmprfLfyp0ndc4G
c/se4E2QMz62yVfobHvGVEO0W8iQ1lPkQmDk0XhTuM5H/1TfiAKfVNvrnx293fAo
IdhVYnyS2kv6qMK4FXYP47lui/M3pjfAoSzuAUcoEi+HHPLlDSoR2NsB5k4ss+7v
ld4bJ9yftPX3oHraENUdY/UuZqL9crxmw6Ac9giUoEHULcSNWx4iT7pUFs+jrudl
FD3d83cvShuImMZcrqix6RKxN75xVRrgyMXqDkQCufP5FDcDAsOaml4oLDaSTYdj
KoT9O4N2ErfiFg9J9G2acta3o3GHJDpaZ0lzHH7hxAN7r4fSRKlInXkIATLPq4dv
3jOQsi5IrM1QyezpB8hh6hoV3C104EU76kKMQWT9azTm1TdQUCozx34rVMgDa4+7
SocSxHMg5tn9eWHvUfz2/HaSz/lTOnwTfmXuQqs+v6M6C/3cKk6aG9V2/+UrOKQa
GIXff3YLMqtOlT8dbsPQiMBmdtczvNjcZIqyh/snczH+1F9mIiQxNCeTL0VPTfXG
oDLZ416D6N2zVw4US3KMObcOZ3m4ROys5vf4P2xsm+OoNkD7yBCaQv00DAZNbGo0
AEV0IifnhvqfWS4SsKfxiGu+dXJum2YszsjKaOxH/DGDkzp5svFXlTK2gn1XGvJA
KXqs0/PYjw3sB3avwT8ME4O7T/EweIwfDJfz3mpfNBeuFWVNHS3hL3GhB1RBbGPi
dCdlrEhGNwPOA2HjbTyh6VuK+fFTNUNupkMa4xjw0DC6+usjqiMSYFMYFE59lKMx
3wqohGY2GeoohBP6oPioHOaCsNHcWhUssaF6LBuQEMT9Oqw1lVC4LqvsI8oPJ6zT
fovW9yuol3ejpeOUO7o2/ZtlHFFQaR6fEWL//vJF/GTFjcN1o0uicrfOGX8sdwcg
4DQpxLeXkoZ55QDfIM/pXM4F3r5PRnhJbOWAqgcmjbrBerr5EvKOCtyKKDbkfvSL
xHoibYB25pkrPr/2TY99VV9gtdiGLrflLtDN2m70NdrVRmqa0dHXxIef8mc2kmbR
UVIbzWgUaeBwrykUEB6f09cufC+zCP4UmeTupVHo+f4/yh4UUno2hCCAfszEMN6W
/N+yOLGE4hul0Aa2m7xT10UJbTe9UtU8yO8HqaOWtZtMcZkMOniNjAW9zOPAd+PR
oKMkQPTeJU0IiyHb0cv7eFIdRnrAR1ctkt3EinmzchQDUrkzPtVGCkySjp3lS5a1
oite/tf7fIvgSESpo7DFzLKfFZaYjWQmJGvXjDi9O3Pp6ThQjcAGJ/TdAbesCw82
SrRBa4aXydqhPkcYoQItNVVUbQdLsIJid6D1m6xmnXAvSduEueZHiTfd+ZSNB5IW
rsusE5ohys4wEPbotfCPshMI1b8WnYfmx+fOiTwcd0Y0B/49LnCGdAG6/fm99OGF
6HXwZFzH4dOnxO7sg3iODWs72yGYf+htZd6/zBp4FJpyMb+y2mE/clcbOxSRQkni
7MB0BXonn1n4YI4/R/Z4YZoRcWt8TIT4EOfHi9tRTdfENwM4EDHhzNSH/dygQnTT
41+XHEqZ3gLSzpac1j1ZT6rsj34R1JvYUeHbdAB7sSpWjqtFNGYxl0q6pHKCnl/x
XkZ5sehHb29A0jUhj/g+HEh3rxyyqZ1BOC7if5amlCexH91PJNss/RnQEZnqjpSd
opX5lEs00iELmzBfDR40idrCiJrF/i1OBG+ZWZ4Q7pVOFDY5MREruBfRM8A02So9
sy/QfaLo6espZaSqBOnMxIjaKwIWaJokcaehGFvJVOeR/+586vohLk/0m/znPXUq
YxUxEEFaSOky/ax2+2RoNKbsqVFWzXhXdFtS1CGulEWIoVjZFmSq6Kogw6uSaJc4
KVAmKL8Jn3tq/AEtjjRIyNLwp3zDPWKq01CeABk+0/gqRO3xSE1ADqpkGdkxg1qf
55sPKY/7DF8AWqq3krYJD8SwNYYd+1jlwCuRCQ1fO9gy3zVNTdcNK+HOWOO+29y+
T1/kKXpFW8cZC/HFgR+MXggs2tXPH9PXpv2OBhXgdlrJVdRv+a+Obo2QUB6DWCxw
iV+mncPzA42Xn1A/pxkd3gmgJmF1/fQzZGY3s39V1/KUjeWcQVeu/9cihNnI4hm3
v0IY1sIGg6Tq5LBgBDdkVSDKphEjJIOU4alf5cT5L6M7ce7nHibZO49CJVnqMfKK
xadmnOJfg6Vb6vCYSWWW9eR9NNIPS4LvKnW8zPAgURre3cA2EI3yJ7njeyrD28Dg
QvpEAz00l/z2B+NLz1rFrb8ds84vOyE6rV8gBWULBSWruwE0YbRM3Wi338aUAWtf
OZ6O60OXFoF8klCAUyj40wuOa/eLISezjXVGy+K1dOh7ZWYbJWgWKLGZ4rsxK814
YNMaV2X9jv9H39L6Q7ZIc2GL8lqFmf+IAoYMnB38FUHAZGXSqSnXpq51U2k3arO7
RLdf7Qa88TqKt8Qu8MgY29ClJ2CYbNaYezeDMn3JJ9DoVFenqGF2YOvmAr3SBN4d
/FIpQl11i3YViNU5m+1Q6WUh76T6AhrEjtTqW3BpGHCFzwXHkJrJXr7W9bR5NUN+
LCerlIO4jtR+dBb88pEyp98Lm3PcFmWFPWdgdb2nWFcUjhMIiJ9I72A4LGepRtCm
fnJW2OTybX04iwOBMt5RiSuhV2mHUngS6ZS2IrzsnxtTvk/LgG2nf5YkTvB15M5u
hxEfAO8QDM/3VDMhFprZ2T5EgyYPvop3TyTYs03I1G0V52xbtbh8q0FLe5F0yPdM
Tc5ehSIX/dsRa1mw+eu+t1WD+umLGij+haxUz15UfqYWyG3PgPWxHUOTYaM1idhT
2JtW1w53h4fkKl2RFyhp9ry/nCWROFzoX4QU4+vWsX4n9vvooS5XzTd3/xZddd3r
BCni93s1vKKrj7qgmcaYknUG6dTHcY46tUsw/fiyxuBpu/hvZznUgj8FNnSYKwDc
ckX7gralqSNMdA7EajZQisyFq3N1Z8X2rMbHUvWRznMqpoaidL0ENNt+FWZ84t9O
cxLUYBaJWjn93SqdCbZZ+xqPHxFTINke28dEdyP1EySM+0m/vSaitC9pVyLuTuVL
MEdi5316sTp8RvqHtLIk9n0+oA41AkJdTy/11aQnCnov1/jQ4KgBfgrJ7Ei4o7GR
zDp3cS//aTevk1CMDaLI3Fv/0qVQpkq3OiUon8ZwcJd3CbEBBP9w2ujntwV74DmI
glSH2ZhQyIJ0KFt5itJ0ZKjXWe49i1Qt/qT4nBRLCUp+EZdXOeFcscrKKod1+NTG
KErdprA9bPN3xFHs63H1TEDsWl9eNyq8h4lakKm2gWRJkhg2tbnK81+oo8NAAjPK
2BwBvoMCPI4ov9WdUJ0SprQU2ggBTBYfRfW//aRWqTi5LNvYwf6xb7gTkmRyO3/E
6MtCwUlPa5Clr3qF9Dc7WCtDNQMrvwpMJEO3aobtCdkGKBMvKT2ye2juERfSEkBw
JobAmKJyh71BY0HDomhTYow+Wp0TlrNzoW2co5mxFNxvKcPPZW7XgimQ592uf2Vm
nsbN0C2zCSsC/Uk1GBO9y3jWF789P/1SvR05kDOeLUJ7OBLXkkmsVAeMt/dXZpjf
WoBsYhsYuZfunF7Nkj2jjZRJK4gTgjvcVJs7GUVzS0IHt7sOIdRAdKcDB7c9obPx
A+foLc84rgZqOV8aEXwTpltpcsywKBk5bHr44flNcxQldHH3vNfKn6aiKg3X6zPL
zIQQQ8KQLC+kObcGSBks6xAYveFvqo+fJkxOueH3LWsFOfLMmWbZMp7mju+oMNac
1rFpEvr39lMD4LNm4XA+RHr7FbZA2565TFLPU2H9GUUACHk0DMUQzArYc6kLdXhM
2cbSf9Q1aGo5caN8GHBFkUxFY8/7Pw/JVwBeSF6+8jFJc5uVrnNMGw8JxB0ZP8mN
3d0hsK3H4lJwTjccYRkxO+O1iieU4GlgYxKXEgBmkk6lKNuWg2Ziu/0yOf2OgJ8C
W/Qoiwey3FA8XWataJfszPEpCbSCHqJA/RYy8FRkv1hOg41vICk854MO45Bj8W8n
+NVa0cQSWETSsaLst6blGoQIPwIIkePe7LhlZFDfkyvVN1wyzdgVkIvB+h7AU8LD
/rPOnS6JEztmNH/6w0n9jyJ9o+dsHcFUNwEFThswCulzw4+6fcOioSRw/vv1cEAJ
DCgaspXRwYG/HBK58BMRWsztwiq9Kg+Z/9VuN5DRXhj5CpRbAnaG1kFTM5lGyZ3O
GSJSC4Slr0glHJFPv06ecjbh1kUVPpqGDz2ZzvAgNVIpsTJz2t/XnAVYFixZAni7
MVPxigSz/b7Q7ctmKOErifoW7bepLrRIn3VjHxNnESYOB4sId+s6ZJGgdXLfOtqH
alRJ1zN1NnUXOIzGWVOoO9w9mLaJW9dIjneZbbweM+Gd30F+v4bkCBJrCRScqwyM
f1KZf2smzNOXvv4gVaUFyCs+32a2H7O6nwJi7SfIymYK3m6v2o2jBl6TvhzbKbFL
4mYbXLhjoG35zkdaEpiakharC6Vv275fx/9CZaoDBcFuusB5Y6D3B6NKT+Y15byL
qRK73vApNuq+RssqhbW0nmU4Oqlph929hd7CHQZZOhczXj9Mr0bKIjvigW0Qmgcy
LElxTP9yCpB/3Z+RgQmVXK6/ekLWSZyeWAhd8HlhL5a4ctztw9WI9MVCbrokWG8L
pjjwcJQMtwId2wiLp4hjQGXfl180wESxQzVu/fTAJ1GfB4z0XWNuaYAen59Oc6sN
8h9rA0Ivvo0WNJcyxws0WMimzuxmMXroE5fR8zj9FdmJLWFvFIpfAOWqW45dI5vR
dmDIlBTkj51J+GtdCXp72aTq3ZXjU5dRptlSwjE7OFFC2Q6o9kwzlKAN7jqHp9kc
8weKSaKFW+xM2Zu1pjQUVLZp9zAXQR5sRULhNKqK6JkA8zJj3awOQE9YBzbFUkEq
UkjGkH16spL1kwk/2V2D8G2KM8eMUpRigRckXMBZR9atvKqIZNPb478xjt5ph1Np
TUm9ucWQPzaCZ6M/gre4AF6higE6k2CKK2P72SOvDOP5AHyj7LvqnAfl4K+LoCVQ
L29cQsTd/qWKrUkG0nMvMIcN8Ev/hZXqqH5qrZPAR/KP/drHZfeWRdjZla/A4MPy
NweUcOpb5U0ZDczIDfamSK7H1w0YNGD9csrbySfoThflvhOo26POaEcyuQYrKHRV
YX959d+nM2rJnkafYxhp8hHqOXOQJFs70tPDpdExpO7Vhat5+ACycYacplRhFG1g
ei9wFMfydsW6wqEERlxVxYb03ft5pkGdmlVghlSiLt3MoYqmXCUVL35fJTn1Gmre
+E1HKLUC0KpFMfXoer8mw2wCeyDT+FyGYOuhEIq78tT4qg9aGRVU8EdTMGwwWplY
Lp767Dd4p7hGdrxDUY/9tVvZq5R1tZhJn3wqAR4K75h8N8rV84HX+FKxdUE+vHEF
j1TLdKcwm4/+Iz2hVixocW5b5omQj468hpz6/LyB3/av9zjGFSyvlDS9LG/3wS4+
vvoGB6c33jhQchI5CVFl3GepILcblFkJkf27d089636dsZeSgexijCxQ7pQ2sotI
AnCf0cRV/AEQOdi8VJ1boRzU8Xo/5yfrWYxWEfqNB3UzoGPfjkM54OhUif7y79kr
aAqQTBukRBqiI6lmYiTAAmJAWTCXRytufD0Q4nM0HDuQV3Zl8rcZ19oqQ/8Elhro
GzQeEPgn/BzZS1NJ5iCRIRfire+RY+CaIbPIwT/wKPJIvoQL6UrAK4gis+S5eDgu
Ha456vA7C7a8TLJS7e1tWu+ckLoabu+6/O+wV1cF3GHcxqrDXzjVsTcWxqGJgTu8
ZhqG5xWkfrXWDexEunMBlDWKQLkJ1RpxeurzJb3DqK5zH+QbqJVcJShg7PO7fFui
j6NxoI9J4tPZIMw8v6qtv54IuP3McDJdrqvlYHGyFddfHuOn1u0LdhP/4EQpXAr7
I0wc2fogM9MOK1wxAaGTtqEG7c/uqHOEAph2hfOYiUyp1p/Bt+TCCMRhBCHJhKnv
/POfFs0DlHgy3GoXCM9TKOP9SkJb+Cn46VsbbE2Z6SgAnx/utCcAlm38bIwUYGNZ
7otgGoUdN1VXPBXsVRoFMJ4srPMVL18Qj3WwuDXJtYbRzlCzBPevVeVzDuDPl3pR
Ga2NDACmz+s5VbABkS13kyX7y9+Qpcf/fmbAzoCaqpIDLKvenl2E4FmNAlLSU7O/
Ddvvw7lPoWok/8C2zVNttlcII3win/1DrrWQfXQqVylkGbgvQpxv8L1rvyFQ22Xc
cAzzMPwmE85t+2UCMEbr2FJCd7RQly+fbD3xmRoaVzih5xN1St3aN4YzekXiqe77
YYYWPBuRQKk2CG2UnYLcJpvSUhOY6c5I/cMedY1ZMOtSimR2y+CKKz24O4hNdh2M
5j0GXBXjoP7rBRqUVqFAGugY8JSYdSJkpaY55JQcZ+qcIJtqdR087tl1OV1VdShS
jF18nlfEmuoha225Nc91WFLIlE7ttmzPWmrq+h5t/bagX/xmEN1f6WRmUglhkpls
18rVK7ObPrEy2kOYkLf2lH80ZJta0bkkZcMSHsXvQiEXKZDu6nWltI4b6vTVkebk
DHYtGkdWriObIPji0oi6Wwwqj0arGRvLXSRgFRkm8lSLAysmJyJPz/yvGCGA13Lt
cxDHXfM56Rcw5hGKxeu4VZX0DZt2b5lg9hY+MU4U88NPhOmqbZ1gBFpT/2zn74qG
S/kyenlWVrUkBJkYj9UOqmnpHvE1lfuXAxoEZKgpVZKJj+6yMibQM/gk+ySwVX5K
ENyn63rmtNWXSR2C7R8L54W+zOBGezRdmn4Rr9vux9hLg2hbTVPgOpc7IMwaUtbE
7bQ2se2RHB2TrjWWs0fntod6qU4dorpMim7jOWCCaGDVpjp0TudkIB4j14CjEV5x
c1X+dhJNaC+kkrcGn5mY6neZQQPh8yqfw0rPS/JuUwfvdOuppqS8WXeHZfUZMQiC
hTOJi+43oAujkCwXE8yajhzOgU/7L82MhP1xDMOm52zqDO+BJZAcz3Sgn9v/PBUt
AaeunyycHlXvTzjZgDftgzwB2cStYre5LnT8c6MauEi55PPTLyFmZgu1gkFmZlUr
mA7B3NszTfzPLmDh61ym0X2QJK13j/CKpyk4Z7ducETxOFfxuXdgBBwLICfgoeZZ
WqtwV1qnkzj/wTjFF4167KG4lsa2xzQG9sZRRqUkXKiZ2MDH28D1DWKOBcDkLEDL
6rgtmVsF2vDn0U8FilzYqooMyfHz9UJaS30hZCope9mZrTnFR6aWyJ+jZhef5mOy
AtxBPTGBxRodR7N6x1CZg55iU74xRUA5KQZZ8y13SxB6BpcGzmx4mtql+vj5wsQP
7FciS5z9i9gn/1jAVx6srAU3YYx/kfUcuKZXBnWoJPBaKBFKbElfbwcfxLdeB5Rz
s/Jr4tWWZz7FIEtyKSSbiEmRedcYVnrU1FgYCHB6Ud6LMuj2s/TpgQiawI9kqhjE
j9FKulX5/rz1UCeN3ShLB0eHcVRNK2jOMriKk6clvIdMMLy0qMytuyZlLba156y1
820nyITipZ/UFwchpmU8vBlwEkO3W4PoQSXjyxO0+BQ=
`pragma protect end_protected
