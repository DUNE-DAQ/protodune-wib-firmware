// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B0AxSFEBD5ZXOVqsrctzPYTXzEs6XePYx8EnTbuYCSlK3OohyzPN2+BwLtq/QDVn
3FrfIeUS1aLvM6Hbx1FzXMrNMwfhlmG8NPQ9fp7i5tZdlDhN1r4f2hNqJIGCK/FC
UhfxVpBlEtpIPClM44S5v2mrhioHq3/rMle1NKiVBpw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32976)
BMM8tsFsdTFvSmTFHDjzmB/GzHpLxbN2na+EqobP+oRTFT/DSEXtcZDQnxsnKhHS
ZsO3gMw0kOwOx7wOev/bDJxQ9EvQzK40No2KWzVzzgQ/F3m7BkeHFiUGgb+i2+wR
1FKhMErO8Q8zYv5S3wLzqrBIYFEyizVd7lgokbXe5nSRTJT2I7v020/gQpVwe7kS
vj7K7FoXJ0m6t6+edJIiY3BIiVMgwpToEVAB49d/kvJCnKKFPB1QGPIYJCcuiWdu
/9KXqlFsXTpbs2vgEhrlKibLu/1hQAvRMvQfx4eoefPlh1V9agZns6/liSBKFzur
Gl+6pK8pUscywgk7fa5vKxQYuFE/W0WxNMb5Cpj2UiWUC9wpYVUJBfvpoFnUes6V
SYBySXdXrMieJbmuww6Z0AZG2w+bG4IUTrinx+p8LBb7qx15ZkXFliSq++QEEtow
Ov630BVPLD8HV/KQy6i3/01euLtYAXY4rpPpLs1ky79jSuAE5oV2femvnYEBi7Hq
cMz34PjMxf8rxkQuilryUDSWkzyWzXvwaTl8AsoRcxeD7Ix/fNFbzB6V9966gZ6R
adgXL5jTJcjIkSO1kzw2eUB13OJEas4Yag24XclxtTUSDB1whG+FfKmurzNF5H0+
yb97aZHAuZiGZmScbstndyel+xgPgGRKjh9pEZAKTg6SP3+q7PGzF3wQBQ7nyI3d
HDItfP/l3iV2kdAg0slH2afeySZFQ+bTBWgbXASP65l9b/590cIEbGdqsM9BLjQI
lw1qfrjGxcSLnGdCpthV4lHTPf1mlS7qcL2ctmaGj+VgO9p2YIV0+ZRsgfcveJ66
hwMs9dkG1wmGSnNelMRTY/QsOwpis3ix7R3qTic6/2JTy5+cA37AMRsgBubVDzZ3
dpjKr9LKIvk89PrrPpM5x6hwNQCa6IJci+F386kcf2rQpsMQp8EgFKcq1zyr+MYr
z8tcQXfg4aeTyBbCa5HcEIrjkfJMUeokddG9pbfCNPGtMBc2P8TbF2LRhb/Jqunw
1A0lQs6Vg8TNKqbcLCb0EG0qWjiW15IZXXgeTFGI+61tfanaUl6KKzL5IzIuTrta
aXGP+TagCgsX9oTIqrZUeLsE+YerUazo9jGeLtS9SVmWDKyClZgRVQPgo+IcxsJr
KEI0Q8KLkTObM3sGnOic1T4MW7jlhWjH6BYEErQgXc4ic58CUBf4ZpS6TVHRMMy2
tbHMwKRMuXb44CsAU0uO/niHQy1eFWXcs1pE2+7EdsQk5QQjL5KwYIS8MrAa71it
W5zmz50mRzBPgufvEdW9VrEzdtgWQkgdEh5RpqEV9FHyCgexeorJKuvQtYmx/aXG
pBBSWSbK05VPiMIgwoSCeKaxcmzzv7KJmZhRcgHzUASt9V2Ph1rSw6AE4ACRGZg4
C/hM1NnuXmXyqItwBjYXa7n1mEO6vpBdfvhSzymMXpsppb1IXZRAUlqWSdAlMDWF
rQkbPoul9GeLiGoCN85dgVlkxkVeeQ/kBtpQuyjOYFv2Yy3HP9Izxzac2itaYIV5
22xXV0XOh4vHgyNM73+pnBfjKw3MEcTBhfd025jraAUU2G2EKoPIrLCbKb2zwX74
htRMOLV3fPKraxDJ32dzwCs4KtIKviQOYuUtHcd6sejf1FqJbE0Ftr78ko67lyHP
gz+eolF0jMu07U53aFAgoVgBBQhMB2m+CaDKteraeFYxK5QmuE6ewv9Ozx55XD9p
Rdx6DshizPQMWDMBMYHhFW9KQNDzq0zDGS8yQcCwU+6L/R0w52k6J/znCuME5AgA
gY8saNoj3OBb3XPQpU3GvRrCLfkJxt6kIe5zU8FiVo8PEgOTNZG08q8RwosJi+W9
2kLBfdlOdtZUALFY+zLXa3zozqTYZwXcrl8bJgTL9M52xeEj6zV9d5dRqQFfMwsv
5CUoPXxfoUTjWP00pHb2Crch/yJFdVPxfoLw2tT2gvFmd/7l8VSsgNOY1AYXwHFq
hG0F8GTWMHOxjHKTXvQWETAzPLVjrRK1aXq0KfVsWaIGhcDs3EXJ+80B1ffMHTGL
MHx5u/5A163jJq2Zxpc2Q5zHMDhgetPrDzldf1UZ2kpIU/OdWzk93YqW2r+vowu6
CsgL2rIIgEtBvvISoIlte85oGh0tIlFlTiIiuhPPNjn4XhD5yuEqRV+w0Pmfd0gS
0Z3Bj45AAtt9Ght8LLyNkNlKcHEcGSw0/sW7mYgB2krfzK9Oou40sN5TjQKDPZyB
inBOPm189CyCnvuzTBobsmLL9pud0P1PG6bcr579HsYeItVQgstnsMrSl9NdZD4R
XAsNlHuqU1LGMStsRy80bqGg4tCcfhiTC2fqgmnlYCrG+drnHuZwllpsm2QfKBKr
jSZeHT0gn7Ia9rJoW6PvELAX6OjgcCbkxAYYSRVwEJIQ7+LXQpUMT1MuDpTmGHiM
/t9wNKDtyfhNHv6mpGRBwTdtqpZZwAPu2tBXvWm3wcmoKPoI0n0Fkx14MumpyZf7
7lnBqTn4vU1Oe5adIxXH+pfJq8jjpctIdAokSQBDVGa2v1Y3ttwVRnUsDhQN1XYm
2SWBxGC6gAtk1h7uBn2JdEmex+NSBC6G5M8Jsaj28dyqzoKYxvPHlq0HPKLhvJZA
T2qoiObxeg98uLRjlgQpRrNJCcdb2XnlYpLDR0A246eJqWud747PeaBoiphKwQ2s
A8LtvHLQQXbpSlVlCGtG5vSqRoAEDZkFIP3FzlQWnKzDkqSjjeGjZDadnRZgEO/o
/dMLDMmF3dJJra8pLRHkxR5XkUaVvaU13811DXiy+1Ie01sYWPpXmenZLNYRTkAn
nRsB43Mhudcha5jZ8RZHamHhC/5hPf2aVVM5CU8pRIm3YevU0FIVVjcTLFIzXKeA
LJnGlS7DP/u7tk+2eEVbtnG3dpwlrUxb6gFrkqF5sbAPVtMx+cCNufc6dL2xDz8H
OZ9M60F80oxlgaUYRK4a9EP6sVQUxiR7+jZyLwGNykuALiGWsTwC0mLuOZ4VX6U8
PP9IVNC2hxOjc6LKGk1QN4nZwXJuJsL4/6waWRlYCN4vxbb7YCzhzEWFq5WagKUB
Vzc5X5NmjR/P92J9xdUu6uu8u2Fi9CittvD1/w09/A7uk7KL4eaxdoqEUxfHvTD2
gTHHFquakV4ydllrVWn1ZnfS6rkpk3g9qK0S0lge2JKTjDEYiUKBNcXF8Eg88orx
cAIL7TV+Di7fjxRkKn7sf3RMjuQk409c/TXIbVEqMchaS+PyHezjJWyzhJ1m7ZKL
yxQaPvNT2cUly+yYNrdnvxqmEbdrV7BM0eKtWrWc8JXVpO3ewD7G8IbjGmH2f/Uo
hBuiNAtuObx+5XqitpWDesKxmk7A2VKNxDtrrl5Lbc8fNjc9KiHwKjKKV4OEiJKe
4owdl00j2VWhWkORreg9PncStBxwA/jnhiMGJ929F9rCzm8bKh9sOwZrX0pEEYDE
AX6qurhai3BPNFHgyKQOUny6z1sLPlOer7hmATRMPPovMoKiJawkaRQhpvFy5Jhm
zwAgqc5ukOOZjGaqTfoiF6nO9goI5C4jkOxi+Ze5PIT09Eti1es8caF6kcR63GjK
Y1CcU6zECgXZOeoBvQWit3frnoVSyc6wS9kTQtqjuS29j8YDKLNKcptyzsFQter/
Fv7lgA9m0zHHtnFJ4n+osby56K9ZF/1fvdGfloP65HlDgKQp3BK0Qf430RJveMmp
DpkGivTA9lXdTuJiHnzh3P/LzQCySB4piuvAH29/Q13h6OrLHqYedUDSRwrvOg5P
me2bsoppPWZPtdsjQSjRu7cSsJUYT/cLzdBmIS7/vt1PyeIAWtr2jwDszKx8WfhX
tAYmwcl4ZlwuWGRa2cFN/oGrhzGSe1dMn9P5ng7A4XQ+Zv/ONk6r5SitBfwN87Bv
S9/pVxc9yRLn3nUVkRHI0ciFfaQ3vdqFOJqA0o65If6+G7OpPqvzcNXAQpAuCuNz
K6Z1+cV4J1eXCwnb1k7+xEoornz2R4ScSZ6/szumcVw8cI0tGCQO1q7XX2Gd6IXg
wVJ0PLw2/MLARSQ0aXBHyqU7r2O/c2TnufpsHDRTXR+4HHxryQKmdzKUxI+3wpbP
SbnFB3Ryk0zII/f0ekeGkFjjpQt6eJ0Pota0cw3RbTtNuc4JPuzEf5Lnxve9cZLt
dhMNdGCo0r2C2xaF+c5R8WhvZ6Z5R7eRPu6mOyMaFFkJFVaUwoY6rUL4EHmEq1Hl
IdYMQOWMwERj/EyoZbAxX937NWfgzLMUm/BYhB29fB+YzKvgKu0bBEgRZ92p1LOs
7GM/+F/uQwHwyxTmmC9b0IknDh5vUN99G8YEVFhC8mtBJdTzti7mMRd5v/0Wz0Qq
hAQFKk+P2ULcdCAA18MgPhTdOMUtSXCbU1fwXJqGOUwk1RbfQ8Yuqvw3pbLrmE1b
UPEB85epQ0SRya7vxSy2AQ1QZ9IKtwcVwx71gJC7aFYm8TgZQRuqdgFULqPRWFVc
avPPrtvn1SZPPAEE1eaoyhbWC/9WXYOuzwH1d93uJ6FfyjOXbCpCugl89yRzfw4M
L+Z9OUlaPqZMpJ7YDVTRzS1mCLG9Mv43WzFhw/ILL5+7YFLpJzwhryo7Y9XBQU2M
YQv97oioMhsaaneMkhZkbeNtsQXXv5GY/Q6GIx0ImdN+ZQHdLZZOzulXiUeh6CBk
Iqg2MUHMBg4BULyZJq5FYz3ObZd62uJMxatKBM71lhQsKAvhQ9ZfSPt1Che0kmSq
diFgko5VSs5wtaS20JViSAmoVEB69fuvpqrtr8H/6DvkT37IQRLy035DIlxnIUW7
a7Io+B+iinwHPmOkx1eECxzNDQQdg8pGcaI71XVHzQnH8UQ0fI570koFkXVOCd/n
L7VXSF4JAOc9inQX5k2k4OjHH5QTSPomyH8MkavmRtQMdQ7K6VmAjSmxQCBWh2KE
IIh05hYnpAajcqGHkBx1IvwmlJA4Nnpi/vVTX3GqvBMMcbg8kLdUyXGkz9TY6jL+
LeL3XNp+Q3XzyJogfixuuv6wtiFY3Y1/tJmMQfgaTtHvzVBie1zmJsspYswOBHrf
N8n2vl/f/Zmd37NK+kL0rimKx3fXcGQmmxGBGUYvML6CqG8MYq4qFDAjaOn2tUKg
BMZsvWCC8VHOLm0yF/gLGCyHhGTMkpZjvmjf5B6IQmFMMfasaQtP4oD2dm0rDJrk
pr3kE6mJaB4rFjf8MpUlM93O4YGwMbbxBl7U2ccPLLZo6uC2oQwt9gZgM4ojt8Uy
oBjLd2ubn8fB1kTWriJ6//Z41kWLkdFDN7e6MdjzUQN6h56pR4SbgUraFAXxbacy
gg/iCnuSOO2XNpj/N77UIhc5GV2iggiY0aU1QFmXrCKQD1k1/64fgDZZsXkwBACT
AfaqFN9FyHeGNYk3y5JdQg42Car8wIg3R7EdC92lLi0x8egTrcolJ59bkr88NPBA
8lmZ6PkhcX3XWzhh4Y6Hm/0PVTH4gqG+Sgq93pp54ryd5to8AmBqD9vo76lAKhJx
APOGxJW0Mm3p0KezekASsddhK21te9+F1DzqSEog/Ihm+e9mk0KaTvgkjqIShXBk
1lBYsTgYiuItA85/Lj6j5qZ+w15Rt3jeSDhwH392Jd4jex3R/OEz2DvviWPOzQ6l
AActr5tiVV3UF97Zdn+evVmCGqYPTfNB7ezejUeVBH9xzJ80jAVum7V0IMDvI/7+
2pk8Qp4Gj9pT8EdQM7OVDmrJG/eWGSPtZe/XkzW2jCQrjKNc+FxUnmd7F1GDH2UA
itNt+9K19GitiJaTFunDuhWYhQgwWsctSNRqJ/Oelx0vfQwDyjHt3rJMCZgX1aCG
uwPG4S1ex96KmPgIVV/QAVxrqnHGRy338K6pjrISesFvOMRLMefZQ89RcWaYx+XM
C5Jqm/MYVbxiuWBNcpy4ALNolalVmwMeqh6vRRKOPeQqR+Bvv9hnZlASM88INLKP
c/blTiQpYdIKEmwIzkkTo+SrneupEangNEXYhNLsCUhAp0eqqjQBD6ITY1GoDh94
BDzJeJseGEPXhPQi27OW5DlRLNN+roD3ClLIgC8VCc97YhPNpCKI2Y5MW+9IXpq0
+X06I+IKLkaRaoHz+SmQPD0yZOL+367A9cA0fceH3303Wjg8HRdVaKWw7wzdl0c5
1dWEl9V/3c7p2yVy4UhChFXKxn4xvoxWy1HuFyyZN8nt541X3ZeVI2jIMhiNKvMa
BHdZxxi0vRMFkA4Znze99zctFsiEvtprZ5P+0GnCyXhBls0c4FnvLU+Gsx0LV+LD
QVdNfz4yyNGbN8uLkqk0/t5lqAC7QVwiNOat8b5OKMyP/CaSB8FyPW3lG6WvRLpH
eWbqywrl3BkC44OzzUx1BzLuW3JTQNtBBIZ4xo23NjOPBV7oT1Sf62om00f1UtVo
NyeLJ5W0WBx50APshHntlUcMBflTC1Y2Usg0KUuin3Kc4XmQG/2t9aqVL0QL5Qv5
1BrAlw9U6BFr5apiBwCN8IEhSjM7Y8HzjfzV+gwUGpQsp3ghZT/nOVLS1YaQ3ftr
GfnNEaFwkTEEgB8cY302haa7P2k94mAESCCxC4vO6ZOPP2uwoxJvJ0avguWTWS6i
LbQ3cMvYzsovwdj34DdIF4lU5hn1OGl8AaMi5NXZzyfpL8cY0DBh8urFtBL8/3Av
++NmdR3YqSVVtgtGUNPqK8zFjAA+QQhL/q+AP6jZ3SKLRB2z/NZYYEQbBgJObY/9
YfqpYBTBB+1tIykbDeLul/u0zB9k6wx0nlgemBKbaEWZ3xFlwkeNlFADGURT4lz1
yctSGjLpnJKbrBmUD8wRRTtbunAzJjCoNrEm6vGSbJ0wYwkXrnHfJwqm3s1Y/EoG
RAPYEh5fm6gtOsy46lSDO4ZXhgx0dQDLDjzage4gKe89eV6kvq7BxagkKH9wpslP
xWUTRxaXP/z4xU76RwsgFMKMJIggQ2kry80KDv7N1Cy92+1OiLLuCBJqd8/k9QMv
hWCUaDjRLCFAC3LM5vVG+yNegOdXjB5pZixG1jtJz0cyjzEvnUGIb8ubH3brP4uc
loWXl7T3MEnqAsqmavB+LsAEtSUy9u0AgI1GyHyRgkmuJ3NOy4CsUpVBfwRkQxxo
V/mpZu3ZpVUke2vosAOKgbN6SsbmdEXqJ/+rzxXWARGKyVtVWIaAHW6E60kMD7V9
UehjMCu8/57uwSZrwQU1LCb1Y2yXj3E8bpSiVwPJLa8TO/X1juNePnW87Cc8djdu
GrF5bWcx+n9u4S1dSukANS3Q8zDMYgderjAc40MxHF8BP5GFFjQKcb9WufibnHS9
qbMZZftZ/4wXurj1x7+H5v4Ah8ehTftYJ/l1plrcS0Rt+ifsoMtbiQ3BW+yes+TE
UqNIikJLI5VjzHW6b8lfXFInWtHfmwx6FVX6UE9u1x9uew+v605mzG/YggUpXWqr
N1+vHV39ZFXBZnZ2pOFT6KLY6LqTZG+WFS8DBVX8PeoZJdD1UKRJIgYAIpE/sJ45
qeZnrFgGmm4xVq19UvnT8l7WCzbfRm+blt+eKLKGUy5P6L+4nMNCF9oVc/x87lSN
kI+JyBdlkS8DnFdjPacuA6e7sYJkI598rg+9gbd13CzAF3fp8KOmMIUddhPwGMoO
1rPZwANU5qSauaEVg0wyZEK4ovHrOQXutgifK+KjrwtV7M0YTvb9I9wuvJwhPUNV
J94uPQWVjN9RNvBdzunZt2xZVcCEWNc5/ZvUD3k+OHOL5MnDOBtFFyj3uDjprwOX
WyfC/JnY0wCfT8U2V+No4K50UteDiw4dd672DPLDg0CjY4Q7B1r35y3+9Q3pEw5a
vabjoAXfwAGCvOTqkrfG/jcxdc3c72cCvCVTIP4FqA8mqbMPrXJFRoZ5lx2nU+r4
0aqxVW6UrLWA/4y+MJJe6v9Bl0OxubGwwrmuh9AnVyHYazQ6ccCQyo/irfS7ev4n
2v6z1QDpdYAc1nBCFMhI6N/1C3TpLGwD3Fh0hss3fuG563EgYJuDm9F2rHfjCTPS
bEolLiqjwWgZLam2rxMYXVJMe39b6Ms6V6ZK4i8dTs+8EoEktVrsNFTdx7td4jQb
jeqyvfX39zuT7rJct8R1JBPGp0v63pzci5IGuFaCab7EJGbp3hsLrqQyifN9NH9J
TAm52kwRD8yZ7Ms2QVJj7zCb5IGMVXurtJSaja+cbDoOi2W+Kb/mJN2584ewK48m
XRpRlIHrgkRigkmtVGytVrA5dUoItpRPzPl2312hlO7vOltBJJtVRaMKEKroINfn
SqstmKRC1pcgMlFPx/HyLHgIU0tIpJ/KX8A8AhUynJS8WPMmMK1KlyGTo337NCT2
dqh9Pxpe3VmGNZAUZAaCQJMesszbZpEHLx7xOEqK7NOeoSlPsLQLlhko0A+XMSQD
gwBLNPq0/K0kTsWj8tV9eB/dFipHOpvPtiENOrPZYFEjBNFFiPOMOjY75KYDpS6N
j8YwTnQQ9r7q9JGdN6VK/B/9KHBO/LXd8haBHjH/RORGY3KyjexwTNiaDt/EcAxa
Z98DsX1AhuO2Dq9ElF5bGSigYmN9Ucz8HBxi5QzB94Xha9/OiP5FccNL1mH+JJvj
gh/3Dh7kush4+P1sB1r8ypytgSzGAcaXrVrG2M7bSvSGtFKRJx59x7Np5IqfTXDD
AlNH1F0XqaUzdr7u+QwDpGIdb7U2IWWuhDpp/d9gaYHBzWqwPU2ss59CPEyNSqBd
sm/LCvI90CMEJGc/6pNE4ynJ5/AIqgu+rUbvLX7AmQueXrmS10CfeG2qEJYZML/U
HhPbYr2nJ2Dea373dpmRzQZtbBHXhXw23aHT/KWSozfJ7S/MBH2cCTwvuz15sOLQ
XEOynoni+WVbkMFuKfajy747f7f5Zj+c4wpbydujO9WUPlMQlVZRWwKLoM3bF66P
4555M3AXPlhK7fva6ms+r1hMM5ubrz+FC8NDMIVVSVOympMhUxMlANkETG21LspC
4JCGbd4NUWrvDZjOXtq8kWNwrU1+fIqve/KRJf/XV1/geOw/qrHyVIEa2cuvp7B1
IxMXgojRGMs9tO8tIzbm8KDsDKC4jlnrUFfx//inNCrAaht5TUET3u6aDPyrG3nC
p+63XELYfh/0P0DYfAuBQj2VqBi38RvQb1OTPTLSpjhtgrQDZWLXOzggjfP/IOOI
opqQlLmf0zfSAtMusQEl828D/masJQNW7qRX5jJMjwm5bfcpsJnpdvIxqmx0TwrW
67KiV4ZHN1GdCivK4eGjslOkRDhPfIB+p/Gq9sZKf9it6wq2p1IkUIeG6OB1leh/
CzPdm1L2ziQ3NJY8RimY7yawC36mWgrzVRidJ0OmQEEeDl2oZGa8jBfapYcqN+KI
RjfHLfmRJHUvKvQtYgh+Qwqp8ip9L2cySldeg0aEct7t9DA2+9C1gJ5tB2abF46H
CDAngabUzXHIJx5vj2eokbjYZx9fTwez4VhsfNLJhHUgNude0NCkc8FZy3kuUGvL
KmcbRl7lctsLIA8ia97phE9vP+J3KA8y219vuv6FCLZsfcx37pR4jVZwp4aSweP4
r1Z4sBE+TY3NsNva6pGvejNjZZouPnTFE//drwR5g/cMGt+zrhB6UD7MsRPot6dd
AAssvVGOhBfASqxDuW2KHz26gGEWraX3SQjbKkzP/yso7GhELopGkTl5tQR+1LJU
m+VeiERB39E8TrXevBN+soXcdGJsUWyCl+hxqlzmlWXqT3Hhx97cvIN9iCgV0kCH
XkUNaxovqPzJpsykQApOaSQSdhJuSq3iGQrbXg3Bs+SoGJ5kiNWfLX6rKoNHhAFn
ENq70SOdJJ0EKFrhZnXtQR6+vvdqo9ZTaw7Szd4MW+VAN+aUSiGJPtmBFbRetrp4
0swt1Jw805VasAs3CCxAT5lNGY0+tXfxNAGxfxhoAh6/QqGUV2V+qq75MSMJfpBC
ndAsTMIL1tZPKPsbk8ZKm8Ka4rlyTHgkAZbGuAwzu608vMk8+r0P/9k4Xo4RJKuD
Cqh+MxYVmvJJN5nW+LPUvwCOV/pl0NEZEF6OLBPDCf/2N3BrBB3qStJa/7U+9ATJ
T56uTSQhVP62md7F/Fj2bZ+SMoAfEiA7X4qbE8Qq/Ddec3hF/0s34bxIQZu3MV18
LdbgebVzgEJ1b9+bn6YmI3057ZsUujAru9uREjMyO8uhsloJVn/ZZWYlpV4Wevo5
XQamjlrJTt8NRoBUUXNUymXuddRhkgPTGAdnycgIfjEWbVW32kio0t1KzYDcuPgs
d4isNasTw9x0SM0ErDBX2AIQ+1Rj8yt5a+s3oJX7pCt1spyeN0gLOVvXxnOOX8fx
qvRMpTgHcvN2g+TWy72OLMCXAH1k9106Ps4pmyrbG561VO4LJPvmVx2GVjLEhrKf
mIpFdkmliV8FeqiLfA5ZSeLMGXy+46BT0Hn3t28bEmbzbAW+/w1m23xbTVc+KjQF
QLZiNeEvKIo0V3+JVxq7HRxIPZ8GbNHIXaoMl+RLYccBVLPBqU8jjfzmMnO/djie
Na3e8/awKwIxvQPoOJclb8dkLOCY2j+52needSqj4kyKvjo9jPR8N2/widqJfSkB
UNkm8Y7rvzKBRXX/XJIyzl2hAY6PMd9CJ8IZPPD4PTAdu2rfG7+DuZAi8fi7mjTq
9cJ5xOghEFimq7iIopFN+SxZq0EON0KhyNMzX3qhsxrHsCRnIWdt6fVqDGtSJ+HQ
z4QRF8QyEll36qO2jHiBBxSuoUIc0vFanBwR8P8nvyhbBlTfz2YTk3qKRh3AxilH
8F7xvvIcRXXGYpdWJk1VISYzDF35eQ7sruJpkc99VYBecjZ+w8Cj7P9EL5YmEwkW
2YXrp7RtjYZ3r6SALsCME+cX/o6ScQ3E+NOeeoRomOdNk7ktgyxVuMR2CwJxQRML
u7VXVPnxREUPnBMkSm24axnStn1Z7vrVRkQkQb1wkUf13kGzojQSWtB8i1GFryih
lzq5X5GI00fiB9BIyEbayppUsPkUTFWd+3qWbh4SJYHCYn+vqMY34GF2whhU25gJ
WLWZyjTgzxvtKEBxxf8SiV7kb9xzq4GYkknLXj69hk/BkJ1c3kWes7anqGOEwurR
3XJqAOkzJg8gZ1C+nuH9lJ6nlIjySatdsmQ+KBQ9lM9tsgq7PjuN1dqNyxpE+Q2f
HshNIARHNmEyq9BI4PrICOg403/FXTDH5vIoCzjDFykMIaK7mKz5fkiCQVBgwloa
vaoWbTURzTfKSb4Wid+WaL6mqi6JTwwjAsVHEJC/5/f5NCL7/tdhNcGc3Y7lgyyE
w3rqSrQWjhj+j3WfT4k361fqOHiggMEjY1fUgvqHxDaUH1eD1W99fQhInhheeB15
Eyjl28qBWWcl8ENtu+V6OR0lLdqYS31VLYLI3ifXdYc4ORKeNMXvvbN2U9HxoK5K
e1mQ1aYUL9aACG8vSgMDE3jwwE4TkWNTO8TOnh+BGUU1Jpg97J6Z9UtN3P64IZDH
zF2PqRtk9iv6qyVlPG+1xmAZij4iPptTQA5Txh5n6/WCUdE2FJQE5uNsefNfDjXD
cjl8ksK8gEHngmb5b5Lb+Xe2FlDRvRDLTvU8C22tpYKGBbfZTQKUyDbA6Bvooy2o
ySgcD0qq20vsRyrw6kVW6XNaFL/dI/TrpZ18w6Lm17BMlrJK1dEyBLgWf1CPhneZ
JAmgrM8hzz3wm0r4n9ejAXCtwDo/3i+4w3xQ99CAHw9vQgOJQR2uX/SvJBgft5iN
nTlFAzdbwbVX4LTUCvbljzLPnpWzNv/1QctJBUNjMptmX6oEYBOovOergaBvJs5v
almCklFetab+eScFBsFXcML5MkbmP6quJvSorVBQgsLai6XXqjvq3yWaLIOxnyBK
5eQxp5XeDZpUKYjLCcqIzO8v/UDL8ZJhQ3ToPbCkxzZcFW1YSSbJ91UQwkAcEyGn
K6PSbJ8MS7+0Dcvp9xciNNwlf/MgdX0zUrZ2FBL1XjKlLXVTA9f6kIrv1esncKk9
j0o8Del8+oa80vnoCeRHT44TKg/opLAmT9BMhCCupDCWQ0UbfFUEFKpHJNuIeWTS
tdxlkhIKaNvuFz9/0V2jVShLp19ZbB9+qnv03Us4DvJ24cEeE37qPcWA0VRGYRPH
YGbPI5D2WiiVGYH2GRkncrAGDrpqTTFJD4IDSEfpZ72/zKjIRIS9QSRnjrPFSYKs
LyI+sAjKjn4FZ3tRnuM89a2NP4Mm2Z0QoKzTyum7fyuuEREor6HCK7RIgHl8h8q9
8HBwRV1H+jEmnpvwy9p2XnzeGOVb1G2zJGpbp8cp+T8p3oSMg/M347Xv8a5it5U0
jMnO++qCRi0CCWq/wxk6GvtvxSRqv3Emb9i1Oj90bMJIpDH9yga3cNk9HH7eN6Nb
OAxcvV4GVcidcDOVkOnJqwCBlwT1qs3OQtXEYrPkNvv/RmGB6+687Cwn3b5TK7/D
6XZHb2ggC4Uf2eeE+4E4avukSHaK04DnXeOiVGzxpupKiuiGCnI/+ttU4pKmWhUM
AadqkXad7v9okxYejwpvh9cfyoXEV1xs9DCsVh1XAo3HuMpZWDuL1oK+GYErR+Qb
1FTQkw10bihvlTYAtcRbYQsmxIv1HnbCXlXxtwc/4hRk/xNpbNiA6Zaz5IBoKz8E
Z5qElhBt519RwYKSixszzONNuTSx6WwnszQh0rR2ltNhM5kblg+GbgAwVQD0hc/6
YRfsnUotachKfUl5VZ52IDL0rwDXAFb8gaMajqwHuJb8bohahLI0LI25QUimeZ2s
lk+GFMMF05nuEOAhAmYXB9CkMFCNZjqSrLuriDJcP5HlDSl1YuoGJz8tCW/Yc5ck
+6dk1w2iPtQRSQ4qR1CW3vp47NyAmIJf+GDfWiCx0UTRwS2OqOYK8ygApk1jikI7
OLQ516WX7ikeKMJMnHqewB2TkNAxNabny+NLOrTYS8+6lPOFzXrBlnjM8Hry1dCl
7PawV7DLjvRADkYc0mHd5OXV3b00xYMCsFTS4xte0c+kg5Skv+LHJzFVKnFdPYrZ
3TP4xPvLTpbZKHbaCnMpuCxnA6g3h53Otv4wZR8MOcsRtHcsvYhJui1POIO9RYp1
JIbJt8CkSM/2z6Ta6b8VAKiRkdUd0QgIiGJexl/MTisfU/wJbvX+F4FVE5ihBYV1
kmsE68m0L6p/R0H0WjlR6AA7i2NYa1N954yBdQ/8dGa9cdUEyio3q579+VyUspN+
xKp6u0QMVznSUud0TOlwkxYcw2Bfx/ZEiDdMVJLR5kCmit1ByWhLoc7Wlvxhncqq
yppP4jYZGqdbW+GNICXdQaemqm+VHPYP+RM9MK3OL9V3hgg4jdPCf1afp4jkbHRa
Ct5qyU/9dBotMt5Kn8oQQjx09hJ8wRRoQlEPQEKwos3uMVq4mhnovXYVzU6DSyhz
oEUZyHP5WM41xHWY9QxMRND4i08SGFMzwpC+iLZEf67lMeeKqPybkHfjlJ/TE7y4
a03+RZ1+5lC0pAfGwrGw9AbgkG+p21bIF53M7rxLdjfIIYDvY9GW/12iqF6x/peG
IBG4+osARyVVu/5Reh5VzTz0QBIT9imbLBDjaQyA4bnOWnwfXLsGyvjeO8hpYEZe
rYcNUJLqqJH+3ckvwRI3DBzfNmRSdVoWS7s2RKImMOf0MVLbmd1Baq5NmvzjoZOf
zEN1E4d3lri0jfhVeNAZmVIHlYDjmPtSnj3T0QGRxDq4TmGXqbl2fD/eDBC7Skvk
KK17ua0C5QdYbz9vQLis7k1Or7drs/5mlcJFSPAGkd1qY/Em84pBf/kP+ss+tdWP
qX9AJ4P5dTaCDCDlYso6Tjl9PfPT3TJJFgWeKLopmjx6vbc7YyCHg6PmHaSzM111
dzNrhNkN4TPBSv+ROwWGCM76QYBSzMGm9esPfXm87lsQ8uLRONtMDEc8WVGvAnF6
5kX117aTnewA37JwZ/Eb8mjSX52+g3tLaTpk7EOEy+kOKpyaExQVV9j2/rnsu2eX
H8tpFeTLmkuQfCHoQRwXbWSRh/xk950zZMvap+iR8gvfnhUVJC6OuDPqDWM9xy33
J9DuRN3QpwE9JPLViu6wYX7pjmhNwcesedp/P+CK6CdfioLA7HcEeYFb1XJ8nlta
NiXI0T4arLPZ5kl73EamAYec7DMrqWsiVREHWKSCmNkcfdB8cR2gUzEvDZitn0RO
uZg93DTGTSIAr/qKPscLlQveYqKzbIz/cujZ5Lf82baWvzmbbHa42d48llHU77LA
lqajsfR3PtXXVwe5ew3WlW6cU+8OAoP9dl1njyG6KPBYuAVobzIh/8S/wuaTOYro
QNwQc7Gi3Y29Ma8B9OpO1zWgVpWkLveKbgGS5TjSLluau1IEa852Kd6VGvgSSXWb
APn1KyY76WT9rjPS/I/9Z6HzBVHt4w6maedAFu1SMLBiaVynxcSV0MOjUP8mKQ/M
vWZcBItZlbt/u5qz3/zoYcQWlmEmqfsSeNSe/IgRf2vY/g4ln1+B0cLO34v6AyVf
/MNW8MYyDffTqO95vOrQra9TvDy4MzgSjctwsrROtaDDHVauM+uZdkoCHru9oKIJ
5CX7SdHPQfeOz4BTsUHQzxAX+wwtesSaPdztzdqFIZGXcmj6hTvnACNBrcHw3OcA
zKYDtdxuCZyXMjH0yGEXHi6S+wIeBM8p28+mw0ENFgCrRcEUatSPxxwb2udRE+hF
YKGu0wcUsQDH3fgn8qPf4HWLArA79p0ijIWVhmNiGVwFJhuHvXKHvIXfoKq3qbL6
QmztGnCoSx5an2yzix1W0DV/A4q4NMX7ZnvL/lDWIL2IIgD5aUd4oEZEICZmsdEJ
cE/n2WiAHYa1hQOr8M0FWhiiMhZC5uIrQwUhkh3k9+ToyC6MKZXL5sxPKckFfpjW
+ZfmSs7k5IHsQ/9dV6SVsFooxzfFVSzKqg6UWisfVk/pB45YbJZzXSEePR/zhDX3
Ie5UiyfmFP82vBGtnEQ0csXUwNt/nY12sgGZH7lY0ROzL0z7vEktRZPw3ohBXqsi
w9FU0zqRwJaeV8PPNb9BQHZcFwok4MvHnA8DRRwfN57e/4LB5Ue/EwXWrR6URoyB
7K5+rh7xIdHaq6o54wvjiSHvAzebKeOZqy+XBhvlO5+03ylyJRsv9XG+zyI0CHi3
t/KeTYvd5ORcROb11Y/oRf7j9jZw+eiCJYxCiDe1fMSVIqIL0y8m2iob05qol1WQ
87SGJSJ5FXYo3jZ0ego7UFKXWoH5+GHkmH/ViuzFTrwxmQvXYHB67c4aI7mbxEOy
FyRbIUzNGKkx4AmGHV+ZpcTgYd6sMjcKrtTvI+8xA/5mEQi+Im3rlevTH+WdzEr+
pqewYDb0RSyWzQO/nZeon+B97RlxozCRz6nO4Yes+8PsOGZsZdHQUiiENT7wrkIM
iR+ixMOqFe8wiJnx9mU9Ilek3lk3xtrTDxUeOlYHUd4aBGzknvP6+EdqfflS1Hba
+jdIt02vLYB+ZTFIC9mdiuM4bDObT7rlxKTcOOLJjyumxmCzCEv2dU3H1Z2AX8ip
7oCDuGDjz79sqnUPMo7LYyjkrehHco9/N8rWI2lKqSK+hW/e+1Q2xPqzo5wGVDxG
Qi/QHYS+mhwKgi3PU5XR41RMTot9JoGcMs6ag6La20Bexe/mr+fQYi+hIK2gkjWu
r5jHymyuH+22XX3VcrBBKOdgzCRRII9bkwGH8E8boGbHgp7LZMaeJ8nAOUJzSSBs
QEQijGt+5wXHIS9uUj0I6Tz5+bIljkA/sxZoc/SfWyfJcSofsYyqlff7IayCUocM
no7y+S5hh+JukOzIVoxbzzWgndzTWioTRg3EpOKx/BJgZN5sp4gITJnHZF8pFJsR
Zs3MTso/oF9u1wzeBrcBtLLn4aEln2bG2egkxRe9qD6K4D7dUpPcsBqtlCE32n8o
8rVkzu99O3mBHbXxr9gEuohU2WfLhdXOGZrU4jWztjCOqZBX9756DcIgCayffF1C
kqQk69K8zMiFgLOPnYU0J1HONagnCuURdyscv7R5uYDyhAm39d7b80KfKdwTmx45
Hv/jb2AiWllLrx67jtAC115ZR8XzRuOni5XYz/rXxSjaRSETof6rcnxJX3hPjR8O
DXnBIyeM37MLWXl7EcrI+QtJSnaDXhdLfoVOYsgELYOhelZCGyOVaxSABShHNKgf
LZZsRuFbGfa5i6aiH3opHI3RbgAKrWPz+NH2Gbwk8eYAPgDzB30U5NnujApjmgJZ
Z+LX1B5cUq7nwI6eDRkdQDRc52qxjQqdRpM8bxpDjZ2HLNJVg00qkxcnTThwdJCK
QI7G04dGJTfkKfgfiYJGNAqA2rSAqywDcAWCywLgTeqgK/+FGYO7PWa7VXTgb7xx
YI7Kui2yI/WaHHtMEwv0Sfqkocn6cdNHuuBPVn+fL4bZv38+aAj1eM/rIxjko8bs
mUj0KmJa4RpyHUHQrn5V3xtRX+m1bdFlEzDVnxZIzjzsbMvXkIgNidqkZOYVgqyX
eK6d15uM028I+Mr4QLlK4sJCnUZi+Nn40UV6KNFvpSWfqjLG+bQBjloYATELIafn
jA6QZti3gS8PUhTdL1WZnQ07OtrJrZcFaelOa4kA7osNGNg12eYZwTxnkgy7huld
lR9iNjWAknnnjvAeFnkY+eymxA/OO0MvpekoY7E3ehFWd7MRvKMX7w3aLw72YUVG
ZeODb5oSk23kcp/TvuhtCE5QNTdxgIOIR15vJaC7tQXx/+43KdjBxsgXgsL9oZYA
+VTb51cZpro1db68YolsaDRtIsgBwxca+c/X0HbsOWQB/2hx0ZcySxtupLWd/Ybl
RRViWH3X6pQFVsZKVvOQFEIs5Kwvrt4h9JvDk0A/ju5P6as9QAXwh3YmZUHEvz1s
Cb/x3bhh9lwz7E1p3SV1mPiYe7IqT2/n5LF02bE+FJqsC3TmGYGTnTpAsv3cw7vf
PTLnRp/GKvlg2mNxg9/93DhNI8RSPq+ju3HcRvMqTZCHVYdo5WosDS4tjGWDHFGH
jPj7LkFtEv1SMxCAZv4jos6VUx5Xb69F7ox9kMlt0RgwfwzBKyAMvQTInf5d9JJZ
rFHmGNNdMwP/7UWPOHU/awZlnuVkQBv2Nv7DpRrUqeVEyZ1p8xtE5PddTE7OmUwZ
51lc2QWpSA8NP3IFGI/tphoXCvW3nXzsdAozGZu5CjyKr7JFZ9mAyWG+IhF8TrNw
dfU9kz6JGa7Un6sHPmUMo08R9Axuvvmn8b8HAmQdrHxv4L2iiTnvE+/4WTyzi/tO
IfiFiO6VPlw5IJiAgYNZ0G1/tYFQWz3tndlmmU+pnShTd45F25p/8MI0zG/pGp+I
Lm/H3iIHdkOOjTX2lSN+to003kqWzzQMczZ+NypgQ0NcPnKp+v3KaIa/S4xy4AjA
YddHUgEAr98+qS/68vIBJ8U2OJSNT+xVOx5YEhm2g277ENWHxta93cBH4uY3eR/F
3YqYmpCHc0tIsg/NBKEOkUFhmNdVjJLDT9ZbNf3LSWsvCdJkBao3Bt+GbOo2kKhE
0PoZdxpYmJL4rlETI5e5L1shol5yn1TM1eTHjaEzG1NLFs6QXSJSb+feYSPSZ6H3
wi6+wkQS5ayi35sMZS6mYTAHy0Nf3icc93K8ygzYl0eMCEvJXbnY/jTTbYa5aEDp
2ZBwcr/gvxha0HaLidsd1XiKomFjRRElb7H3KYFejvtosTkhMEIWYNbLcUK2Dkpg
2gKKllKPv5Fu3keAxrCyhSOaxiaKF4UiRLwP8gFN/7oF0+sH/AtMYx5nMR6LQ0M/
sM2en0kvCN8cigpnkY3vdmuA+2UATA9oKub3KLn/Eta6yvhwYzAxb9veb3tFUUS9
rGzWng5zvDAjhzFQJ37gdAWbMRgOcQpHYz1H9u7LEFhJXP8tndcrdqV6teV1VIOg
eGX4/WlEmMIPl0gdfLROlynMZFLSJA1rMvLDWvnxmVQnqkubS16nZwFNDs8SiTws
rI5g3lh4qZpBGtEMe3VAvwyW5nsseqrGdLLWmptlE9BqRDeNs3s0+y4tn+7dcA95
8LgSagnnvTLirCkTbT78QdJq8dY3fmz4vdKrq0qwDNEq2w5rXdiSofnExw51fGPi
uUCVEHZho+PuRSWZMus/fg/cTGbFR3aIzZs0M5fYkE9RMJeQvPsYgu8n+oQcWmG0
CROHKwwg+bVN/eRLUlsAu8nWzKYmUuN9Tk7Vdy8/nnl+0HXt2/XkVZILip0dlEda
+F+H+74tE8/E9Aw7KTbhKjpYMZ4Z+sCHa3F0s5EwOO0+rno1DNEFopgiUGXpQd2T
Uy+zecgqZ9zvi+XKQpUdyfdVTVyoHioYrcIT1cZHJ4cep15yTlbOrSB2ihWtRBPb
N7cNTac9g4WAURq0crzLSJD4s4oPpd7HfK0ThObrX9qph69zfhjpUVKeg1JMjjtZ
0n9XUXwQKm2HhTiQUVqpcF84JMNe7TsOobQK7npSGnYw7lKt45+8LIllrOLyvNH7
1C9+fNIek2q5uI/7UCaKqJSpGoaC+oDtnW+CZ9XDx+nzXSiJOvXRmTI4uX6F035G
SR7GcOT8+shzUj3cSj3WtYcYKmrdqFt+D8zYBAlVqJn0ixjLYTRTi/hY3tB1Ctgf
qG2OMeF6bnzsoGDNgoQN+ozriWRr4Bja/zBc4RtV299S89bsI8HnFp6H3A8lzMtz
/X7Hv5Yt1/v/91vD4tDyazKZtcNbMKDbcde+UrVNfU0FOi69J9sxARCX7d0ejz+1
2hDbzqoonXTvbc2nKqkYyAzKzaW0/DnVanBpVUWIWAjPy/FkgI6nbL9e7dhcVL5u
CGRxtXKTNjiX3JSW5iJDJS1qejWghP5dsBfoxj2WmZpaoUevgs/U43YzzFrWDR8t
jWWBRc46e5zw+LLTyLR3Lsbk/XjUTavEXY0yrzhLhZpzN/TjecRvrxsRTmt89+hr
cIlKOn7LyYWbnW1grYc0p+jQz5z7ErkjpbRxzhmfr5CEF+Bz8bHJC7cSha8Vg6Sx
VnauRswDmnjbh4k0ljtzkPotBDeH0wzDNVAHWAeMTobSxUqm84E0RdGBiMsFhxpA
C0AAejbUNv4uQwsy+ChlJaRACccFUIsy6h8m8ux0A3r1in3zhXEuxlNKjkJzpSY+
wdiw2nJcmm+s20yoWaS8b1Y+kULp8P45Iannf7AyzjrQNJ+qWDVYIhJ1a65Lsw/M
hxcchuYhXz6fWdksW+gBpK2XkqTaGLpmk5+UJ0tp1k9DtUl1GB2Kmg9GPPqlZRoK
5VwCUHFWQJdaMIypweSVaW1xsDVJc/iP7cPUxTcL8p+ULTXvuA+gR49LwFh5p6Iu
Cmpnz5TQmzyevpe0yjajrFKkmLAdTglgbOnQ6R3MWv80cWINI1Wau+sKz69o0QsE
26nVd/ZA3qVvusS61sx0HVesWA5kEifwwR+yZch5y9oRYRre5u14lpPkGSu1/d/e
DtETCHKzA6xOEXJhXLHdyOnGfUtBKyDRQmLM2FeCXsc0D2yb4g1aCv6Ucrd9OVgm
IiuhkyYOb51WArvQsc5y0IuR8G32rQNeoaYQWC2WFgaVElixYJE4TQlph9DkTvhg
18xHZe4vFF16oviixpWX8YbOHjeR8rx0UmWDi8ClFSJQ4RLRowsr0E5OdCBP6Ba/
jZzgJ+YXs3Oqo8XYOImFnNHeUiOwC1uHUrl6nYqq+QzHXsypEUMYPxfDKJ3MotAX
IltfUqCyMnWd5HxCAMmSdxqfK6QFqff66c/aFZ6tQEmcnvkA5ZHst3Rece/5eoHo
onBZviJwQjxrjx5/S2KiW8gX3rUsp3nEGngtwq2uSXpEsV5YFhpUAyzBYx0kOz/W
KAOgoiVAIGE83i9sph2oqwWow3gaw7PWc6/d3bPzaI9zNS7hfNRNVqcbmBHq7bUz
fhRqm1VpqdSM+OSvUH92duVobUza78gjVKTB4gn/oXfyjdcK3ZSbUSVy2aPRkTCY
5Pi97Khk/W7uSVsupISKQ6mqidOZ0TsHiAAh2LUirjCYBpOK2mzfbu45OIbpqMFL
3dYNAYF091Rsdch2+mfJONDJsf2B9+oefID9Pjqdaad3rW16RafFPy+8Fu8/gaV0
Gzwpc39MNd6WG3pLNfY+waa71bZXrn72k5gbUuUvM117WrNc/QIN9PggGzbIJgZS
/wvK+mSInZmVYqN8e/6QMWhozu3y4XUih/M+gzf0Bm4TREKdfrpCsPOIPeWzVmcC
jKmbv8NzAKXUQ23M/YwYZUxE5y4Z+O4iyJjjAUVdljGnJXINZHyCq3JJPj0sneRQ
b5lf+AEcaPTxCCxFAUukq5G8x5IsPq7CTFDS1C9kPlFp53e02CVWP0CCn9TNqgv6
rWEaRY7kerOj27ILgLshBkel69VWdxk2idtSsspGE8FSlrh3Gd9D1HLjUlYSwiNe
EICdJjXt5o2CZPDySQ7678ZRbquz7qfyKKdxY32B0pjgEPf737ENR5D/4GhhmLOK
nWJOlhskdSJEM2Lojlv/bhbFho4OQ6D9YbtL+cH0vxTzdRdafKZU/UICwxVPhT7v
A+vJElg431djCkEyOBNHHQcAlwASiUaJe/itMASp4SO1qC19rm3WMPBwzYFb41pD
KepBPSNXQBhAa8r8BHaJczk9Vf/fIzQa4ou7jEWBWtJ1N1o0DaSyItT3CRTEEA47
CkWoJPQFWt+jGm4v7AErNYnKeIp1BHhnjGwDDZA1SGPbAjoErViwt8JNvUpYfUxZ
pgeIhBuiR14YqD2OELWdm5niuPavUOUeklGMeM165GdzC+Fo4Mpi4AQUEZf3D0i9
n2t/I50Kq28jgS1D18FtIHju+VBZ0tHbTEXnW050zN8vKoh7i4D+6fRlSHbUi3pf
kxT6yIhdxobq/966TpPg1erT+rVNGzdJbQgqCRm6DZARPIONY06bakt2tIPg/Ko1
e8qvQ15wu8+bF4grolCMOJ1i7QOh+ElD7vxDfyzJZRuSwaQVMeeoHmQSZmShk7PU
SYOxAnu/QjUVM0iZ1dIeX8rZpLF08A8eqlkOn6HW0RpwibYqzAB+oZYC0CPckkTy
StmCMWEn/xko6HbeDzglWGhBWONb2eSNAiEpOkvJmucB4lx1tr2dYgdc7mXhaOoI
2586LOAAt21wGU1PJNHZKyX49wqS6/CMHkPnljMcd6u+b7xhopY6iaSMXwzE73Vs
Qzl8JTBM8Q/+EQag5GWsUnem5S3XCjLr/eqZXE85PJR2wqRMeK/v+wO62zf2eODZ
cU4/ujS30rSKFcMMDFR8PsXfj+IRiakTAkN/GUV92bazxUxmEdgU5KrOeFo5bF0C
rGW+CH/+pl+qyXmgGPdoNJBVWnb5KJZH53seHNFKsPboGfATOhxkQTEpohV32WGL
U9vI6pZWicnw4c40fiD5k+nFiZwbfmdVdVz30/HkV62r6GnDM1qoSkz0+EsHwmtK
IZGI/Gh5u2Hc9QoMt6P50IU2iM73EEdlwu0bqkzqBcMvNwI65E6tyRhvcGiDUhVa
XxWC8VwL64j/GKFRWbz28IGWPABTk5SspAQwRizD40SddSnZ/nQjhdaiVTxlQUjt
r4GFVtPBJDRsXcLXy90QLMeaG0Lh1LARvQO4kPXqECB7FYzcmJXRpS7XCUJTmKM4
UT6oZitdFMWjQPxB71aqBBECAS3o1jHCXkfv3QUJ5uKuY2FViX4wtVxkHn5Pjv3z
IgwptjYe8nUURe4u2WQKSMCp9EErp8YMIfFNxwPhxKQO0pPKYIlpl8h/JiAfkmg1
aqK65MKWeXUxrdN2AZrTXaV1GdjOzwAI2SmtQT2e5P8XzI7yB+ExB0SgU58FMhZE
2opBN9vh33h7s4ZmTKegSNKG2jJaUf7uWuIXqjg7z/CK8D3jAMuR9zwA8xYRR8nR
CzK0C1Cx9N8In/Ov/98Qx0elNRMCRlLRpXURRy5SOm1BroOMCXLgYlE0Vk+GS+Ee
rLIuFRlFnK6cTEARP3zFZ+q5vM4Tbx8+mSjpykLCstwBofGiQwqCQPmEOJUgK1vA
YuHh12MONReRck4lAuPg2IDc+Nfh8xHgF7USm5Gqhm4Ped1KBYglklPd5m9G14vh
Hp0dSE/2UBFlFRUZ/lzFCl0R6n8YeTS0ztMz/PA5Aq8v2FPu8NOCKaX/Q/9uvVx1
NrNOoSo4hLPmgegPK8AxRqkQJDSle3ETVfU0qvijpHiifYLHZyrW8gi24We9vX9H
/6rO1ysHu8VmA6hFXM5IQeaFsrh7IdrMOPs6gmryp4QB0XOatBUkJgfaAt87WI5G
9bajV41KoAlCer3WH6qQlYD65wbsYd5QI3Z1XsaQR7BlcEVIb6BNzGtThn3YPwz2
byIRHhIGhhrXwrclUbd9f6LD3B2icf+8MzIcxKI7V/+48PZW6LEJnJV7ZkH7iD2q
gHtVMg/asWTImd5xtSUse1YVcDGBuRRMnpDRP6/6jZhKxh6mHAUo0y+3mYSAm8+w
ygGo7+ahWILNias+ETVZxBN4yzK6Ec2v6XSSfUo0mLAwZW6AXu1ZdswN/l115JCy
SQZtxrnn8uVFTG5CzU+/icWSY57kKqctEYepVz8ALYRKpLr6nnYGKj051PjUd1Y0
2WhSwRDOmmcZWA4jZN8SNSFGpSea3NBNY+n9JjcglPzfqCjiwYtnrz4vxwtJIDSe
n56XxM7CwtmUBrw/LdEJOm1SqzPjPoOz0ApbIfjJadixrGJoKV28ljthETGlCymz
2mICeloYmXJHVPBSo+woUGXG0/pZ0Tdfua3sBvaOcRamEknN3JlUpo1e/trR33cb
8asuua3gkgxdieX6UN46q4HsG7WRfD9RNSKmfpAIo9Ix5eoeUtYRm6L+57PF/wO4
LfbNbLBuJyTxs8g24H6wRYCEPCBx+VciQqHI1nLjXqFsgJ657r9qugGcRJHew139
83X//bPBvCcdZj1BHulRBkk/tY+W1ZZwPt9p9SoQeOJsU+Go/JKiagBkTxlLuhlO
T/N7EoPNamo5hlFZumINK3IZ2xyxjEUCdbqPFZZo3FdQIklwOdYqHzsnYa3+UNoO
rFAiSwWyopItDnxmYCExbcPu26ETk5zHY0TUHKNqqguGLFproqXT1pp/yPIpy7tJ
cQfue2uoRvpFa/sCxlvpMVzHUq0ytEricXhpERRvWC8woIW9tVBSDaWjiueJ9NBe
+UShS715GvITnTVWzeMOWhNTwIS4GsR0rJA4H3A2utQUy4bW0bIoLpM+9wW9mRsf
DHBhh968bKig/9G67j+2CBlnm2fw4CHl7Ak2qS92iH+O4hPAAPyghFtQJ6UUy35E
N5CTmgpr3a1va7+lv5u4BrD0m2mXl7EJOMS0Rbm/5MJdFvZtAGZRxw4KmSf43hGR
48Kv0G9oOoJyGod2aWiq2y3jCqtoqqP6e6vuQV8LQMgCbfXLc+5gfHnk6+OWeuQu
q5hnt0VZBcPh8pTbhvQmYxZaW+BGMEZdtJ8X32WrtUPdW20P1LX2BFJEk4VLNDmm
RGm3k008+xznrxj9pAZB0tAgDzhTdG5gZLj0XDiYXeKbLywN/Zt0KonB/q4YCPUT
Lmx3qlv+i2r65MsSSyTaDiHaeWzeyLn53HcWo1MdYMQ5Rzb+mYdmO2qRw6McsJGR
bizKc4Xh7/jaoFyz8hoS6HRda+4fbQL1BQ9EQf167vM8HPNDB6IAov4YE5VsjHZE
y8CInLMhKK6S/o5xn3Tehsk5qHwUY2lGXc7B0Xwsgfj4Z69KDstNOavxgW7m8UGK
q/qI+I7MBfCttSfbXb8aFrXW9LrBYy9AzLo4dTkWwCVQ8Qh6XPq+br64S+tvR3S4
GpA4vernoM1TePjQJCofE8BKJKLuXrKkQUrRCE8b4WTg3vcPrl4AQuXzbchLNgmZ
iBAJH8ZK2L0u7Vm3uDFfzPOkKBYJ6IhzYCduj48ILCOlwlXIJLuTgK4yPXfm6I7p
wR0/8L5Xoou59rMNFW3Ln89iRtakGHQG6QB4nMFfjVBW9MgOZSz4cy9uLixmr2rQ
B0cCAd9kT3Km1OgGf1QoOuH4rOAoYcvFVefBCgAsfMjAmoi9o7Z4ys38PCu+oqxl
CRvaNAPNwqOFuEjnZ63g1w2+mXf17fCbhb74GQnAU+gV5VsJrhfeawiC0AXewpYW
06npMxCDXQELYlkvhNeo/vi4E1gwRaDu5S4Hl3S3qIcOB66SBwoAuWQxct6nFO46
PyYZCptiTgUsyR8cdrxNEpQjfeP5NgDJuuutyc6yttfNucN4LmyvL8E4uiumqK7r
rDgRT89yORlH/q0RKiQIgCwUj1KtCUIE5leEAyLZeAkNZucP1c0X/3zgzZoR226T
Rq+zPIyFlNQ2za1jcF+YtQDpzRqsW4YPc0NUKYLaQT0Ia+3LkTnkLmMSn0VEpaWg
66REBhx+JlKqNi/mK2XEPEL8rMT3e0oQYaCqUwX+4Mx4THIXAHmUNwSmBOKJZlIT
6jZIOHTOa4ptBmlFUwzRyw00knJt8rHKh4D/q0iDI0BFR+hZqLAiNu3Xd68rRVpN
1KeXzdDyuBbSp3KJG7wqHRhWE/+tPHQhV30OSYwdldHNFf+7Soh/+yGe5YPHoqpo
ynS3gs/jvbP0HrkNWD4wlXjA1rmW7ok/0ttVL217Ms1OsisaSwVh3ZmtGI9U0R3n
T8H7alejMWOtTU69mBmbnhdLKcQ+GxcX93cGxiQr2YJUxbyoKej2Vv/uMYKo6IHl
rZqyrjHNpdYdzI43/uhruJhlDNauQGAZBy/QP5+J9lNhrE3WeQFkUmGoQY0zLbJS
3kIE6B/Kg7sOfd1WFVqfLrab/l9B5PZt6VjyRNtopfwFFnqUNpG+sVFFcCgiSQlg
sFSrHZiNCI/ggRwECSMKZaFwiIwjvQufQl7+Vu1aljtCUe5OEsPCFD9sNFQBmluj
NJQHotOVILK754dc8bLCQ52RYmdUD44dRtw5LxONX7+80MCwKEpt//tW/4jIwE9v
cA7+DoASKokli0xqdXxyTz0Mf0Ifa3dk7TMISFdeLxKawTkq3qxxujUVy4h72yoi
h/eTNpfnzFkwjI1Z6Gt68njghgx1xkylLX0AhIYSR+BsERZq+6S+3WBCiOWcnH6N
IvpuVn4bbYTLpGEcUkNGuB5bW8ctyz0igqU3bVGyU0MNJ4l8CJ0DAuXJ97dTGmX2
XR9BWlC9zQD99EvPhcWfM10NQywuT41Nr3602yuvLInwi5k+lKZLQhzAd6llWIYY
E83p+JLCcUrmjkG42eAIGyixwy99kOJOm7zp2hfHy0zAfhbt+hJuJMa3bO6faexx
shhkjnTHBfMBWzNggVp9nfiGvcaFdNrbj5rgYispL2rLuT9+NJfIYK5k2akTzB/3
gVWTNgaGEi8TVsqZNxpIE3OrEYW8LOmeRyTfkJzfF9g3swj9ZkP1rvcPiw2V59VV
cxaCrtmS36xX8NLzdPXd3rq+wf9EE4h3pV93UvvBqJYlFdmiIDcq0lq9UnToE9o7
cETX05GMd3SN2/+8BsQElwyw1XOEuEez18YSKQpATLn43xlCsR9mPK9hw9+Hx914
ejb6vtBh91lBx0dxfIcpQ+Y2PY52Ap6kpXuVRXOHeMbt08EoMWqmzHE+Rl64Mc77
RcS2fdAwY743EJ247aMbn2QGlGhp6vFJvtAbEqFVppjppD5/ye66zjWBya/IYDbV
xv/c7+da9u0O+Q9F2z7LwnU57/AvdkpX5ON5DNef9nvhmqxTy4qDBoPAzOocfGUT
6sJED/qWgkzeK5idHf0aGaDPc5v5JIw9eCug8bdvjpaDqiVjNi3VH98BmTx6HTYo
MYpgInntki6AwVpHhVtT4B1sK+OSam+b2i+alj1xgDSKf3dYOe2SoPLyLj0xRj+I
vTlCav8Av9Sl5U1NIPfVV4p+NBHQnZP0pKFz4OM5pCDK3V9EmCLu6PuA541jXSRz
uyVnm1jTmkyslraSILdlafdtvFiCaNUfHdT+XM4P4Y/LppIQDVWua8/cffp6vTW5
UxmqDW83ouaOZ0l8lt4sLKjbR7gCduNY/m8aeOhuH6Fx2RZ6qqB4yo5rJgRXeRN1
/bIKMgGLaDDdXHo50tz/eOtMoA/BAcWmOVyu8Wy7xy0ymwL9NXfEfNHD9aLpO+Rl
tc+2GsnVl1rhW+w8b8fUmFKibYTJ6ZOgoDbJMhRDtItRPpzKzqz/iF7ELAOk3jng
mNJ6clR6ukJtQnWJVJ+DPut6qY++ltvLI8sHosULoEJhu6I7e8EMstMsvJidJw5f
TV2kE5SqQtNKbcWrNyBAwOf266ewVmnTmlnrSYCpZg0u9u0WdsO05R+uAiJXNfFG
MnUccgZsFUuiXWbh8aArsO/0uav5iXgsyp4dGWLpDOJ+Set1ieNqQY4cR7HBKgcG
BXyDjL1swvK4AsUWoe22yHkPGdz3J8FBW7RVU6KU99ifRNVLbMUsOcXvI/+OgbTM
v1LYWvpT1X+LnXpqcEFaXBMzYthiMwTVR1DrY91x2kRtaxHL6i3S3VZmBlc7FH8X
zDTlXVkPmhPrqmPzWPZlFbwulHDZy8mEZrMoKAmRTcLwC/gBJ5LpPxUU0m7SxdbF
YAGys78kS4I0HgCe/YZgabGkwS6NsDYKFEjoSX6rK/C/Bmt3bVEFO2clhZ3oRdXm
JKUPuySP+zwT9UMq8itztehncNqdJBLppdLa0Hx8e5Rg4jcq4XqN/zujdJQudfc7
F6kUUtYYnpxBiO3neWrxPvk2WrIpFDuOxDScrnup95GNLsIbiNh6dzqTviABrz2S
d0EGlVvzPMCbJT8BhMCsVxMrisVsw52dhNe/Eh9LUc1Ct74ZfKRzaZEpaQrhakAp
3rd2THUNG8YE6B5OZkRW7DyzQl12f0w5jlex9m74uvXRbrQjwJKFJve0OIBdvfcY
mNuZsuLS34RUpeHLzruvS1jZOw+bF0BywLi5FFarw+JLyS2RFy7m6SItYPQ7bhKG
9aGTSjaKyPtbOksWI6lZsh+OPc3rqX2MCnG+YHMZomJOF41LpW7YFRdpk4KfiuQx
xLfZuZ54qfNPPaUe3eyXBpAXe2JhMORJMSooG4Z92J6ajSVp0wUQVaEYRPJSE2v/
XOuoWgyzo5uqyp1Vu8Vutos6E7OZYkxgsbdfcpDZKa0DByOQPX52B4seZORUc2kO
CFqmU7Ryh65wG7tuKtQTsE37/7nqOzWg1c6uxupNIqyp/s1v+Oili886XD/FLyQN
TGbClNTNHSNaR4ldy4R+oCqA/eGx/JgH2tFQF7xTiUxu0/bTj7VUVDyLBJ/S1vFW
h28UEzs+3Ul5G7a07csD7A8sMxjoIcb85M3SYG9lqYRmMW6YCtshKtILzhYC8nm3
PsfP/XTcOeFImBGOodO/3ACxre8fhs/rCpPIvvkSda/g3XQtn1xNeSTpHn0bNk3N
Fzc7TH4NgpTgzrUA31zg0ZJp9RK9QVI8IIBAm3cgdYRuuKo2tzfsumKjYyKm9F7L
rTjMkj4yU2jc45yQEFbCwyqbsZf+IpUXVpgqvC+WZG/d14qsvqQSY7Z+XgLCoj1/
HkRn9G12et0bcUAiGyDmfWHyZ2hUuQFJxVXVKgRKvGnN8mkBV07+nbwGR9bcUqp+
Kb01hqR/eRXykbju2HF689jUNaW10xQHkQOM8JgbzKi/B36pCSX7mdKdDdg/UpJf
xSeSuy2l61QrzwzQlI/KTfBmfLJtqDlXNx3ixL2m54ylP1UXiNCCr8t01pYod60h
jZRP/n6hifmO13LaLNRdWAyoXJjHKna8dc/k68HEPK9zphSny0QGm23lwhtVKaH/
S3aRChm2y5Yj+o8LOHpF76+0yLJ6QFVrcdIzDz2kZZ9leJo4Wzry9p5YqFK+ns+n
KtD1rpUdqtPLgQRbWPG907SKgX3FGUTEy77vmUkdzceYExveEtVEOdKrjkb8o0w6
97TM94osbUATNMlgtRTYKfOJMEXpGKhpYYc/VPm1ZnVuRYcoxIP70Rr+i5J5pDSI
SOccgBbfKklqnjRbXI3C7IiIzDrg7V0Ie9YbgPAfBcmgj5DdZ8wv5WZEbB2aZsgA
HMKUeSjiUf0XDrnx8t6N9kA6rFXvPrD3hgu04lgZR6nw0fy0KVHYsjYmXXGzzLPT
i7ZBcSzuhb9cwxFOrjw/LK1AVzDIdtXXAeDSXP7dJIauMChnJyCbCYZ5qwzM5vdS
XQr4zqlqJ29AY4/OWU2msaaBsC6ljZJN+ieY7djfhr8HpxELlGz/tVXY8+QN8h1P
F3N5wWGs3t8jdJYWveqGMxwIFLb1MLmNVDuYeKEHT6GFxNRlR2tiiqQBJ9F2Sb2Y
zxgnSeB3XdSWUA7NuWHMxD+na4/YMh/ARXCzyGkpJP3Ubyl77ebZDSgVXq5XJQ8v
D3ffXbX4SkJV153g4OTd0adE5rKIL9kaO+2+2ooE5FbNUHU15F5jv3XUV/QfTapC
Ng1nIe6u5HEeA0WS/lNbbzQfFNuY88ppi99LDUF5gFqzBsoVCbw3N4Xldn+b/UIQ
KTzWSw505kuXkhGmiYJUi+FhvtniFpomPBDPjEb2SX02e45KAo4PfG4uq9ToiQm4
nL1ugcBURZL9xU7LLn9fiV1I8cwgz+8J57qyx9eh1oRnJWJ3lT0SvCfx9MubsT8t
joop2K5+XjCzSL+S4FURzEpCiCYY3SPlUbnnJUSnocT88O2PEUZustqeFJu4O3A4
CWxeGt+YTpXQJRF984MUUBdn5Xs11Q8Uh5F55lnggF0eqAaSeH8quGx/tVCq38kF
22EXSfSdGhClFpUXv6wD+tqzd4ej/oPPkuer0wH89pGJABBXjJY2BfsU8M+xptZq
aKLXJGHqHsW0Q0NW0CtCIMyo7cWUK2HKk4AlohHDM2ZZbBXMLxaq5ymjgn5P7iJR
ccrfzHHVdbRJlsyb1cHpgpLCu6CZ9ty4mq54inTwqaj71sQDltUD4eNikOE2gqVo
gMRG3CSGX0Ebaf70w5AMnk2nGLnOdDZeUvn3xerITzYbS2g3OA+7KLPAASCYXjY+
m5GMh4WzgC7MmVSyvLZKwmIgU0IZqZv9qa0AFOABWepNZO+4eI+crts29fd76AIJ
UbQxwStMShJAiHxcO0QF9sn0YvSlCUF0CPw1e1TnEJLaJpCYoce0rXfkSkCY8pfh
fbUPDSQlwBP5I98qJtXAm79nIa42O1ggJSY19bUtl1rSZ7/ksqWPYVM1fkUWqXp6
5LrZefJiU7T9GtxFrNsLN3+drqk3nhIY3VuIIU8uYR+YtsfJ8e6Jt9KVtfkDhJAK
+64RbAaoAtuSOR7EVnXjC3oKekPkJPisZkzqjZnuoQhSNYRpYcSkVqVcwnhYWPbl
P69b6ktngnTYx0z+SxZ3qbfmcOcwGdDxAAA/pDYExc5wWZgA9tVVjPOAmf/ubZkt
f0IzwH/vyVmPSoZqs8cIp7WNyQE9DqihzL8uDw5xXseKqX2jhuZIR9B8dFQgrsIe
zSW0+pjNU3AddOUpEvkdxr+nRaTbehqLr1klebD/YBNnW/lTqvPYiJ8cC7nZzERS
SZkEgke1eTBViIVuQVMbhC1FCCFbhFAOrFkzkLWxddegV6Jj4NXYaFqKAc0uBeVQ
nlVNlobcsv7dgTJTBSuEsDLzKTGWSEr8+lNcjcN8P4IMoKmvK6bFBHEqnlXV+C7C
LevtD+uQD26PfEBvHRmEV/+Par1HvfXFn1Gy3MS+2sF+3zgqJ4x0HyS6DJGvWjof
AMk7rPjF5JitVqBT2gZ+ibIe/FOXolY01uFgwltFC+yZlw6nSYkSiqr4J4276nPW
aRRUpkxDWheVcLAXsPOxS84ozVJjL9VJz1N67j5lbLbi/eh1mAb6cXVkVZNncBAg
9kUcMKkMKSXZpA/j1d/xpWOpKaHNEMpW0LdTgTArj2xYn9Fre6VpConh5ubr6I9c
iOiegIzRyTJVNCP1FG6KLtlbto2IGspUnUxom3MrlBKv/rBAHhnCm/7jwiSevccA
7YscSdoyjxcZNSz3Bi0qj7GMKi6QEjkEo3KlJW89BKkt39c+hNIA6JxDYzi+m30y
n5JTQwjmN5kDMPZfe/L3K+PtkwTXWG28abWtejvIra6V9GRxN0BQ43KO9hv2kn+Y
kfYGu0TIbwmmw8PIcmTdl4RMqRzn5CHgfF+hB7i4LVk5xn/pNCA933CSyvpgvfjx
RPKiepbavZM6f4UlOjOuGH+1YE+jroZqQ5uVHz6/SF68dWAovQ5BxFB8Fqv6qdqG
gYO3ofvYys+/tle85E16CilU/XcMiiQFopDtRSCJb9BI7Pq9ZlR4rZKJTE2fQAa2
FyeClJTPmYoG9Y0X9cJf8bvAoL1AtCTvL7NbUDpoPq2MhVaEmmuPJ4Vgm8k1/7Oj
rI5K2mmhfOo2n7hWYyJPtYAxJoyTv+oZ6Wg8Qewzx2ZRsGZhdg0O3RZJo1Ssx6Ow
X4w9nX6kcGTebFnYKVhXcj4nsqRv7IXI/9QKiu4VpFgD8dZwiY5wBcIHvcbBDVAH
lCWngbmD3E+w/2p1adXAI/ZX43rESqOCjHGaXvw9xVSGF2x0gi3VAUnDHS33Drli
d90rpR/bltDcVlCfmFpxX/BYwUXbdO/pqNWlhS/YqYKru4qwIyVH6iqrM6iZWL/W
2s2Gj1xWstLgYSAemTyUB/AepaDWHTW/BL8Iidb3CcwVrpU58zgyjZTsYtHJ+uTB
uTe3bPOwbKQsUbxvqivcuk/6/6AJW3AIOb9zDXj3JLZnIHLZOQX7fOyGIGA97ZoK
I022JcpwnDlsJPASaaHEyPZgS7aTDHQfvtOwXfvD8jVrhtDJQ7tt5p9dZpxqwzr/
83ZtTCLs/WK5uSWoJ7mif1ktE8fb4SDBnrEeBA0Zj1Hm80ktdernh4ZjiHHWevnD
fx3yPa47E1QzyblnqZr7zYaRkR5Y2DOW9uVkii1Z6BhZ6f0u/Skv8MEUDnvILZao
kwZiYlWty3QPekiYJAAYDcHx4q8oxWOOOT7xyAvM1/QEw61d1IINqUBYFXwom/0c
G3a8QJ7vYR0yVhled8kwEz3fUcb8sYUhm4BQ1yG01A9muqNDjPXiqfZdGt7CE2+p
RBJt/rpkMdtDdTioaptH2rUoFYtwdtvLZ5zqXbBvDM9gByGNjopuHDRmtXawly1a
u2rWQuPEHSjlT2N5BIx8YfpZTxP+J+1i02PsrL3A64njV6C4B18C5QdDAv7CBfxz
FXD/bGwY1vFEg+SGyaBOqFKP2jx9KdESfubD5jYgE6WvE2cM4COe3Or9Oo3pCp1m
NGVugEbcm8PfsoRXwKpPEXL9BHjnDTumCYRc3yAH8611uYJQaoNWlDoPFt5Lsg6j
7BD+hoZFGOOzcmjWbvSMEBMRubiAjfKfGOfqu5gE2aZ8q0MrqKvh+BIhPmDYHTEK
ITzSAkLjw10H4TxxzXs1TuAoW4sErNdJ6yrKOsde/2wpXVTVyoDpdvTzplG3nUYR
955FWmmHC8bNF12cuZEsmfqHAtnRkNKivEotnAoeZqkMNumztA28EoONerhD++TI
FKh/VAMVKmU5ZYSIXAT4xch//1vPTiD7kgYHEW7iCwBO57IQlBgs2+YYDoW/73IZ
BVztVRxJl2AfTEjtqYZ1eOAGZSLJgRjVjiX59EeDyPWh4SQKtvuh8pQqpyEY/51N
tOdSY0409UbIq0/uzvJZqQu4Axcb59JqlpxD3ji6XC3K3Yrodvr+jY+CHouwxDGo
gIX0YUzSYlhg7p4OQ8qV+AQXSVEImkMzy8tsrT61+RcocICZtq+aktGK5MfTneb3
IFjiQXd/tCpGqc25iP4EYcxpd9kTO4pmhsMTXWpJ6L2nzUzysmneaaHMtqAEbKZt
QVCi73kbDQwANTa0kw+HNMbQ+T1rgxNFbSesPrlwGNJ5WcTyHxj1+3F57f+qvhQa
l/VMyfkSCfOr99qLZvrDG/Me9eHNQB/XZQ3+Ivl/TS+FXwUZ8rpkv5XIc/Oo0xx0
O/tPnOxuUgWnaXBlt+qmySH1VHeQejF0bWYXjHWbVoVLgrUzrJ636Ugj/ph69/c2
Pa3AUWMxkPfx1TrFOalP1ePiiOcsqwcJvYBDAOGdAztoUs09HXbjEuqMm7Xw0m6j
CIeQ884Ed3M+us7kcSJtNPfFvCE2pXe6Qv5pLuJhoyC45gb3IZ/p0fmXrDM/6SHO
KVaIT7j3KuOdH56QoghV2ezdHdkRufPPNXsAy3OmPNItgENvjLhSeAV17zvP4vcb
T5sMOHb4+ahKpvDE10ThZZ90QQbHf2pE3PhqJilL1r+FqX3j2ZV8dlc/Lc5r14Gb
KFqZFQbMPwr6uUkvA5YAmZsDl04w+rQ6QyN6znfNFDE3Ew4iEOXTKU+kcaCdIs0k
tizsTjKrQcsqsEYh4jZ07r/DFz3HKXOP7tmhpAFGP2rHTJOcGJGiHuMWsdpzG6QO
Uncz/wg2iPGNxce18Cut/5tNKFvI8QAq2VNx7zZOvepKJh+bZo5MHmau0XURtRKT
mxx3+fImK0kEsL1WdwRQayLFnt3OPLpdbobW8O36xMod8z0IdOjz9VSt7cJtowT8
KzmtUo2Fm6jMIsQR9ZfXgFvOk8x27bKVW/BRqpFsKcLMhUWdEThp+bXYKMQ6Sv/v
mAuzTa3DlVoIoNSDbZvyYz8A+IGASusdFk7XderfO/2FfT2ZUD+QroyVFZweSr6A
zd7bZ5JoJH8fE4DG61p9+b3L35M/wDBEpXtYfTB/RWNfu8nc4iys+uYdRLvGRHyU
OkDIaUhymX+0Bd+Bc3BU6Eb+Ab8M9QGpTkiHwxiVgnk6xe6elAUuu/PdDiK3PrSz
OAmuDWYI/dPrk4ZwJjAsjVNEipaEbXUoCEvWMxKg3n3WHwy/U+Bx5Dah1O4dEfcK
+nYP0VCZXA2eBRdKju05gq+GmRVJCEzvQxq7jUlsmJ4bwlt3+KHxC4VEg02XJSMN
RzwrfS827idynxUPuJnxapHQcCsljXtT9sa6Zs/N5j2Y9Ay5POw8iy8cQ5xXYc9d
UuVhFMNf5AYfv3uUpR/ynT6RNSsLmTzBbCLPgqtYMuYCQT+Xti7bR47qfVgtCYKZ
yVbJE5gJdZGnZtx7M5mVXZzQ5ezW/7wZDQKBax3yfA3QxkQC/9mORbzH9Tv80Sp9
q1QwybUtJg6CtTrKPS9XoJvuK0cgGzxgeS7SIlkfrYCys+4QrDp3Ubqf+84/vOYV
MFtL70j4pNNG5SsP80ljQ/iR1wfHP7wsBWPujvvH4ELxspe2eiOjwe59uGCKMzyC
xnKGJCfwXwNCJMbMKv6kRPSrZCX/3si1UyHiqhiJ48ETn7MLfrZ3SIxk9nVrU9Wz
r0aDIXNFOkyl6/5qVz0IVx9PxKFT0rJeWvyhUO6RjaOtoa7ZffuPYLGXaeGJh9CS
dqYK7MNBm35GWlBNH0o1LE9Fc+CY+DGFApxd1uWVvxAQSuQakx8Vtpl8R2e53n9q
6ztwniXrK95FYq4uCMCFzMsCeOF+x8qPUyzTyQA17G64P3G+1vvAgtI6EtvU37QQ
7fX61BllRDg+635cTgVso6Pd98hETLlmHNXi1FBjyFDIC57Jv+oPzLjdwji02Wnh
S90h+a6QX6jwiGF8fT1Uqk3hWD1ket3czDPbCkDakUI3SGzgf4lZXSilojf3s3JG
e56ZuOZcsTWFHdHsB8+hwGDBXjnWAfY9NJdzNqbDRFlFlggsBo4WRAVOIhyX0h7h
uc50QLAd4OyJts6ieBhh3j6ZGZrS6JYCe/M6jlP3ge7R+k+WypqYoLqq0UGOVQlZ
KQwu2HhAdVlvDrNpIawU06WKyU9ckj5vpY3wYLoEDgo9Mgt0GgTJUjseeRP0WkK6
67NLBqlldLm7mmAOLwHTQrfcijJTw9FJVgIYZMH5vvR2hQETyFO0POhK6B06MNyK
c9niB0VY02tvsAwVfyBAMO5w86XMwjg5fPkV797jsbgghsBcYz7ScaoICFTWbVpW
pTJvtCNaIXDgedD4BK4n1Z0TTwJsuS0/KchFNx3i04YPt1WLmWb2SyVtigV7V9N+
6ITOrR8u4AO8GQjd1lccL9CWu+u0m6dceSPo5A3VlE9STJYtKtAdxXFvlkmZsfYd
n0yT7WdjYB7AeFqscBBKJhjW/g3q6aiUXsLjp22YRat/ux2IURCoYGKH7NvYLI+2
BIkjyvleXNa6ux99k7qWXAjlSozMUH7hinROVnRTWIDQWMQrhsp92ZeFDMCJnunq
m3DBZg8xy9LqfLj3FKQEoP/g7wdP+GLyZEK0onKl1+ZFHkT/6Q/rJVO5UhUxVIXP
InkHJ2nT7JgWRXhcJ02bvD6fOaItUvu/o1UxK+t7GKm1ECjmgLfS8CvUPbb0sAP4
f5NgAulRWYpXuDl40TuizZR1Y3Y/ZbSeasqhHG4AknA9p4neFjE1IcOag8ST87yk
23+2GcYeoU34X+dDXahK0ScJqrSf3D8BV9w975V21/U9YDikNUDNrPIN3zvlY7U2
xwDE2UmkDfd91cxidEflqwlZMD/U75FzEVSLQyjiXO6OIvXfJRz+G9ntj7JJ3pSD
SaWIE6fz+EBnODkDJASxnlxsKFw9KpnA/4Y3/J7Yxkxf+FCF4C0OrMXzNExyCo80
GiorYK3Xz9Evc8bmtUNEn3rcralYeXTMoPAV+cJwb0BF/KDEnuaWhS9YymUtrIsh
g7OKmNWrYp1s7dkl3a9Si2JIqodfPf1o17YW6czsvrw8P5Tk38Ew/WLdPAJiL2NB
1Acc914EQ49LjzsML4P6zg+5HkeTnywfQ4KWrhQQeMyGdEs26C9CTtmxVwzadIM4
iHwmlgc5MVp/90fbgZU4Ow9uXvQnJqoKtl5JZh2Rc/16R/SAy3ncMKTSYzi9zBKH
QjZ/NWvwuZ6+9Y/rJgoGp3ZRTQhsNHA9NwnIbjE/s7GCxf40WBnW5H0IfjE7pUei
oUB2XoQlRSBhT6Mm12sABDTJcLHd6clWq5CxG8TxEtMsIn0dZSyBJ0ctJ1r631xK
yGbQu0mgpSstf8EjTh9uNUqSsNwoOQeingakZ7DhqKZ/5N1UmYQPuFSrwmzHwIxQ
o8X5bZ9CNndlm+qsvWfwQ2Uq39wkzDo4xq74HkdX+gH983Cu9eQrWYsvdSa6g2RZ
XH90Hpqdil9+wdYOPO1SbtOpDNqcqNKlMqfUVdhAwb4xAFmd6NJDvpLf2eFBSrus
HbN035kqGNMXOQXIa8Ge7NX9aEWZoNkuamzkHHa23qxauuwzQdSw+VC+K9si0An4
BRwcwmjxmFkLisQfKWhOB7DhjcYPBBIfTV6YIsFh0CcC4l1dlZMO6wURWU92SZl8
M0TZarPiN8iZdJYiaYYgx2flSWz3qeZ5AhgeQbkbUZx8YDSY/KNOgtnnd5OgjTea
IPCebNJYvUtlmgABSG9bt9/v+o5KNXD8MlzU60zCgo2kLfFw4sm2AE+cWDZKVitU
+cjILSKeN4rr/u5a/Le4CkucS35k6FDV7Pz41/fLnyHB1ssWa3qvH3GZbEyLWF6o
SlLEOKzJi0VhnuVy1fu8sljGVXCwqajBIjii+KYslFRSrmXmzygd5eYkpO0dPHHD
lkCVPpDEyd19WmqOMabl+oz5anmm2Ke0pRCAo2MCJblIYCcaaAt+4bC8LJm4xL/t
EtLcBaR6HfJvORjzzRHppPG8Q/namU+eQ1EdLaEA0FeURj9YkmoV8RdotVsKEq7e
EjIW3YH8/+MqX7HXU/JoBUE88OxMi6v/+8yKW7C4By92I1vaoVrtNgUNYJ15uvkD
4Z8QGZ7fZ2lOZTIq+NdPD9UYztVgQFj2daHsQ7fO0YtVd60c/iTMu4e4Bzo7qmaq
I1jFBlYaQLmf2+V2RWLcu041itMZUaYRPLxw3ukSLDJmNZ68PkLjcXJuC5HZ6LSt
Rjhy8kMlErfMvm5HbJT+q27I33BimofI1TF6+2EvXRC8Umnq6Bld2hOx6O8sgJT/
ldJ4c+gDSLE6c7BUAfl1n0OflYIToW7pTHyui/4fnJQaoz3v3JvSegZSdzpOn+xp
kQASNwGTMeA+JldPuKkGyIYyS9iSz+4IkBpaSvurgOfsBdM4pafx1IlYAeM5qWyE
dRYGvZ7pUJwihyj49yp+Jehpy55yx97DM0qIk/11yc4xkJR3Ei9a4N7p/Fwinkz5
8DMzJKB9OIqu7VdyUKhV+3stpFQZHXogJ7Mj04NMvvObtAGu+jOd72wq0uNZTt61
KRM7p8n4KV37EuCHFP04rbkeb3LtGoaX/y4x7n5cIbTCdjBxE4S7LkCNPYxuQObZ
EsL2d4AgBuhYIFh9iB4FYdxEG/vZbQ36sq2FwTF1OM5C8bTt8eUVSlyjPXjl08OC
UPMseb+sNGqHCA0F/iWGhwR2yaVHUTvC+6UGA08cxhQkPO4wnClC7+zmmFK87pFV
IcrfMyk9QaVRPzJ970siMxb5JNXxbPK8z4LwwZAv8qUlfJj5mwCiqsWiHr5N7Y+e
80Mhf3k3lcYQDE/SZ9yQNZYPGnedqpZnBFdZwdOHt+DqFcANvE2HHXyev6j6sOsQ
W3rBfDbGx4lL/YgSrAPKi+o0EkyUraCGVz6s4S+wXlSZuxkCUvqWly6EUDgeLERZ
HWihwAgKb9MA5lRjgDjv2Txsm5+Qikl8WxS21BzU/YXNo+n8O/xenKDr5k4UAvKQ
097XJHj1eU1JodGU/rTwmKrkUSzDMs2sqtQKmAjm9uxPS/uMUqZmv6uMo6dpuPAG
m1vx/yjSDwjTGk577aMPzOYFd4wB57Z2865Pvd0iyU0RUOmGAsBfWu+rpy0tHCrD
1H7HwyAq1c2Z4U+r+OH6aMZm6WwHNxdxaRySrge4M+JrsoiCxOEtE11INPokDHm3
KC8z6XMxoOhkllYjuAjJWxfp8wxa8667y8MVeyRYAGPy/y9NtQ49+0Q7JcWBFUd2
Y2y0Rn7WA7k/JWdmhDIQHUK9JEnCr88fzXBJHwZNHOBUbnrXY98z/ByDuJsyYt50
HT6PW7xfrfao1hXnqj3DoLg4MJpdEaoGWZ5CyJZs3zXiC9m9gQ3lqDj967Qmu+MH
TIzVk0aRVva4IgVzsO0ScboFOF8NnRIzWp4f5DyovwQgef2Cl7OGYwAzRiJQEGxq
n5mD7DdR/qL5R0N7gNJo+3yqkW0cUkPZA1qXZbr1NgliFiHZJedcMzr05EqaSI4M
bOZ5/V0lV0qEX7THLFEadz7fym5Mkf2eB+AoAwtvLKnGfrmurcWCSMj/9HC7XfX2
zHneFWBw1NRqYT4ic5EJzwhKO7mEAViEelv9q5xbIEE7rAiiYxsCtl2oy1X1xsYl
1s/Ag+Do5w4HgZjRKdVN/smSp+MISaHLAm3sPR+VCNGLiOZQLQztAY7a3GBL8PEq
x8qMiJLbb/KKJA376reG4PZat5qL8bKa8anmVLHFTRnPaJGOCQ0CRmwI/2k5j4QI
MLmcZdfqm4kP6hrF8t+VVMc7unAQIQYTVxfUoiIrwgNf8i5gCN+I+l+Oie83cIyX
0BD7pxfz7agDJyz8dktZsT3SvHWxo+THYFtpYNVv0tJaQMoO2FUNZqaazz54xvN7
l1AayRn6sveFGXx8tnoxhUjAS25hFM9CNJoWTMAUF8+TDI+JJDsrfPHzQ8qcIxut
VIS6gppZLNnN5X98Mt5BSZEv3agNSvSLqKGSHioA8aCt/D9WzryyRReXDTFNb9sR
R5qTJjqtuM8/ar5Ptlp+F50I8XY3TIVBP7hgRIrAMU+SZIr9qY92X2eeGYJUDhQe
YtJnLQmGMqnDt1ea8xBc3cHkTxcTWWd5myy8tlY4FM0dCmylORG1dcbdN4eLuVbj
f9Fd78klu2tc0KMejm6tyFAkHF4r+Xm87SgI9Ebu250vUNi03/xZChvbNzHCaJ3E
PkSxPkz7p7W+miNWSYcTeudjlbIi2YE8vPy5p8K56yq7rFcMSxI4VhKDziQytO1z
mqyTz92bmGy5LGqQBbQ8mY1JCGsRIYFKioCm//B06JcI6O0JYttYZn2zUC9ArEdI
PNLi1QX/Zt68M3Lu7OBdTURokzMFevnCqR+zwuBiuHERefedFi9z8MFRz3I+9S9q
Uw1ONrAabfsdfYI9hywxuxmYo2HwS6mC7ogFmRfxyonVNJuMMec1ORvAjSKH6dQ5
MDBz/7y+9Wuv90upqsAYvy7jH1qqfKJVTJFhtq+ysBULIndX2vEkNTnPKPBxVO0A
7ThyH7kgo9h2noCccZWjt7Ny/J6tUJXQ2L1w+FyxoGo8HmCbi190Q5M86G1QAycC
i/uFOCW9TFd5Y13g8469EJgzDWCHTuOUOzxK+jjoduAx3SlFi0ElU0Dj68XZxI9A
3dBnog61cYGW/NTO+EETgtcvDIW3PUv5Dk+oX40EhDXlYZDs+haMKJad0Of2L6Pm
9zRbhZpN+eIuQ05XxuH8L+p1dZ1v21eVqjNoaU7zdsBOPlw3SZlv1w+q47bJmcGS
Kpx0iwMOyUf3EOf36++/dGlwhr6m7qVB3P3U6EjH2ALpwHe4Y2Hq5DgHZ9cozlDO
oPP43xD1KxyOH1Y0ftcMGMJsMS1Nxk8KH9zc9+TkmjJZNugCI3MKWTE7AznYNYqL
pcczmJhDz07W/PF4f7F6GH04q1YG1KD9Zg6eYhynfmu1cEfaL/tajGEeW24nPLxD
HsE4cdQrZxAhK4+VIzBLfpZFKtnVTYFpS4yBpXcpFpPBIWUmlMZrlsP4gXV63cvH
sYMM9OdSahJlMeaajQZmMbRGYQYL3D40SC/EOS3VWeSVx0CeB0zgm6ICRMmz+YUP
U75IntpCUlN7WBZcuDNNC11dWqfLan8OxBsl86h/eVy4poHivLOLezn/f1r/LgXE
8Ed3dyPSyar39g+zJdtvXlC7dvx8NR0UyW3AUVDSRWP4d3Xt6NsuSCe7EioC4r/i
EJ9joa+ddme4QG6J+fJx7hDuFn1xWk+8ETCrIqmg8jFRtnU5UpfILpC6v0nL+XVa
Po/Tcj8+e+EQ8QoY89sAOTyZ2QMNVOm3HV8Kj4SW6brLrtDZx1AUOfN9ce2IL9/6
L1HrUMrWMH2AOgghTLg2gJ0My3U9e65M0oot7wsJ8vavOZjXarXttJ5JFUltRstj
NS0IwSkL0YgzoonMNxqLgu3UcZsvNzNF+Y2+K6fkio7RR+GKu7KbXZfowe/yBU/n
iIIUl0D5pKSiwVv2MrqN/Vv0RHL4IOq1kl1DqouFR6spELW0kIk09aKJEy55YMnA
EOE1Hi33k/WZ09Lykrvpetd/QoU1ivfmj9dPHQ6k5pmW5elGGbM/AfeDfZW7Ipcp
qoeetuj/c7KgDso8ZV3KhYZo6esfI8cj8fNI/vnq6bTJn9IAVhcEp8CD0diT6lTX
VgQ1juTibyiqKmciu/cnLJLTR8kP6fNxF/mkYRbal82wYpODp+1AmX6PzXa2eNWM
YkwthCjMLpQYRaG+mrnR/9vnHEuECmr6V+JVDYSdqXolCfpUDo0u12Xn3bSMGi+m
CNI2hLVFhgTLBpCVZvdjobraul4HXHQNmf4F8Srez6BpXD+DkxxWN1wJEZjrGpYk
jl8XaTDldJoqtDIYX8nKOPKlhVvehWkBB3ewJ1fu7eJx1Yyi9yus3DxUfxUnCahg
Lvr86YlxIwyE+dijq32eV+bwJ2NV/y2jAeuVWXiPvZaCsJ4fh7yhUzxnSUbHm5VP
VqUW8ogtwD6DCnaRu16VLUlLUu6HZGr6S+/m27RqnWR4s134QwkPgPFY47AmqYAF
ucMvMNwNuePcqXTDG6pznFAH/HnYF5Bw3+n2V0jTEaXy3KOTbZFxYLDOj2rUJpOd
AbbGwPfxnpPzWbTNmkBpdr/Ohdx16lsRDyp4wDNTg5v4s4pGFLd8RY3m7GFP+X8y
FqtT8WbmfLT7//i29AJED599d07V1fb2lVcim/49ghuy+Ch+7UCNVl6Y/ue2f83v
6FLyf375EgSHz4GQ6oBWfxHVHfGrTrsjABVkI8JzUCusinWZu5z6Y3SZLH7K9w8b
oHDEryw5y4/A3vkxecXSU0tLGelRGloY5Bj5c3SnVo2bUg65pe+eMROvwZ6EDFFb
zyjRdhT4oUSd33dmkEkD0UTdOsUAIJMkLfCiNUurPSwuPlIwUlSgIgWTcCdAhIlv
Brvsg9y6e+1T3D8CWEaL0kGhmcI93MmALJ/4x+3JjVdfNqB7C9Zl186v0eJeUoMh
IT4JNnEPk7nIweeY0qfjg4v83HAn/4lGpIIUox5myXuSEumkXslfIrwhASfTicM0
kLrmpiH8RHHNM81zBVuvrKc/watB7Bg/Yrjvwe/mlqbK1faRlzEhKtQmeeW7UlS+
1Bxh6GarAArVdyemlWjao34qdYtti85Jj2Ct+kNkoLNE0ikcH2F1+fTOsquGo8Hu
Ws2bAWNzYAD7N2Cs7mYvmkEgu3AxmqVkvz9aHvZeA5U1XbLzKSTIdTLpLebPx+PJ
+HFU6Va0DsXxcHBN1n9NOnfmOEbVZ6GtsjzvJ8b8nqJkbzQkQsUzwVJRg0MTddM0
34bb3dBYE8uS5GB0RhChWSO82OOx5PjGF1tVnhvjz9C4pgxlYd+hiHSJH2HjUX24
+kiC9mjJJwNWg1QLeHoyeU8ekx0+Kk+9LO5GkGsf6mNbxkCHss1/iU80ozT1sb0p
7kmvF9hEWc3PjthyeIxQWQSY8DZXXM7O48yAVRXJVbi2g2fWuvkMiht/Ac1TOvtp
RjjyyB1nnwW0rDJXSRzDmvNmjhwibOS93w1NCzYggGw2yCJoatdZMFc0ZnP4H10p
tPuUTB1y5uSOArzViuXAzYTZ3iEs6wxVGadkO2qjEU+LX3timMvpLR9apMiFgOaD
rpavPpi+4iVPBq+aVHtjf1d1yNCxzsZuDoZYmEedv+kW6+13JitD8yeVN3YO8ki8
BAjt22w8vGRpGmiBsSvUFjeUOsaEQoCCswcgwAiBIM+o1aRh3RAIX/Qvv3SJoJwN
qZBdgJPsJRAo82qtw2fF1QK8GieacikrAjuHYtWOBX+C+LllDdQYZvpau8nvhNYv
Hzh3SDXSULrnJm46R+8FZu8j2yVoQNUYrQWlAdT55UpRrHtfGU/bO+VaJbFUvreV
XJrPhJKU9fw0ISLwpal8OzvTjoHc1b2oOcRJUrghj4N7ezDx2Sstsw4QKwXsuGXu
phJzs+v2wqfy9rgnQYiMa5S0Yzsfg8g7a0R5iv5Iv2/eWVjopm6MG+0ap8iDkxOc
lwEiZTx7WdEVUjnCpT9Z5E5/BvjwhnT5nuEVTpmU/Hn0tmQCnhRG+zlf5fLfxVlO
J/y7QK0+NBnulcH3Mk1VyY43QZTJ6qRI9hpaOX57kd+1oSCZXH3Ceis6AYa0i5XO
0gJCi8gYqOOmk8+ysyUjtY5+j0ZcCyjBhl01wgTDCUNI3CvTSLIog7Ln6/GzTqnH
Gjn7pnOhFzfg+DXjoOjPzTW9RVbEPw1+nLvyc8UI6qhgiFBt57c8XbLPKDAmXea6
o/BHC6bZFJKEI5epsDL7x2tItv3wj+EtQuBogGv5eGKLJjNNRgkQnFA+E6a/mP6S
y9Nd+0v4Z2aLF/6aaMwnjSNIoHwteUAsRfrn1ue9LqXRk4osjNh9mcwbnjLnZ+tK
4QrXKKWDu13JMBSsJtPVgCJTiZwTaGgaEPQmVwTmaM3nBZKFAsWuZ2GX59o+cFO2
u246JlEgwJ58JjWKeUIIcmsBYXzlpnPm3viz7yS/rZ8TeWbqh3PtHxq2piBsT8MJ
SH0BwVyMxWXPUxdYEUd+pJkSiwYRJ89h1V7Fl0vCgL/WtIOHe9uWjKOvG/7OjFkZ
WKODv+ypX3DZkfYC4j9vHDlyctAUYwJUNAPQfFYRNJ4BUm56nhVNRj9Ttwc51IGX
uvcmdznbL+dj3h4IAgQM1Cr7uJq5HBSiKkAIa4q0vv7uCHcKObojS1JaNyv5EvJo
30exJP8RNw+L0s698+lODZA6AY6P6upwzeZmgR09up1ST2pI2LgnV5218LagkVEC
AYkdNaHxrmgwQ8Zpz0QtrxJ1yZwFdwoHsx95M+B2DjdyYDWKIOIhd1RqGByaTxw5
s1oBiR+/T7eeNfZtwGYF6o/ZDN8AQvh01nEZjozVtBDuGtLihKOUBKwJwEXCAHp5
3wjuuDGty9DlbQ4GF8x8gfSBAzs5OnaDuVOojTliCJm6h9BmN6+n+/FvOdpYYrIn
9Y7lSLaAX/3JskN0EuluEYARxEFdSQW8Xp0E4jhcNOAKUxnfMWKTqh9zUAbKxNlJ
8flCLvp7inMrw/WT0rPHMC5lXLpJCfMnxwFOIKvcokI7JxlZ67A3OTE1ypiiC9rt
beXRcIa9cLklFe6oDYQbMN2fRj9+5QIt4B+FWtqIHuWsEPh0/EhcXvHxhuh4FYrm
OSd3Wxo+nDeRzRlqAUvfSrNF9HZrcbtO+Y8Z42Ht9OhGdP5OdikecCsv8J8xp4ni
XUH9RWE9nW1mK7nwgSzyyqrFk7XsSUAXzmmTl+kkQSktfLuVuX3sEKIssP+6NFpB
dkbrlw8+hheefnbfxnYccO00p3g2sd+VFbz0y8Eic0idCLwkIjsX5TV4Rlfco7eR
kaXZ+n74rutMDhyT3qNqt2AC8XdauFRf+N/npVRWFAXz7Xj6sKAu1ayAFnE3U+C1
caopmhxwqz3vjv76pDYDoy+jeDiUjeLOVl6V84tJ5uMKFh6PknvssMvGlOsQ3uP4
ds6GrwD2nTFqYp0v+iE+7gBibP1AraULkfKxI5A/RcBZMhadmuwmqgmJGbuzhahH
zl1H0oLTSvlQLa1tujcbDlaAbhYG95XSBkplyBdqU7qsvBxpQDrHsq6rKLxQUjrl
nfSA3is80yFWKDEggGzD6LKa1h8BD3p0WfA63a+EV3I47jqQuC9CFMFE/gpeLjHi
GOpjjj6Ri7zN6JaGB6rfqeuYI/W1Z2v1em47bOqd59VJWaJCNDuDJ5OQKdkmaTpU
MVkoaVenkcZJmy4L1VNcY7zp3t2hWpt6xpxaroLj/zVAlaP9pgOlSVy5pkV/Fnk/
pcQJAeFYlUmWm/TKqW2kgfWwauk7BEJIwulDPM+UUT0fyy5C6rEFHpNoCYjgYX8w
IzQlShlmcTH1d25QBPYiaqDQn3V+7Cs9vpgJ/5wbfQ8qpEMp4xAmrK88xqBTUUVf
QVsRl2xMtetZTmx7VmlDbGTXgxLv0aTK3VYKhX6k5plZoRwn61ZtQ8fAr6vIC6dj
Mzp2X0rJFkmHHFvv9FV9OIyN4YLCuM3ZerMIXT70acfymGzHlW4uMvAye759G3yD
jRWxISUXrixtpCqsMyATaX5YjcfeyAQPIkC6clDRaM5RATp6ogIQybIcHp1axiaz
DV6SUUd55PyrHTa5tAvexAR0JqizfmhtWjqrZDmJ7qkHhoPii/UwH3Y5XKfObpFC
4qEtxdGfSrGngbu6gqyaFlwnNTq+sn6fjchSmIdvpaxuv9IXieN9q/3Lc4IrqmmK
NMCYcneNWQCN8N6FAkNsMygDxsTN2Y1sJT0lgv+2P92dpA+gEgIV45DezqkZngki
gtT9mnx4h2Rzqh6dsM8My6kPljXJnH3g8Vn1cdvTFm+uPviWA/rrY/sf5Guprzds
dW/+sTCl0UGfwbi7572PfdB7KDfdEqeawXMsvHtSePZd9I4L45tjm+bCVegkzKGI
2I+yXwxgMCcwvHjQT/BlMuR8u+u4fdTlyS15HP/CHaBamRAW3SYVfGTriEynBsBZ
qyvwgchI0HZkUroKuBCbXj5TLjPthRgoIgnVvW0HU3tMUSGGpjp/4YYsIOOx50MA
xiXEPrf6Gy/ev3i8kIuAdskJhLktvrH5BcVFN1hpOXHAuMS/SEtNncq7rm/m7CtF
PTANZPzGT0UNUF5I0BA05Bzw/FXX7RRCJWWErCsCYos0D5EHQtvuU5Dnl5ZwqIzE
Isy4OU4W/QCADmGBbLGK2FBp0WmlIrVCHOkhoOqqYMHg1jpzeeVlD1IvbVMOXp+E
Oe0r/u0037J77S90tAL4x8OlCbwFZLCglUOCH3Qr9UFla9bnHsrDMVmPNyOxY45L
yxVt6Hu3lzmEBK6GSTNLv5vQIKjEWLgP3F35VMZqj8OJz1P3ztenGsw6ieXRe0cD
`pragma protect end_protected
