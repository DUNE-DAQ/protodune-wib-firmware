// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n9wE8GLn9OBMLfCmDGCMgbx+lKRHPuDaGwAdpZRMUhVu/CsvTH+Dipty2hwJEfCD
8HW59IHNpzf/NHRiiL5St+zWjbSr+MllHn4yfceXB8dTBkCihzWpsA9rCdVlmkhD
IjiYfwsObtP0054TG1ZBzyfNdZ7I3xxwZia6R92i8L0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10000)
jvhm8UIdSKfFjIKDizg19vrAGw3kBf1bTR3fh8LiDgQbC4BzDHKxAJowSU9+c8xe
Z2z1YcFiuD4SM0RSoSKn0xuoXeznsEiOnvJwsyvJAGghc4KLC+5J79A6nGzbnqJ/
koZte8k4UxzOK3aLCB8mX1+cJ8ZpCnnAKKYkAsUWhYbp/qUuwOivOYzGon3OllTg
Lj0merpo2IzzXOLBwo/cDVQG/hEI9GY6c+onI/SNuXgcfrkFvSfazCs1yi4tv2fU
VMaEbq+N6y5eWskGdGIzB30IND7liVJksNfprirZMTM33+1ZCWMd6AnQXZxv+SQC
Ndk+LFv99Kbm/M0bQtttRDd0wMaHr65mi9/LTXCcqKw2ucNjmzm89XUeubrKbzbJ
LYtcmw6DVNL1kOzhcPN1sycv6hsfYx1RxVOqn2u0sNd7hYbp9OcS96nlmPL5StzD
iYFv2F1KTlG1SWXzYElRwOzHYwleB7AvTVcwEEgysjJoxcOmkgizZgVEFsUBtCP6
/jBupkRAjoFi3vK6YFZmuPj/IoCOSKlPKitl9QqnRTudekiKWStFlbFRmgUbTQL4
gEfWu0dU9mjxsifw/lIhTrQ5cqjkedAWqt3zdmRcT69ujW7nKZS2vmVExiGZUTsw
0QqMGL1xarASxMeIpDbuMDCIv7N8JsBz9fYuU+pD2RGRHCBd1+yXsLmqX+bj84pI
fZ05ovN9ZeJatSg72p1yBSNIJYP3P/Srez87qOkIZcurjmq1BPZEQUItnegi+t7t
1ok5YJ24ztnrzVZuGrzfpVI1cEnn633As/C2OiD6db7shgLd2mcUS+MpnppVPwZl
hrr4M9Opf86KvIR3dTExrdvehc62inlhVKVUx9q2JS1Y3z3d44tvaUfJ+WpQPkBe
48SpadZ8bzCIWCZxHIeS2FUTKaMXwYMZx7s6/kgKm97K8cM3/Y8vfHEK1tmE4XKr
oNP6jfu4Y0MRY3AgVA9bZvbcabz551Yk++OkHNfJ2qOPDmrSZeo1Zp3Ec6VTsEfH
j5s0Ni66Ema89xegJXB6pFjRsDkO9MUqRRzBF5pYkLd2Xh84ru3lzbMlsCbsX7qA
6ol8/QFvMGY2Dt/Auaa4JYZG2axSWWzH5iBl105CDQ6jdUVBU02O+ycZdHkQLU2H
W43NXUP46HU3014cRT43VQzDtZnmQ9zGWe3wQxol76JFyadjLqA2drKyOb3bjg6h
GcG+0FXh79hdbL49M8ifACAT1rfpzsj7oj4kjjHAqYtAjnnoeSZTADOLjGyAElSU
Pm9SyaNYlxESE06RqCgqmhKmjCx6+4BWx21PIYtguerWNRO0a6pOQN8p1N9aXvmq
pKzjW43K8dJq/S9CllzW69pV98A3en0a8izBCx1Pw3qLeJLZli7SlDUFdyQcjgL+
bN7w2BVTJrWW5G57M6AmFA/1ANT4aZPGsWKSKPFDIfznXgNruS8h3gXI3MhwixFd
DWuOO3zv140LgJcCiaZnSf2H6qNdMjtHd/2QuboJ7L4zzkvuBTCjoNBoZbHtCV/S
eKqFyWY9ntARbzPKtqAXSASV2MFLmpTMwO+Hxr0/nqi9C+KA+WgyGNSMLscLKb6J
lCEAl9TugyM0nVvO2hPPDwmArJVX6ZOhec5j6QqGeDQICvxNQo5B1qZyHBzFwS7I
4d1cNrXB7vtg35g0G7kYQeP92pOjTPwNwTdimwyM4PGb2DxYBBYbK9uLnbBUmiRX
dYzsZcnDsuTx41lU+3b2VM2jle2k9Kvcw8sxFfpcfl6PBDmxPfHVt2YBustonEc1
kIjsKUpNtNDBQ4U22RLLqZ3IwPgKN2tuDws+8cPH/lztsQS8Jyo6ohog7I8+S+U/
KSkhf/HAPAJsa6Y4fuKh2jS0fNUjKOrsR8LvL+PSXIuQ7MZhjucSrGQIqraQErxz
MxxxADuPfzPHcQm5Ekm/iDx4Bn8bfek7Rvr6vcDPIttCO2ix5pqN+joLJEbfTPCM
x6/MrcnsLXxSycewPAuSU2UEjQZrPWcT83SajC/AnejYscx3YExMbGHOxektVsuU
toFOuPlEa0FR4WzSEn1pswmfNPolqNyZCsnvR+Lj4IiotVvqx4o7GJ4EGQaSocT8
BoxNpLTa3JCsiUqQ8/ot5gA2Mjng6c0W9u0f7os7uTPAnsYzXg9L1w83utTS812s
Oz5qmKaI5bgBtB8ZvQZcMHHPD0v6MkOpzIedLYYULSJFgkqhoxQEkKT+6f6ZYnsS
EYX4oxRgx9BGALE5RaU2BmBxmMRgDzNo6G/IE1ZEFTGsaFvh5r1Fe/k9IA73oS5S
Ek9GSPh/B5+Hxl0DCdu1Y8YWcQtKUlWktHz6Ntv6nbvA+2gDUN/XDa9a9DN+FPVm
+cvsXwFt7tnW5m69BOOZ0Utgjr/wvoUIRZEtFnt4Bv90xXPhrCAbDsxUZw4bKfbs
fqtD4GImiL3mt4aVxt1Rwudz9DMGB+qE60PJAxzYkEJvUrzB10KHB+pTh7XWnGEc
kNZNH5Nix7hX5uEx9Y3Ci4QI9jMGtSqJraQRW3SD5uC5WZ9bmaCEXu1hwFEtuW8c
MIzOPGzoFDSdbgpQjXXN/1lVpV7ZPQ3oc4s7MEzpyfGN5O8p+6JbP3Gn8BMZE/BM
csyccqE8P/PWHEVx4xzzApSgZxvolDu2wuA3/jtmh97WRBcXvbZWFavpvh5KvtVG
LOQWxg9YNh2TiLYtr89aJSIo1W0b57p4AnwEv1YNDR7S0SzU5Hva1dqrNxRghNny
A+b9JFbkwh5E82hWT6pzTDmScWIEPMUil+3/UvfYe16ioWHkFLbbxt8sImS+AfGv
sfU4dBncJhv1xi3E/sjmjEeiIFNjxU7YvNgjPenJHp5KPntw3hnsYMB4WVXS2/UF
xLDh8NvvDuHXYkgXI6jOQQtSYTm3Whv45OjxFr+v08p/K0hgsC17XQn8WGIrOXcb
n2n6zcpMuUGkdd9+a2WNKb5WdHskMhhe5CEiBJKS9+G6jHlt7gT2H86Pa1j/ZjyI
Gc5MXlEIK3rYlXSW/pgC7iZ2PLTD4euJSPl0Yq5VBFpYNjtj/vpMr9WgDV3sR9Mc
7e2lRz/mkCOaypQhnM0rUWnn/qAeC5ARQJtebxODpomUC6LLf6n7Q03R9aixNQj+
CADjU+cH+nqXmnx6bHKZrDOqxEYTLInR5yYYlKP+eUQ0enYwOq5bcVOhUI+cBw+h
mKCCpJtckc9oiNY15owXg/mrWH0Hr6EejGeGqkEizljxBsKp7t/nRjcCTUmsQNCX
ICRXiLUj/ByffjHIw2nOnIiWh4XxI5Cn6LZIep2JD4J3nx67wc1GS3pCtW+n8ATO
AbMXxg5XLzwI/1fDv0oeb69OH32UGONnxzQ8/MJKS77SQh3eImQr3Aa9SBZy0dpg
qeJb/Nkt+3iTF3MN7gw+Ifes8z9auv7bJdHn7rBjkLJ4WR57gqfTirondwyJAbcA
1KCNbOOB+/LDoZaXVzsDZr46jCPPbhwrP3IKQd7e2Hel/OG6l8y32+GgZPgiTYLn
9f8uNwJRIZfvnYtuG/Hie5aoYpPQqz8dwW2NdZSzfnVgdRZhVJN0Cb07lav8k3Xe
DGLWgVUWCtgjTo8Jrq6B55o6N0xpuVeosNBFz2N+zrtmIaZ/hKb+CpiQ0EtivAT6
nbSrKTmwSr8Hn8VXqsH0yBFPrVD8M4l2NWPkyOvPpNsEbErE22QFNfNlSi+Djd9Y
zbT5x8lDrzmrQxyUHHRu6L7MsQbjk4peP0oQp55R7SP5z4uUZcy83FfS/k8Ln02O
PEK+epTCC4216g0vDoUi395/fbMVkpwhnPUlxIv+DkMPG/4Y6G6W/5eN713IDjH3
FsqboMjG755O7+C1LBe63MpjDup36ktCZGsXflVMaUp2cgbq7coHX2UjoaEWIn8w
+3pe5A+zyQ+MX7ThB3MxoRFVuBA1f9zX2EEG+VOCEyIL7rMnuG/pDXu/VjEDTXFR
9mh1Lf33w2Cr2wQzXMKe6uO9lwWl+eD4lHtS5yhGukXLMCOnEQpFGJIPDNELdDdL
mrDHlp4xcWDi9qPd+3FiKhaEaJZVJrjYpD8coXp+aDHt/JhtUs+um/c/ehOz8EhG
wyQmWHDhxzEy8GzNJwnFOqA3NL5CRH00yymp5sTwtl1WgYGk1eVBRzcG9hPelnpX
/yskyyBwJNecPqNPkzQ/8ro0NV6RaA3B5lgGklbKJXlV7kw4RDGjmpRVrhSyplj8
VfwEIB7r6+K9FszufxJV3x3jNAdf3mUouT572jZXDTtceaymvwT1aYfz503/JYYk
TFaITkeAdHfz9YzffcJRtqVsv9AZIUcDlLWceonHTVJqib5S/xprnKIy5uVNMK2h
a0Qr0tT+1M9XR/kjHKxU/i0/zthbJUtIqSzgryp8rL/ynes+pPASnprZgI9pRakx
QukpiS9gEGw8cr1QZYvbg7bywK3EvMkpb1wqCyvBIp8UwYGHCunZsQXCelQc2i+i
k+uYo+0mjMoxvTFjqXyED/Au9rnhZ1w54+MfA6VAPESQOht6u8zkfV1bVrMQcXaQ
nG1gG8b1hrBt0GdJaMofnfFaMdAJSM/iKkKZj+CxIodcWRKlHx3EZg20naVl7AI1
1bR6i5kJ9YrEn3Mlu/7sUnVCmXsK3PtX5tDp1BSnPHl3QDfC9nSvKMsOicEgrNMT
cMSrmVjKYoxDE9bkwnE4eQb3TTUUrJ1B4PvE8EizzrfRr41cWzsbJOKvZpmDscXL
ec3Tkhc3r5IdVkMSjxqdc4Cr0e5aIeDwwZs/jevIA489xieqLpvXSmai7ST1X8gS
GS/JDNZoiiIRGvteUwd9wKaiZvq0flN0QPkgt7lVct8vQ9nwYROjXEspuAjyZRdZ
Pw1bGKbOqtNSV2aAMg2OJl2lNHjJ+J19+sGTf5+A6UZCWtRZ8R32ulRS+T1CRVwR
fcDGjWAjoRvPDW1pkRL2EJdV2Ep5KU9QeEA2XzmOguQfyAmnL7O0/5PRpvTBBwwp
uktHHbA12AhcAla3Gyc4wrbqhJedJTt7c9MNRjsb2yPpzH+iRnsfqO1ap0f67Yhh
hIFfuAuJQ0WrR0Bftuztu8WL0B+XlA0zXWsB9IRLY1Tf9FNM2ojjnJd/h3qQJLlz
uajseERmmfvyPyHGz01fJ03jwpYYzxKCLf6znxtKmbu/VDYEhEOT7gV2dUYXh1Cs
XY3PARdLrfLS7fl4y+0Cu1rxo9P6UsMIMXHryS8ZJ26Yc36VzteVtQRw8yBGEsla
Mi5Vhnq/KK3km/Laq4UXktM9qyClpIJ419FXYwtj/rcAo+bTpwBUqaxi4Z7cnAD5
fDle2Ym0AN1cOE/jOO4J1yBMJ9l6d1e3OEYUqszReGBAqoeJ0pN3tcFZ4WI2ZMMq
1AoMa2JmaSGNqp18jqGgWK81ei0eLWU41DruJGkjC0b7CpgnBgE5qDBzQciDIF+V
iMzVLjK1HlnhupcghA847V60oGqzr+FuHbQxmoOC/dlXKBWlUeirrIApkEUM5ga5
nrg/HSnt3j+CKxV6t041brz/nxBYOjMnIesHF86sSB20XibCwEJxaZpxdgzBNu/4
assNhOmaHkg6E33VFrautyAKfn5MkfJdD6IqP87Vz+Qp74SddDzSLlDvTSFgrRyv
cfeQ3hPeMQOmXzwNWzLjtOBJRe+3kPcYTI48Pbl+KY450VJex/iP03Ut6ByiConq
Dkl4y6GaZzmRedO5Lak1/guSdT4w1zs7re7lvVcyiJRWij2Tsi8p15Eavmym8ZjZ
FyVk95RBQq7qpBq6p8LHP4A5AMO7TJcQnA6+b0BVA09KzVsFURL4o92J1Sxrq8pW
itgEB5Ch+vTR4dWRa57xDfw/OdYiCN+/joBICbdT7CteTQRbIyBxqg1re17vVm80
lI/fKKjdYO9hKDuyhP3bioEwtg3nr/45J4Kp8b1RP0Lfwx3xqWGJb21GCcMxJvfS
/bdLpt87qwLYJuVRA69F9PGfWHviQS6QYZW/SzzZcxAsOayrwrXsASYksZdAlm9Y
sBKvbSKvuylxPbqsLBhbHGqFHsmiTtwStyFDZohnyGYI9XZgWwAH5zRlIBQpnK8X
2tGorllqCFHDbL1oSSWNdAIJ6tATMKGccKSXrMrq6imwSkY7ueNf+mgNcOVtDXV1
aewxUjXhZmDu3yR6D4w4zxHNrtaT/pSZHEFadHhNbvumebD9stouLn3T+lkWQhpg
O34RmQcks4CBVlzdCl2CZ3D77WyEznW85exD6ULCaSWLEO1XZu861AIrhMk+Vzkg
kv0m3iegD8XodwqRJLz90WkRqnv9jETl1Lao3aGWw7tp2H55tiJuScJcouSMKNV9
+jGOizfTsVsK5uvHbIS3g1DzieCYFXdd6tVEdv3RvzsQ5T1cw0xlekPHZPdVeCkb
lqP30IpS6EWkyY5NkOA4UsuJOPHK1eJnoA7GT+tnFezZq3yJleFV1/S/rYtueyCF
Ri9rZAaaCvdNSdT+lhc7BJRngd9fUVYa9pRAllWKcyTV4m+ZjYPZiptXbpAr6DA9
mFw6q7I1GTBzxDL/mjAfPaTWAJIIWyUXFdspPkmnkAJIOaPj3UZu3nz+Q7WW6w1H
QNVthb0FHy7r8N8ZN3LUv6zGfUT9spGq0Ez3RwVt/1Gxyx2fMjppuXdHMye5eThP
vIl7iQbqPrOxbMeChp1T/OVKNc54YEOKKNnoMQlBIvTjO+nhynjlp8j0ZsUTHeR2
lTlUt7FlAaauCEcUhMt8HJ3RRErGMdPqBNHyKiWtBUHX1Q1Lr+ev23SRlBy9Dnr0
8Zse1k+ql8jfZtwN3M6ncbTJkAIDIPIeDkJbwPX79oa2TawxLRBZEs8nP2zgIZF2
Wb6Na/VeZ7SdX+abvAz9rkvoxDsNWDSuIOkzDIuLqCZNos5xngXNQ6wZMHbjJk6/
MviGSXs6DnorFefISU+aDk3+jV3vkZEkwfq78cKfOTNKe2CzqvxTQWHrL8xbqB/I
Jgbk8wm85z/+mA3QwQT1T5T01T0pRF7X5lx3UL71rrYc2lOkE7w7XOGmvM8zeO4z
ReOQzI0gx1FmajvpZJGg700rU1MMQ4wgcGa//fvgA5np9HLxmoIGMby+gn0JbEVg
/UXzyxEwW2zfBPprDkOfaO4naRNI/wdAHkh3rAr1QzlOx8+JUPvoUZ5ELLlZbCnI
fFGPdHXT7CCfqdmuoiViCU+T98mOdsyrQzetJIxbjHGa1n10Le5OOX5YoHDUXJoZ
0Aw260aMJfh1Ww7tO67P9p7p3FjxWtL9omVMfm8i6VSY/OUxcf6k5DwxMY/n6cST
jLlu71X1pwaKONqcwMlYRRShZKdtcOl8MnqIgHnZdJLWPLyoSRoSSPMWynVzfAcQ
tQ/o7QRo0dVJgxqUXwKu0BSwm1R/aa4JWbtQhevOa9mEYOjAJP8hoBEgRNOzUCyH
iCquCH1aCdIsvXa9hA4IC3wG8jmTVd7CZ34S4OP8ZWQz6pHfP8CqEDOID8M3KBQa
cx0r6S1e5rTKQzvyjTc41YgBZ4rXC9YuIloHP8CqRpLeUrN0uMyvGjA8XzJHURc2
rYNjzOspe5XvR2CZ5gVI5eo8B+M2kvT3mPX/jZtiKydlATsdKKpJQrLhU93GYWKF
Zx3uNzw06hteY8xHuY7xpPsRE8wq2i+eXyVnoXMA6b7tdRPM5Y4P6CB2LMF0T1E0
vrqbIJX04F0dlj22c0rwoVLDFHRTWZ469j9Hk1Q+JFUi0/R0VTcQJwPiQeM9Y5yq
6fB5unNRBs7slkfKU//khCeCQ2gpG7M9G+ilq+Pxddn0c/IbsvfAaQhCFqkcI/bo
x64xGiKx4fWw7CMG6HvqKEDu/v6b6IMlrTXV3m0f4vLLd3UyHz3LVF7KIYsFJLra
vF0GukU6l/a/tRtNloZg816X190Jlg+kVBO2qya/KjkpbJ3oychsc5ECksjEBvgy
RLGZZOAGcymYUx9qmmVU4HMVzw79hGNXRQxpGZoCzo+Erb3/9SDrouWRmydXLayt
X2wzpDDz0TLakn/fa76fzm0D95kyb2K0/wwbZk4LSXfGRi+OsjwwvB1rIbXipPgm
m0aEJpKDi8p6UnN6IFuvibQruRvuuWz2V0EW7p+kqVCIel2Wx7qQteOviVXFb6Po
TOInfwpcAxM6oXW5DQWo2ovbq93fH1uUh4kP9LMYk3LixC4tUF9v3rJ6XZ1nhe4C
MyUbOGWVIDfkmB7YyqwzmJxrn+J0fBuFF0dx7qecwAJRjXmof24FTuGHYFdACn7D
jNqDw5UcDiNqUfnl7VKRlpiAdmFX+Kje1UfTo5mTZwAgxDKbP6jp17L16VmcC+M6
uvtelOGsk8klvWs6I/xRUVch2NNgucp1psjmwg3a0dGbxZ+sACDIcSJX2zgT9XKa
K/MYJwMTNvmN5lBQ/Qq96WZYZw3xd1Wg4ZOt9hCqKLmeoBjr71LzWXo7R6tvOrid
G5NDDUY5i5DzqQLF0KVTYczoQ+bUkOBTdC1wlFKODQt/sgBUIsEkz4m1Adp5oQjU
6Gl7D6uN8yvotw7QDC6cEY824qOoh3mfTEEszmf2lVlkMDg4Sqm9wjxk9mBVHlA1
ijmmjv+Grgr0F3vmynbDO3cRC9e1ElSKjdnWW9ik6ZTpk+cDOLQjWacFteGo6JYo
4mxyYgN7M2Cim60kl5Ools1TgK97EDmBq2mRiJkLAFE87VA5yoAzkiVo6jV9Jcoh
0k0GFamtr5lJTGPdYeYoncyTKHZi9PMez4ON/COatIDRy8q2BtRPcVfMMaYcwdIW
8Q13+IAeTr9G7BaTWL7/KinU4zku/4K5KZhgOVfLvl8Wn5X3r5wspy/mE0S8cENo
brzLDLCzwTsv4UbEacpC8aW2RzC75YMsOiVsZ6h+bdpEUkFiJE/uxWYX0/cI4AHF
uopTds4VlJ3kiRza8wE75uthx0Dy3D+a5q0yzMUm3O5jgKzQJ74LHzB4QKKxGC9L
fAWCkazuzK3eJ6wb4JUybIZvpKxJtfA/cE/W/bXigVex09God/mT6leAlBtCbmrz
xhHzu/sv4kkCS4qmrDzi0Zpsrd1mOuUvV40PJtwj00R1RJpfI2zt1Q42Ew7ahBVx
Hp2EbkK7okI5sW2GYOeXEnFntF8t9HM6RZGrRbigmzWsJfbSox9KfYM3Tu1vZGOd
RQRHADisSIgf2WKzYOJ9vbjrGMpyhr5mNUHUK2zCe1L7Io0lckiitpykgft3ZJ4O
tLJw6msg3fhyE3uPPGe3vZ+6YEThD1BDPQG18hgXNVpgmD6xabAil5PWPnUo3auL
UMjMwYwdntHS6JeSDVlwk++szNz2NU27U4An8E84MeLc38jD1zegVAx+6eEzDnk0
0DE7opl+1vBt9F+NQQucMiOjhs/e83UP1eN3HE+E8msb5T7QM/wTFA2GPyFdn2vV
1UspldR2ILp+GNiaKTFHgONZxpDuUN5FvDKuShhWKtps5aIKPVKQ12De5Dl40IrN
7I/6OMLZ3xpIueOf8YdmH+OLKaBHLPA8FWvUl1EjNGo0QZxslAORWEwftNfzt7GD
vNGEcPg4L6FNhMCfXRGuRVFS1YEVdb14kR98CZsBOaVs2qJDueDG958CmFqhdEnZ
0/YHhsvhJcpagEsMV1yYHZ+UqByGozFmoTlu7phILrtcy6/Veqq+yRb87fTsj6mS
yRIyiFW1dMgZadpWIixGg4rXly7VKFr7SFPxhkIFUPTTYPi6A9/64dOlHJsuBIbt
UwGK+180O3NLkjLpbzltP/uqlw6844vm+MZHlXyTs6DQ6pmcOP7HuFiIg0kLwhtV
S0ykKi92GT+SXsQBvL4vP0HbodbA0qAxJyIcTPxccoEktUuwNyUv59Z4p9fRNLB6
rSLMwmVhKltFpQNILiRBl2gqEc37gNfAtpeWh6GD+JvQuN9rxSoFWnNhsTwo7R7E
Tf7NvDJtU/EmeKI1TczdbAih6dZ7b5PBxDPRty8omgY4H0Y8nfbjFqNMhKoH0DKU
BQEI/hE7UFu/YuRfGHmqteUM2oJgGP7FH4izTXj/aQWMDNcOgse11u2v4xCqgpWb
PRAzWao/HSHjspcR4tGvk06gO8zeki9Hi8D9XEsvHqCXVM5m7jipgPyV9n8OlrXN
76wuan0LccsVQFPvopoNtLHzwGXGBPtwMtyQLdA5U606vYCZXqmM5O3HJvCg/Jb0
g4ipNuSniVRuaceE+muA2to/38pjRZSgPhOKIJTDDCn6QUkRKddT4l85PLYO32c7
Et+w+dCM2UoSt1HQKjJBvYQ7ozQ5qe8CvNPJeRwTtgc0736prfr6ipQiHAL1zeMi
smLxp/1TV1FY6TZVlEoL2EHvE69TMK15HyLAcCFoHaSsu5/cPhcD7jypvHXpI+RE
nFDb69CopSS5+noYVfAtV/UFvhCGAihFN+x8WSFH4YgfiraJj+Ik0T80D/cJ9RYJ
IDPJnTX+Oz/a0X16LppSbb2s9t+5gczO/4Q8fltcvy2+j4GeYA0CpSI6gey4LZxz
ejUf/XNU8GQaxduSqpsAyVHABCT1FzcsogZMb9QlDUAOwNLXxdkRKfrB5cXFj7AP
yNHQOBoFhsbLkaHggY0xUlS1dV2mX6Rz5ZZc1rpg0rr+pm5tLFnH4V/iGrCZ/p/k
Aj7rJlE0/IPpfhhsfgVm7muAaNBQ5qc+t7uD5sL/jzac1nYKxQ6qxFR6kQwt2KrU
ilXzmUmuI2fqoWi8SMlpOrZnkjVsRI8vRMzQXls3U5IWNcW9AizUyo0zRK4TZvtA
HU4ae+L+xdae/itfs3dd7f3AR0Qnd3cJz4Gq9UC9EeQLeV0WdIP2EsJa+YWzsXt9
ds/FgBz3vjYT90URSORG6NFagc3XOlLULEz45ZObaesDs+/hL5qDdwMBqzGzceio
SonAXT3DmleqFjlT59PPGgUgT9jJE/PDGmCOY1i6HvsUd69S8ojkTuaVPThjAK7h
gP3eSenbHoxlSxBMVaCCD5gL8xPfyRwiAqEoT7kcSpnvmtNHrEcRDJO/kMteXmpI
Iuwc6NJBfJvdFOuwqaTsNg5XoxNshFoXPmnhp8ed3C5Az8TyBXJioItDAxeC6rr0
cmqPcy8LWF2YgcNRf4f7yJpQrK0NP/Z8Goekp2y2rHs4AWXkwkvdBNfuZglc4Whl
qgu52JP+VgntXBjzlxC7HmiYhenarhBzKvghURNDBlbl0YME1Oitrl8PrTKkfP7k
GOSTbpnPO2yHW1t4MhqkhIJsbvEEyWABeJKHcxM8pXPbpnx618auFX8eUtbu5VFq
7vF4DFx3niGv966z5zJL77EVW7zdGxsNXiUSBfPWPFYIcXBTc4IAjS5Q8dA5puM4
J23eTLR7XDItoAGd+7jB8vEnpjEqhTIGyDY6LFGYV73DzLmsyixIXmH/6gR1PCpN
WG9qQqtX715sjw0Rk9AbGenk8ppv1W1U+CShkqcKriAbw9/amnmedBBpzleKitu7
kc+oqd9+g+3qkgE/CXosatFF197LC09epa4MBywhZD6piOaaDE6qriuhoZ82PCZk
B/kNFZiDYQ+EeQLqg9oNbDcgu1hy9k2xuu1tEFs80lr3bJ6MFNIdtC2OfaUiqHxb
CfNRDB6ijSCKdMj4miC/fbxCPnQFyOfad++kh31NDj7tLFxwsSJCm6uscN2PkuT1
+Vii+mBQI/msehFKn2Y1ufLW+wtkUI3WL7Ckfqvj7vXn7AOyiDV8Klbni1yoZUb4
PNx6IyUJ0yeWbtn8/n4SJZfqkp4jOfv88xTXEYHE1S6BvPPdV+T1uhQ/BD1njqMP
XE4wIPxbKXw9Uxmdoe0QsACWmSNAyv4KQX4OFc1ouJlnxqvihI1zReAg/kVbICrh
d81IY/3GasEIkvVqGTzX2AGiea6XECC10BcM6YgunT5Os5VnKZS66EUa/7Hld1Yg
pwIQbtD3DGFLNO1xBt6rUoalEKmghoU+9FtFDhzExC7R0kNj+rFVPLPNtpNMhax+
PbXTKn0kedqtMnpmJ15Uol6F/E9lY1reJJxbTXwEa+eRUOfzjJYD4a91T9jvNBWm
0XdGpbbfH86osMfJwLQRdti52rOjfz7DSEMBrwQwJT3AJkItSLpB8EV8o6Y2/tc3
FhBx5/eySHP1QzPCVHX6eN8N3VhhGPgGHXVSW2wzMftDCBGpMU3vOCNd3rhEIcgm
m4W1+Q8cDRyiwF2/leuGiU4zglXHhWFMk5swesx6VIUWDryqMErIF0W2HwZLI3BZ
q1TOX2jYhYZrTX6mapxh0zpiuK4gVJ/C75wRC+iGE4TcCoxexruy5s2pRvo0WnTe
a76bNHrAIVxkM1Vf4dAPvk0X82SQvfZrL71LXCK4HfwVsqH9z7kKA124Enb7ZPkr
9gLE2tXd0YmauYO/nD2KTWrYDZyeOPIHNu/TYko2Hz4IqmL7SXUJMlSeb4MK60S4
jgFl9YbHRk27AdP1gwjbeiG9UVZxcEI1Pc6BGAvezYuyYMgeI5oo0ZoyT05G4jgc
JAkGieSZJKZGHQjPGVQhSFwU3ampna7EFok5rIxG2iOd+Knt0EocLrfarxeo2uRn
Wift0zeU9ON+xTt8SNFW8i8cTdTu4zxxDcrZwqNznr63aSdZotuxjHrf0n/YLTKs
tt3dhG5P0m66N4KpupiFY/veoKK5PDc8KYoLy3sDP7x+42JbPN8nRQhl4tLnzUpk
YN3XZY+ydu+t/PU/e5LSiZ5qlPai+Ap0Nf6x3UHtQlG2sz1mr3Twr9kSnidHGFPb
mbtX81ZJr/SLjIGvx/o/RAJuPpUPoG5atd95bWK+Z1IfQ4NXIzlc/8iPkNtmA0dJ
3nMLFvc37G7N+IsmMHE/3OJTvlbwvzLJlW7Xtavt//+X3D4zH8y6vEHmEsKGH3Nr
w8F6MySVnhFshoq5KK5wqSRRgrt21Cc8BFICenfU0CcOilbJJ1RVy9wjhX/NM9w4
1LrvgT1biq4Z83vt32Y9TwmeHPX7DNhXNk4Pg1H0lLCrgENmTescbXU+ezvQX9YP
v2pP4JSladB9jmY6d4VnNMkOkbx3CISXL77+h43cRFGXEOiBbrTlNk8j8gK5JTcL
p5JLxw2Kl8aMe8ABFaMum5H99VW/VG+yj/7IvMWbdbWFTZbdHyzPB6tC5pKDOLpa
iEZpS0JinZ1EYleyyJzVodUxsEw8VYcC2NSa7OAhIuyvfNXDrMEIUZk9vBHIMfMV
ak4TX6xk8W66wC2buWBOR8BG8kNFTGDnuX36OHub8H0J8onddA3rP2B30eVlAWO2
M6yuphZ/li9KHIjyyiZkRor1pnadKtOQ2kqJpNz39ycnzSXxayLCh2P/NahCWzTI
M3tfaiN4GcKYEyzBLUUGug==
`pragma protect end_protected
