// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vit7rnw7gHdDTGmzimH5Ik4z5qvUTZ84pJw3MqJuuvAeqykPKxHi0V/+43x6oktl
dviiHanXWB7sslSPxiL01/gcBJ/jYXExfaU65A3AsZsP5sYzWuIIVe4W0QdGOPLd
s+W4rLDv3Nh1sDlnEfRBkupswwmbmlho8Rfcfo6iSd8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21680)
NIpwCZ5CxhXFR/JuJIckP6c21kBs2ns3A1TwMh7UUTV+wDdxujH8DuQqmmgRYDdi
CHNO+k6UNBNYcpoT4hQhc1UCcr/GUXL3Dlfplt623bRc4TN9uZwb6s+4tnYjG4NJ
XlV9tj0e1kjhhPBCQ7YIe8VIRKja+zcz442W+/rYGS9J3w5gAxytBB3FAlsOxljc
c0Vt+TOMTzco4PEwFMwDk6pR7Ol5qHtUziQmpK1zBbGs0VUZJVqqkVXpz2+kcf0h
4dQZi+F1luTL/HMD/K5TvB6ZQ8MSGbz+kyRaobCr89yuth2gl34c9fgTHu6fd2Jy
BnOQ2teez+GRh8IaPQoUHtO8N4614pVU9gdRpNWK+dvHcqDaajV7NjNqTsDISmIS
u+mGjLTChgYxiLCzbrxJC6X1Jdl22D8INTC/V1ruaTjUt6eGZzhICgUn/lE0p6hc
vQ0cSGTbjA46HHYQrIrzq/dnTrRzvvbsE4FL+PUS1YvdoQ9x4laWJmQfFkNdD84r
jUp/DTY3ttA726qyYoyukY03Jv895pKvkWQgKLkJiGx9hoYBk9E5mXbpYFXueqEh
/bj3ngnoZpcLyVy+xKfbFuwHEZZaYbKipXxzkj8gyQu+JZWA4nqKAl9PgGVi0n/A
t30nF95J6rvpiUGvpeMqx2utM0wYhxI7BvanYAeh56K4TSEM8KmhTrrJXYUKqBMy
ZOZWaSpeYcOaaD2jKFl4GPldptuzL2GU72dr8KWr4uOK8WlKrbWeUZAgmMMM5LX0
EmA/B6KcTJJhUtndUJMfouZqOIsR6Ian1NIOEhjWgWr0sxQpw9swwcp24po6m2NI
zACX6s/tIvPbHkCAQ/hHCuDDwyzDAyMrEtKb76rkAxzyMUQEYZMun1kHeot0TVjh
u0/NTqWGc6NR0dJbUiNRSVRt6iRX0ZfF2ZuFqtlh5amhWabXWJ5Wbe8eAFgnMb97
jAVAiGKCQVPLoJxpJOCE/bNF5JTKSRxoewSCYNnVBlWJru8TAqK7e5wiHJ10QgMS
09pyCKsk7QINUI7IQ1xzfN0Qss+R0B8KnUp9FE0Ss3ZQLD8y0TAWkIZa4Z5ybCGj
29KIucKsgjWbbVh8A6BhUPPmdsgGw5YswgZhfN84cfApSSYOrEsBcb724t90/zb7
LZr8eY/5JHf8dNiZHF9Tf+VTg3gb5TbEQCkJRg9+8rtzsBh/TEkgB8FDf1tHoYUP
endu5jUd85TGJhW6Rqv0dpbTTRLE+JWXzuU4C5vfTEwwZyyWf9tVnHw1ywa6Fo2q
bo22Q4gJgYzr6MnnbF1x0xBJ20T7sbajOQnUY+fh0fPYbHqXzj16oQ/oRrCk+OJs
qP/Mdvx9IuPdgI7rSNXf3eMCP8+4DEHcWpywidwrWNubslq7ivw+yikr5cDZiz1n
e/8xTQCC5ZRekGbLjOh446tJUqpu2/yGnBwv6h2hEfmvJWOuzh4AOmbcrPD7eioD
Njww2FSQOVP6978mqHvQiqMWYefemgPv1DSkf4zz0OT2/KZ0eWYFMB42J4rj2CiR
J/wb80HNf4JT7yVKdoAto6DM83/VoCwtfS1TGgnbYQXsWXTw2HrFSm7tvXtwm7ay
O2+UQA//dzfB2CkLyd6/SnQo9Qt2c/iKBQp0yDMTcWnH3Xt9ecLy3vsRgVuSU6px
X11eRrfrfz7oOQKNPSu+cBLpJ8CwoBTipayy9HThsQo0tksEx3RlCE7U4IcqLFEl
taSCkXdrco60VdhuQ2vZjWOK7E7PKf6ICJategG1oipKtETA/sDg09EqZYsOwrpn
1xVm14u72ZFSFo8fgQ3tVj2E0Yro2XX0HoeTvLdreLxOd4U58KAhq5u/Hi18S8qI
2zXcp5uFNJwjWjKFmgjlk1SJpvMGeeOzibM8vak/WgaPzt7OVDVMu4MbQQKto0XW
svVFU/GjQwbKZU++AVIbspcBf2Khi4pP5DWYp9zVqFU/psjAF2vtN7DCc6JhmIrg
URoLoEv1imUgdJTHIuI/0XaUysIz2gQwBQPkp6RKT/Tocz5zb9O6kq0LjgSpVjMA
7fKpnazBtoddT3eW+JXI6p8EKBygWPIdL7MBzHJ/TobPixsGU5BdCXHq/Gy6J9uJ
XGpET4UOBU5K6TvKnxKI4+6a+UfwIRz9QgslwcS28toPmnH9InB6TpSnjBcWfYhD
rw0kWCx5vVakekPwQxj1mcrqewSmh++oFdnc1c1CR7Ejpb4olLF6tyYQl66dL7Dj
98yE10509RzJD9C+WJGnhLZqIrfRDNzCSZJTNuGHLcQfRJqsxzDU2VuiYMF4RVBk
IlieGiGvLw4qH6hPa/jHuaUlbysgbGgUj7DGxlzlyWzFK46zveFumCdqmcv+ZYmO
GrVUNlKH3dPDgR76nU4m/44k9Ss/BP2666/cjomt6klHNve6zBYaRqnwhgX/1FKv
FwKOEdW7kxIgLnxmsnaFkjOwGcYw6/kEZDmSIMnDHwotgyV2LfUfxvUvenKdaZ10
+f4mkv8M21Zucv56HgQGsaPVS0u2UNfkIZgx8SNZILr64dpqp46Y2a2uoFT8scFY
Z8KHrHXmTItlKZcB7b+MXsqU3HovgH0VnKTRdAywfODUUmF5Gtk29wG+pZc5Muew
bnvsuB+PPSCOLW1oIe+Ocp2TN1I1+ZBMejEBqaxNEpDzo52oRyG0eYa/7Z9Dohhr
R/+UmCgr8GOw8z/Racz5s6lsLIytxVRrCVMn4e9B73ps8xX1/B/lGqQeTJe5Snxj
ZkmEHY849DHJi/96Skko4lAEke+xmycciEZTyW1CPHkRyiV1LdZarOGfOifEvYS2
C0fxqg6Jce797ERsVRkAIcz9mlTf+8wDIBSkSz1llxsk+FZSjCnINWykAhTa9Q0v
FAVHVfLBoCSjdZ67hlhtcnRqWbGWH09ijy2SS7rX1l/zzQ2N4mght1X8Pehz5/3A
0uYoSuOJJMZrCMxjZ4ywR/vQ2ZqFnBrzF5hndVJjhYRuX2de8m5PGvJJ2oBcsd3B
yk1Ejczsrckruy6OfWX8m0nH7P0srCooKxmdbxDUVlg/0DRWbpfGudHmPnvmSsmF
bZwFcqfn+0s77+EUFYLZuDti9sE1t9bw06PL2GA8UnGFPNhtDfuSLGeEf/pAuPXE
nliVez6kmwSbwrTXmAD8UTsSBRIX5rf+pFZB02OPrrA74/hNlJjZkUlcr1zpud2r
xk6u7RPDqNvIgAeIOkCW15LpWZLgzr2lPVEmAsxBuM1LZ0tERwkoQweUz/BnYNUl
tzwstjKIoGvucZk4G8ZXdV6DLQpihuTMrceN1aaJau+/OZ8S0JypcLgjN4qKgH05
5gxFzJqTd0dt1CemHzWZ6ymOQixF1XOJtDYxWaAwkVW1cgPKJ6vWhG4MPfE4Wr3K
zlOJqJRZxsJPlLk6LDXXDyvI4IgwkGxRozzv6b7XYQnPuLaalr1i9JBL6NkaovUP
TMHQixSn7tR/jqfU88lVswg+/0oLFY4TN6m63XoH8ZShOk+l4eO8XsUOqoT8HXv0
bJTE0I3Gvi10AFwC2308b1oXIWLyqhpzWgiLlVdA0bEi0jtAnMC+5PqnDIGTRJCx
QBECv3NZbQE/tkZ8EBvsmslOlkla1oNWw7w25/LXggtk59Cmu6KHP+aWZUP2ZRYC
pJOH76S7KAwBOfXG/5mCVc+GFqW3eYNEnXuykGTsLuNwk7/sKZ28Ft9Fi1m8Ci8R
NBd9n1Uq0XyDLzX+gs0fVlCZaVz59RnyDTJerBqGU8XBRjhSmwIWG5kD1722/dZA
SFRK94BBKfUBwrv0CKNk9C7tjwUw32Cl8E3JFkb98GyVExAR/CkpS2etcX2BHqA+
9FzZsBtYLWJbJ0PWvVbzROXpacsupqlWXcre9sc8QKTpH5/5pMGsHRY3GjtzR0Th
llpgrMaUKSQ1nlhP4jMx8J0kk+lt0q9PKACLk16uGauKylqiOSxFL2Az4olHMRU0
4GoXYUUkHV0pYd0V2VN2/K0J72NKgmW+0CtifCegnzz7+rOKBJwyzNJ6SCkuggGX
bL1xegDYxIz9c1oMLdl+Op0PPDdTtJQ5joCRzmvWjbR1HOIGM/CwJ7nT8NvMtYp7
7sZg5SzL8scPSBQRrM/qGmf5zxj6xv4t27+C4ld4hxGmwg4uMFHEmBPMAM3aZLz4
cX+KZgNaeE+KENmeww+Ni7ImUIcSLkm9P3jlawp4EE5bOZV6DRRd8Aktu8bHiTED
eSXomtRfefN1ClESpYJ3t7NAI/eNQshKIEZcfK/M2UCCpH4BKtGaH2hUlQ3GEn0c
LfGLkbRX8v4WwR43qn/vfvXhYjAJ7HMldKywHyUntItSWUIf2CD0LeEFw+kYAosg
MtA8BTZMkSAAFoRhkR45zbv5ylPh9WFoAIHBWon77/LqcxTSh4ckO8s3TqoW5d6G
AGlaujUbamzwnlvhC+TQCMjHENP+geqq5MpMShZ46EuRmSUWG4t2WsuTKjUemJoy
GOnJdsHC2klujO8kedOc4VtN/B8b9yffZp4cjdYUc7bRJII57vqEUtN3xaNNpedF
P2UvADed3eFUfWJPAMqPzZnbAP2pkfY3AghyxH1hmmV2YTKpk3YGeo0soEQsp/Tj
zh0JUIhoS9pNWujwsC9OeDRBhDoHnrRQ1JIuFzBfB5rmtgAD4t6RiCoMTihPYwv8
BuyUH+x9TTD1W8vUDH4yZuoUKa+JHX6efLYHOaWgDYdwrve4E0NRUjcnn+CX4U7c
d/djzS4UkOshEZpZR2OW2U/P88llkfCpPZl6nuezreB2XNADS3JOc7Z32cOn3WHJ
0674XDT42jxmhL43za6ibyXh7Z/gYGRZaS+iwYygWDORy32gxGp4CpvVDV/wey97
uWtyBnziY94nsoUKSLJlj/fjp2I99ZptIPiWI8JUAUbrCf3OnygMDkm1jDMndtX+
ifv4QFnfuHG4BzXuwFnGlGSo0gGNJR9E/laYAUbJXlWuaYDd8zP0qR1r0Xf5GFSL
TLidghcQhlXgcx4nfeQWAT6YJP4avmurOS19b3MMCanOzkP3a/CQO2J5Tm5XKjDY
QpxSW1KTWd6fuBLfaS3GIelyeF4pUMdJEofvhhHOLXnmXzRYeDYdQXV+KLzu57Xm
H5gK+sbzBDq/mNmddTXtKee6wuekN9BJzM4Ea+xEubwopUG+VnaJ9JU5d3PMMy+x
JY/pJ1iyAbFIh7z5zcrTsJL22iKHZWXZfZ4biaNcdQgqBAFNipYR82TiwUf9ytw+
z0w4eKYzmgzJojaMUn11A6ksF/UBwQ1qZ6/t/sqEqLH3maYzffhbIDPgMLOxYxGU
r3PJ7xUD/FlJWQoZiSmqZe5VVtFtnX9BRus/b4ueOYmkUbAGLccBA/TaW5/2VIlJ
654y5ruJZf+WoObpZ3vcaAqNzkXFLXlLasSbgVrU98bF/V4SJmSVYTg0CoZgjHUK
U7JYbS9ze/94ZJlFGWQdqzDrywqdHeq2g0GjATFe5r1Kurg+E0kZ8mQvsRGKGvAy
Eoxrx86ppfajIIDyjJZPm8IVq2HgFwlKT1AWSd5BlCxDFdBqhB4p6C591+MWXs/7
EJCUtqeg5AH4a5I6NMgzV5R3mS0kXwVlbDN5K9HTDaWOVufCB7tAHJsWWPqIiPPl
+bynhwcSjVCxZTdagkdaxxScvNW4Bei4lMwTlhohCfi90HSc/E1aRCGkOdP9L2gO
Aux9gLXTQ4OV/ofLQJdvXOnpm5csiC/EQml4D0xfGG+SFBIoz36jX+UsW2p4J38V
MpQvwvXRT8DD8hoPpo6Zyby4iu+Fot3oCwUQNsS9UQtLCIVSxjOwwZraW/w8gDV1
ERJG/q9afCUaDdAA8yUi39uvx4xFDvvNmqOZ2g/3EccCPXnD7FX2srLTL0kPf8yV
6cgmWpebx5hlEMLrumTu2SkNtnXSbO1ScZLtYR5GC3FzJmGWkaRRkGrVcjiRJh5n
KRfpR8tD+hFYzMNAD/LFtLoBIBJAV3Qr5/1z70Dk52sUTowQ7cZ1haDq2jaBMGRZ
/ARFKJP+W/GWcYRpBbCLWnYRs+8uS7MEtllQBaxUvi/O2V5yEockKcSOgAquxLdb
7NQqqzpmGxMk3u1yAF5PG+1Pqw2vbpmexZct3BCV2PaJRVo/8iELRNB6zB4zbq7J
RgATZKecGE5oRhaWzQ9C/O0rbawl0Z1NByVOSkGe/8LpUF5worqnGI9+MQXwKyXr
6E0JjlsnOPRkNp/wgRkqk2ePHvVSuc81hPGHOZoqgx1hoN2FNi4ZCC8k4gC99PdD
YFhi7zoF4LILiAdr+kcM+XXD/KQiQ75pFxETxmqGug/4kF3OcPPA1aQqWTahTnCJ
snPMj+zCrp2civgLL0VvOPRgz2v53syKRSlupxVjqcr7M2EMavGqYC2jlR8sjjrN
Hay6SUpn4TVBbe0Cy7rIefIXTpAAPmkuBdlbTBGc1S4tJ5mm0+/s6ajclDCvY3Uk
eReFDJc2plRemBnS0yA5KfUiQWPxpq/mTvUDeEwW4hc6lrO1WfhtKZyvn/q58gSw
Cd+6TR36pD0Q+QMD7PE9aVeGIuhexTDUNSSUVNmzbKMywdsPfi7TkeReNZ39kRLJ
NYMZe1Vzl+0GA6gF/zvppIRj9qBSEopQYilt6mThBhYQc1P5NdLpIuwEG5bFMZZj
3QCgcgqY88a6Ns18dTi7lG6v4UmJZh6gwFFe+e2hHSW7tZlfDsiFzPrfe7v1Y0GP
qReeLw1OOJ9rPmNOiP0OOYx38xyZY0btsFOYrmjcaHeFqi+exKxbuyDhA/qwme81
Rvxuz1hrZh/PWJqOVUFAyqsItRMnmUkfvMJmoC7l9v+P0rRUYE8vLjDogOn0DNxD
T3amu+ScVggF5kfpIYueRM8Az3/Hw4x5OURY5aa4+Mwp13iC3zcIc1HQS883uqDh
xBiSiqTpHbOIPOH9D/tqq5c5qrEGJPG/Ye6ExUPzU5J987KklMs6eN+cesXJqyRs
tWuNKd7+zEgtUw4RyKaNbqOr4Knuy802N+LXvBWvWLTey2p9GwVMPZeVhMIjhpj9
BGkk9gOulP94jAwuBYsdnCeo5JvAaw+4kny+Jte/g6M7+zQnDZ6McYBao3Ubic/+
jfGEwlkzkowe4Ftx8p0XUSG3LCSvQnp42qSl2Uj7khmavbDF+0R7Bn0zJobDQutt
p0MBxgmB05/fzige5E88ve2E4hy4f/dnTA+zaIUkUuE6DI6dr/MKYTsxx9xgIotc
Z8g5LuN4ASFH4exSOxUqbl5/74AaPjBHL7v52tfapdFz4DyFMyM+tWaCoRqRPgn2
UaESQNTLDWtNX6gyCBbdJq3RDooeSt9yjCJYygobTNzvCc4sMlX20BcUsHpB46Zu
eGtxIdXX+AmluN5G3yFHYvE5Ncvd81UyUOT8E/kVOqJL8/yzb88ccMz9Eak2WWeq
1K94vhyOjTABRxOnAulcHUBNznCg3NYCce1KdZxveCmmvFD/UlQvKUR6XuYMoM+G
wfw1QZcnz4VabjbuNJ1T6FXxH/wA+T9WVn70lItDsSSN4Miyr3VbFQx1Gp2KVhf0
Ahcg3xcgCbwnzI1e7bbnBKuPX2lFyu1go1QdI0cRB9Hk0t3gCQCDc5Cn2R/s9Rhi
yArqwM1o5+YuFZp59pBUnjG7JYxxWOhzyEwHmf0PcLOlpZ9zU6TCo/s0YVaalLQZ
WIpJGyq9UUU2JbrWQ/ZNt1/EDPAHcZIhvwy7zZm+nm/mcQX1GbMhEnisY7IAqpkT
QPcYSO/NAnlEHehxjmY7VPXNWkRNcb+Hrqg/zpQXvavtCZ+sZTvSvRaSf8gsxbxM
Nmkvqf0Ywgs2QdlQfx1XIJD40YaswR69bVT24tKt3tygQcIUl3dxmhMT22qm4bpX
Hqt5E/RzvzKh4OI/WL7MQ4cStKo2LSw8MYy8QvO/wHEI5THF9Tcovyqa/3MCkeF6
t/BVNMgj44ompsRupASFuytJoBYvoMxyCPTV3Q6YWhsAREkeI2tyPs/q/hmSALQE
3mbXc9EsLL88eYKdQQkCyGdQ52B+Thw6rWhF0A1xghE3KbFETTNNzd6CnKu3QUrv
GMtSyHBfAds2UeytN1QEfQ7S1xF8MieRzMI5W7euT1DHHDJH0bicC1hX2HBVmvN3
JLXYmTU6QTQt6o9QD9PlAgHovIC9ytHAvCIhlY9X5MMcVhHyxgVOmadpZPNkmUWX
q5KUX+VCiBNjn+vWxRh7yFvSf6eQq2nSIbs9xdsXu9KM55jZPcK3arngBapNGgTa
DHuxZg27/vmpQkPlf3d52LNnNSbg/vNdFXBULGZIeT8Xl55twpApAGD52VffZx6J
gUGfKLgfFalMANLVCHVr48O/tfGT24bioxQBl+YGIVpuJNhMTxJLTrbjqu9kznBO
P8B/usXU3o465uJ5+tcnK4cphLQhOJmtTwt7dNxTO10Ly4j4/cuksxJ9e8UulOqk
2y8UHWmwmcta4WIs6GR0i9Wxd1cwXn5aioF9iUQcuOOhn2vIlvg+BCNu4fLed2N2
hV0eeAdLYvKz6KJC9Lweb6HpWpaWfd2AHyw/g1rLwsl7SBQzHaT5opOWlCnZ4+LO
Jr1n5rBdpMVzile0t5QSzryfV+Ci1DcDPdyJxH+XqhTMYzbeuO6WJHfBikx9n5ke
l6MoQbxFGCafnhadfmNn4WoeDD9jubNx3e4C/NFAzh6QBCnbP/rBPdEZP3jYBXR6
CBwrJnhV9EGr0sD5zE2nD2KD49W457+LShUIbizryXfik4Fslr8ALWWmKj1TctI2
KlJYREuAbGEGAP4I98vJxFx79dj9H1hHMYW8tmfMqQHb/a+OJzgvJmjUGXkV7wS0
wDzlk/j5ehMyI5G8KAl690Wibzojwg4jdGczsj7veZEhGZSed0q12JgJrvOGDiRA
eCf0Ppsl2dQjHk2MtjF1OkIyBuQ4RnkftAdgmr6iPHF25UacH2RhX0It70aBGkWN
i2l4IudZM216TQU9St6kmsAlJlk+EQD8PIjJNVEVhXTFZYTQxm9UlaZpNQBpBYtp
8n1gIMjyYBm5Wru1410bcv+1+8auL6D7ZHHdNiflFmgOB2IFxeRfmfsJeydxt2Yd
eEQV4JmqyUlx6iC9ssDo1LEukjtYXjqoYxuzt2RcOjbUsxMnGrUAjJ5vKndMWtrA
dhbLh2ZtDDd17oU/TywT8ynFpuzyERHqivDMsTLSsKiMOqy4yS+53HSPLYu8VgPJ
8KFVlgIF+ryZVwBhIdgjTlAEE3dQas9tU+/5K/Tt+sNpw7O5vF67YyE7+y1Gk/ZN
+ZwiwHshpMlVMSu3MXlGDyTNVipkvGCPg8LVs917BGWZNmr7/8d3e31C3ffbu09H
0jMwlOw1Yz0idk8M4b2KKQdv1qvHY76wYPXFGmw9fMgmL8FA1Zq5r5FuObohGsE+
w3q9Y5axwWfl7dlXxCHLG/9lgo0LoE0JmDOGlvj6Jjx5hJSFCpznd6RFYPyx7IGp
bt88iG2JnJfmriPAFNwMrHj6J6TQ3DRdYmxa9qqS2YnCf6PBcjrjafKJHR/q6G3a
Ta/pb8Cx54XmYvCteve8afMcP94403u0yg1VfFym9KL5c8K2/4Xn0xrTuKxLfC5M
eFH0Gbp/Ge8BayVpxNH8MTAOt10vdqWuFS1EnCAHocisCeDBZcT8xYQZb2ygqdcD
XFUYPzxKN15oiwjsobRR9SwFPHy8LUWC+QrwReZyNuDSzJLpKf7T8IlcLr4nciAp
2F7HdpMs6eETzY1wYye10POu6VpLh2aflLosYDvc1rTK05Vcos+PQKkIUVxlh0wZ
ssKCKCyvJWtG/oyziu8y1g6nWULK6FtQJ4Xhm97+QQKAq8Zd+BSA5Q0U+i6sgvQE
vzSVdCBTw/BZ8pycNjAmA4fLRkHWjR55hd53BtwIyviiQxcAI1Rl+SKpo1HCK1gn
olZ5X8J8HKSZwrwcfng8a+qRQfDotO5+n6kPWfHK7d0uk/HEJpyl/G5q/icBWRbY
CCONfQ2jJGaJsF8ZG3/IBTNKGEIM78EdTwFTszu/1igS1bCWg4kWaFNVuhXLigAw
zuFzctCOVk0nu8/nV/2gt4ztHUl0+nvFGYPoCoZDcedq26UlwddB0vTNyh4iXCgU
dxqig2QWH8fPDb3UC5HBjj4jFBkThpzVkQpAdr7t9BAircJFnc63rH67IohfezuS
nf0jQTtpJy0twBfTmg9XS7lPYgSrnejSzywI7C1Bcmu+ROUOJ3vUc/GHmM+ERknt
qBUWdnUih2Zpz0aw6OELddlTaSRfz0/VOjGvFs+yOv38Jhh7D4bjsSK6giLhXM6p
KCFOayWh7DZ4WJfngS7HU+kCF4C2+TF0Ok7I1ZBCWckcpd90T/I0K4EM1RdBIatO
CNORdj63dBQ0uFkC0NMJotSUSFprHY4lRimZA/EubGlhgv/NVpB4es7xDwashmQf
KM8rBs9TFR2qyYQLNPlCOtwBgNzMK49NqH5MrYk/ckCpdLc8mbJtmMg5u4ONVFj7
um5U9vudBfhym8pyNqtqYOirRmgMKYZi/c7sbF3tdvtMmxVMXEIln4oDHsEo60hU
rXVqQa1dVATK2Z5dKHTFFAb4IzLQuXZ52Ql9JqLqoX6EcdDSAeCymEPlQ8Wfupj9
c/rkJXn2ZJZI4Pld88RL0j2Thra1hBzCqewV/vfL6q/zRa/5gXiyQBC7Jj7b7ipO
wWJ9kxGL6tyH9egRe/miQiaIczLoce/9k6jsHCaguz9BkMp/cc5wtCU449ioIUv4
3OdQ9xSz2aDuFgI+dNf2GIW1J6tMi/3tnXx8X5YtFobatXPU0Y56o9bn8vFan1yC
s1OsUMUBM2YseukT1qXXj7ETLRV009r+8lebOa3LzV0gMZ2o+om5GTKqNMDjjh53
ykgWU4ppaAlQIpeYHWMpCezPYvHX3WwSHMe8AyMj9nZ71uaU/Hyj1g8aMF86esKO
Z0v3Qpvse/0DvYz+NdWJEEbjaVVFJQiIW5Ho0XnkagB7eLyV0Bcemsu872k1WWQs
DGq+x/E9V9nUGogHwFQj5O9nNYt/Fw7zGxV9D8/LCITkBUdZMmtlWfJ+jfwDF9Qy
wpb3Fj8siIQgu7bLJPoJyPtCwJjGuGAHGkWgvBRgjES1X/hu43IXkkWDkd7VK3eM
ZwknmZoqoH9BEvXjrOKHeJ66VLdaQR+ofPy2Nz4WT5H0r1H7FhHiFxpL5eHG/iwi
a74VfqOk4s8r4MbHhz7m/Y8ZdHzZftIolelqVtP6NQhStQkkLwptRl4jdc0IKsIQ
+V8oodXlyrLY/wuKdoa3Rj23kv9Gg8U52JOKXW0mv5uw3/ELQ0u6JqhAW/4HIPBd
MYzwtFR6FlKOZQfa0UQcIoZHH4yEKDJ1sc9dXQTfZvz4J+B3ZgP0OUaAL4utmAzC
ozQCvfLNTMSsj4LMoiziVJFZOiJTBkIVnNxCooAuJY+wxW1XTxnrX5GNppqyvxRa
u5Uu/MLIQii1BldiEKeQV0QbGTAJGel76BWU6BgCeGL6jI80P04ag3QXMQ2fovGc
F4WwfMsjg8pmLfwc862a79CWBA4pgvMftbzrQp7kGWA1Nw3LS7UKnEXrEXEveSan
d/5dhXpZ4Elb/eSXaobZyuUcAkbZL2pQdPQdJlf/ZTZBYBIMUsvygsDjqdNtxl2n
piKc/+VjzD0wNLEtmRdi7ocp1KUsX3EAkFA7Mnbf5vMiWbDkr2dWriSv0s+xp51l
ob15EnLFXPa2J9qUeluSfRPfy9M+4lukdtDnRPjpbrfgeL7AIDiTk93qtrotW9RW
mHKXdaAE8eI6n/ZXubqcCmvO9WpYJ1wxpaoZpnZOxlcl22qPLUFJEtvxxvwfKqmb
CGpSDF7GSjRkU4JbLxx3Sb7LWVUz9RT8kEduGzBWZz8gKHyHtAT9w29QsIboZbIk
tpSfIZHH/L/KXvK6Gwxc3qv+Yej/95E7kXgfeKFmIO8VCx/NNCSL1RxFlzlhYEKe
MetpvheMV0gnseIaIA+ZAxMkJYzqB2/PQpJKr6ZA8npWTh2203JksmDTX9wnkADP
Z0WcN9MmTLhgdwa5nlGcTyO1YSMEJZgtH65Mc429ARotVIEmhK2T0NVFGk6t8mxk
+qulJCMqBydgWm0zRwtP1CC9zzaPHqW0DA4zfPpqOi+WxWvmkNL4L+RVI3j5q0cB
J1gWmBBebsJRdsHxJo2GkMwGs2SYAo3GuUbG+SuuAnnJNoDBwcS/P53cL2Wn5kxD
iQlveIONsxWnxArN6Uh9BPuiOwcCw5rT9J+DV600LCYNxHLXK9Gs3AgerMb4DxZZ
+mnVS/kkYe/MO81+hE8nXf/gfdbAxJ0NUcOmd3ukGJ8FkIwn7Wj+z9j9hjrsn6zI
aIVe9bUB/1MRQUobCYF1fcp5l+6U9QdZsB/0cXIAKZi5RzmdUOT/oO24/q7v2UZj
jZWjFAct8qmq7HcQpRZMN+aMIPvxjI3mda4vja/Eljs2J5xyTuz5bmIoJ787u4UV
gtTr3d27YdDS+BqQVBZx9Uzv33nURK3CWorErUGFRoooljRha7x5MFraa6bENibL
7B3gJu/oCY/BGUa1j58Nl+ohX7ZffmJKCf3eyWkAKvsSA8Gd5lLmd/o9rDVNP6jf
DvEl6uiGmLHXz4F6eBspUdW6+Tjo7+G55BbyBhVecf8DXSxm9KKzUmiTbQViS48N
RJtL1e38UHY92RGJruFRwMKafozRJflzVJZOWEcyEcjJuf2DKWOtTE5z+mrbTmxi
vovQnZ1ncO0VFaSyENiHKV7GptCvhsok2P0DI0ECQ9mvmuoX1jWWwtKEv1dGSIL4
8cmrIVkmS7it1ulLJvejX4wqUSuah9hvRgKhoPQbPxRs6foMP2nWGK0JRTGnqRIR
m4MviEIHXfQw1SWRkodJtgWMXtfYooEA1w4ZHxolH7o7StWRfovQerWaEch/Y2iV
IUgc/am9UCujYUVwvk12/UZS5OGca/wvp8zQ7aKAy8EoaIDG9H/+8gSFT3tGKqF/
GtGsbokWRAzThab/4eBFFr3sox4a2w7+FInCJTro4FIdXQxcj2XqlTX3RxaAPaG6
palWkH5bSRxAOmzQkoPy+4yhWWmaczyt5m+n2LxVcrjxB71vogpTDIkJuEWPjc0W
H2RULH1qNLK/N8h2I/GygwLdSuq+ecfyap093SFAC0a/gPYB/P7vWiMQIDR46RXH
dmKCxQUFO6gMo4F9j666dgo9OszUvKij1iGtcx9Rz4AhqsqH9yK11pPl7T6nHXES
3PayA4YaL6eWFqxzpmVWe+fyk9nbY0ek+gnaE2bYRJTpDnSNbPtOLT85AhxnDO1G
/AVCpJlVKcawPtyXM7OEJYmijtbkkizAvNJkvaP4ZMJD22n8/WvD0f3U/GBSEUq8
RYe49grkcZGYNqg0HFPSZFMdl7bWz5xzwXsbBW1eZDfjeIH3eBEWWVIaaW0DCZjx
7aBlf5U8wkgsn0DYuLQHcTjx34QBhmjTTSonFIR/TbWXeOEh4vWMppB1YvrqTMc/
N1AKg8/IXPEqB9Q8wCJ8PK0UbTHuQLHPO+JFe5j6F5kzyJyIscXuQRvpovbMVOz3
MVXBlve1076arwF2AqP911dsuIpRok3CVPpZzsyHkgMjf0g8ZpcOQJvU6uslHTGZ
obobKtGvPgznIY+E3T6hWbY1/xKI8RfLGCpJ4yRnlMqkOQOw5ZEWYFofH2Qnn9+z
nE3KoITbLhmoKIWAVkkVW/bxmF2mwoBbL2EvhCe1EOJe7y4pexueXM/Ehqa4C0zx
984NLDPQMdzK73i7inQIE9sjn4XvksE21WQCtZDUb5RhXBoKIug5u3xyY0Q7YHRu
7wT0h2PiMdGRPowt0G0N/j97bLd6rEXyIiyjMLuJd6bC/inLa13OvpgXU3OnWHQP
fsmddkOM1tisuRIsLccg+7sBLRoGRu1J+ttXu/lWU1p5DoZeUvNXvA1Ve8+yKCkS
5wApVxzgVhUDGyu3R0ruTiQEeZ6jcN1PF2wntG+ZhWuXehozOOtqL+HkK7PeaoGZ
W5ftldDHF0PfUXmhidRdxcClzQIL7hIBWFqNhg8rbO4MosQzHVEKAjaDd+/DfePo
um8uB7+tCvY+7zJlTaMQFwvtWxW5/gRh4mwUlBMbRoIdMTMjHlO2zFjHRCshA9uu
SNf1GN11ecwELhk3S3vPMj3rijjLiRzUoOMbmj9RfW8t6dtvQl4nzn0t0HLd8oBJ
VBlpXIZNSGhjy/UueVWr0zrs87xC8NdC0JSkGLvUVua91EUTSCBYBbwXpu6pviv5
JVgkhsx4WlUyuqLQRT3an9MA6yOF1wDwgnRCQj2hG8xi0rzyjHAZBK52zwK3xIqi
zKxgWbdwYVWX6L7vEg0Os8HZP5I4sNmwAkOZD7lwhGg/CpXBcoTbxqV6pM9RACbh
QwI5Mpn82g0up1BqCRQWESWsGa3jWjO2apSVC7MJvoOyNMKn9MIeQx/qNpUc5+TB
PAK0je+A4XCoPVXmhkIA39E5T8PSGEyrZ1ZpePMOXSaVD+bB9MbJ7RdBknKQeHq7
Jd44HdtMBHO78Regb29lRryM0OjSyXMgh8C9qflj6Su5stywDW/3b83SLlJ3dB0T
P4c1JAonMN86tqtsAQcjjLG7FkinBnubwRBGEAU7iASOjo4f0XojOK9NJ856BfLi
TF4TsiShkEeSVHalahAyvUlkGL9TEjtStAax1E1fITJy3ExyHS739zazt1HMmhlR
DOzZt8hlVEpHbcsLwta+w3UDdSUGMfNV595mVLNCcdT+LsaOzapbAHVbI7dD/V8G
8B48llSZsjIMQVsIuc8S1mUukDtRol+CGTk4CfhZO+2ONJydKq51lGwZ9lBk1s8s
Ctp/y7dchLfO/QTLxYfwzILLNbiFC5vRQ0tNUHp+aQoF8W/gCKx5Ko/0Xf5PxF+X
d7V726eB9JjgROYfTxihgcuD72O1xn0C6HCIPiR/Zphl4i5WyotCU3MQOjCJav18
SihDxdr3MJ26efN78i31NADtkim53fQir10gi7DQQDIWDE4NwZ5q3mHjjZpUpvUL
zsse+3N7MmEKcgqz7zhGoxzoClHn+CIbNSDqOd1IDoZY0OGxgqnGju5ZCHqpNDkn
c2H+/OOJOXrjWW539LJ3mr45ABWKXjozIu5C3RPmOP2myy6smRlcCW+61BqMCSAQ
w20qXTk0EGAAHpuVGvQhblxJUw13c9H7iaGoVcEiIo0y4eyiQcEcA73/L4TxUGtk
5XIU6x6dpthMNTKuXsFrT2rBdTEzg9NPAOjJm0imqb3xipW67VS1VJZbxsk8+SKN
PqxL2vBS7hGYWVgr9uvZx+ZR6IfWUGOnpkSqo+HsUQXE7tMmCNoWUQHA8GQmsfqH
3hxCBuWCFY3I8acN4DJ5Jak9yAP+dmOMoI352p3VWWIFXfP6GuO635aW0nIZgCR/
uIr5Zk3voBJ1LLqJ3MD/ZWqiWY1Ssm+xX7prrWBgEkIlr/wN4nb1sg5O3Zxt2oZf
4aEvrNocRtliLCPVSICUVse1ofsSQtqLZtTdnsJPaIWWIOr5pG1MVx/cYg7cEoQ8
y/jKbvP/IjPiNeBPX+ZW1Qy6n09yPQPfNbw03mSS+dKtLJliQgBtu4kwcCHUGwXv
KIo4jgEBQ1Zof+94eyHHRsb4e6lAagS5S1RymNo+FxiJOU2rDSy3PkptbKus4KiT
dZi78dPGVuF16fNIBcJwz6IU8Ddu77VJS5GAV0TLNYV6iTokpZ/W8F1nFJu5yGMg
15d2rnaJcjWoKyccdtO402U5zOfPenFvOv7Yjbc+khmsaOPWA6a36Vi0NK6PzveO
dysQ1acc1C6x50Rb8GzDogtfkcnMiWg1kAAZG4H5MkxDuND1wsk8V7H+rCeUcIds
FlkLqRtQlMr9YN/JUnlL6xvjmBierKKrNv/RliWHO584buu6jLmkzb64Aq7iqKMd
hJ5/jVD2lPMlnkaIEmv0lT9QnHDlrZU62nWFadX9hPIT/IOOGfdyqcUBp8I3ZtRY
Eajqm42IBPBhFNdAyXi5gmUDFhii+IpOSEy8S2nRHjPAeq7u6ZcjpDoOuKpCRFqX
dSTBxkf8N7HpfQ7K0LH9piloidcnQzng9ERKOElbLAJtJOhgQ2j32SfeH+UjmAti
Zcrwq5HOf4pncKZRrIeBP/WU0OSSNYv8l21+E2JLbdy2SJZCHYU9qf8NK4HWYTfe
x5K0aFHBOeR3koHAK7UNfNxM6prpC3xYSc/c/OEH0L+FkmLluDv3s5zTYUeQy3rC
GxfSefacR5aEzupPfmWAnBlSJLcuQMPdOBtD/9vBk+ccat6eMA7IloiuvVh4CUt+
BxN/JUhfn17HVi6vJCKC41jPWWqc6FlSckbvAKdIEBs8IgvotZiaCQHdD7PNRjSE
NZCzyBL7UyIbbae/wubzU7G++9dGIQiJJv/E/0SqgcDFQMKKjoUfOeYnyTbCBoof
RZdIygJSUZykZJ7EChvbZAfwrR2rY0QJTmfqwhq4kzReSpyq+G8/wYgLDcu7FCBQ
qHLA4Dwufs8uTsKrkEC5zAuY5r6ua+OdA1UO5l8pppSmTiQ04div9b5aRn1ehILV
H923atuCdtygIfh5Y3Q9CGDKk3M6ddPYIeDCGzpzLATYFB2uf2rVpcvccjARhn8b
NGQ8dWOJSmVAfjKNe6dkxQ4qmEJyYdjGv/XZ9K2mWKNguFv1PHsHqEIY13CrPmbP
xjgoAubpSrpnK2Sax94ce2Syreeo/tQAsOq60f1f1Rog4jtw2xvQHH/iaKbu/ycq
eEU+PfT5B4v0kN7hd9esESKpCHphAqS9NAC0aTBDye9bpY16QQnAgCEB97jZCDw6
jtHUy+L1wEBw/+xBTA2+E9aH/DCSQK+G+zcKMfcW0nPar6ATa2yDL80QhdnNunoB
L9iX0Fmgt2vOl4XHlNEfIXIh4Kgl82WsXuScMcPVi5qkwwHgzSx1lkTKmTLLsH/L
SIlYWgn77CxZGghI8Tj8XkRbYiWbyAxsXJO88vUu0X0CgR5tHV8xKJMzTkDDfgjP
W4SZdiEI4VtBdJO33SiZLz3vTkTevhb1U00o0TtmXupAt7AOHcivc5BQMBRWTPNX
t/XIrLa8f5TtXtEBqi7BL6qDdSKSzaC+8dIsumV/Luscd0N3hgh5bPUdD3ytdwaO
WRAcXGof+Crw/hunGvW/oB+Zs9UzFlRLCwJAzgdoPPZFveFLFhB3GHk7Vr2lSxjf
373n+yrRpYAnTUlDmYga9+EcdJb2fBcqdxbeG/mxqPLAyxFYRoMmlGVQSuACpB7l
+gOvAlfDadDZV5qUXHCcd45y/rr73WgdltEj+0yvK45ttFvSvINhObeMvXil+cVl
eJpRyppoEwXuVYvZdrDRW7NLXwjcDFrlUhiIrBTYy6SJ998rY0yswmSy8PeADb3w
WbHYrUyQB04oRzIEZhSKGyMrgst35POCGTyWtGtQR4Hxmag/x7LxyZqUf5nfSnyK
i3Z2e09D5JqzIfA/dm55jgmlhs2iRCOIHdiN4eE93rTnX0/ES5wjAc/zzFRluRfN
v+MURK4qdyE0CE2s+PtJE/DBx4prFgrr+RSBgt69c369qFb7T6VcXdCqZEPXgxKk
Nm6ocuPuHKgIBqdbEfbkwN0I5Y9KgfN0FsOAm7LkekonQfb6v7br68hUsDTarJfM
h0yHbbRS0upC6CdUCviI5GlcKEOgoTyEm5W+YdJqt/m4uScfMprIG8IjtsysyZOL
RvgLhQBpPGS0OThw7k0Q0v7OHaKUB7NRU3xMhNFYoOrAreKILL9Y8yVH35gDHUP6
nm5a+35q3OTP8bylvoQqxif8tfEpPoBHK38fprvu29vaxAR2Yt1eCdrCg1JGmI/Y
rDFqs4SwDZfnXPOhfFrcUVoGtLhYNK6pfJqxgcXITMGgeKX39zSbOXyFh2a2Y1EK
qI43YKV1vj5wDAzON7tf22L5QEAP9u7Km9SPZJk7bY2uZIQRgnhOiBLJ9Zvafzfh
aPnWxD/sUkM1OU0h+OxMnYt7JFB41CiMPCL2JJ9VudyUWkysW+iYgdVwkNz0FIpI
79DPmiL3KNU6IWwKQtFCuBuFI+RVGKBWrCxevjjvshfQ+3ikMf940qr1ZRpRk+eN
JeSUbGW8/jt+pAuxF9/z+sYvy8L2A+05Qcg9Uw1e4M9UH9C5o8Lr27nX7UBJFIWp
c75h7hOYbK7pXfTVlfJ2/gkfHe/ydR6O+33TZY4cddMYgpVxWnt1t2LdB6qV1BEI
iqb1G9dmMfKSzMueT/Chr0HQpa7+HffjoUFU3PwuemSvhYl+vvbjAPIKhcIsob4r
vwaBRFHZK0tz1uVLRQTWujyHVOOrYw0WXkHzGC2R4ctSC43744bV5TwbB/VDnEd2
EQPakJjui2oybJEDuW997vWiJLtjjQCGRIaAYvnULx6+qNCbvImyhDo6vqybJc+M
3MLiAQmIpBtwkzI37G0SoFfWJ2q6qF3ZNz+SSXQ0PLvWW8Qq3TdeBKnbgftRqOcz
XaDJyN5gr146bBK1yCDXH9xspWNMXiLzhyigVOwXrFyVR2sv/Nw4LT+qt4xSPzna
7b0tfHoOs6hN8yRBxUie6gJvL44cp3zhtBtFKCnhNsVeqW+sfeBQ/b2FNGxBPoTg
6G4E8dbjkqtDNfvbNpwRLQMYbrmDnCHWuKErFcE3GZDrWjsNqnX2hAB/Y1OoH+Q7
912B9lvClnVnnBChtldXEZn04fIujA2AUad5gBMVTOcIDCKhtro/x1jwWxqS+rAZ
RuFFLZVVVjyNcFG+ui0b9JkzTu4oSmtvxtFYV95nT0nidQnKNA4wDYKT5IKo6uqf
t2oQz37zNFR2LzX+TQ6cmwigSEOXOEZcaNfeNLM/sNdIKrOhhZk7KElzzp2PT+yw
MDejgTKKc9QapSPYSLIIfJ/A/rc25Ouubg3yNN2HhnfRvjhEiReIdJNurA5LEDJY
sPFWJnPjf9qfITJzCDQer7bBgo4Zd3K6YexhsHa0SFx2aQCKN1f1TWnx5ylKtyEu
ZP47mc6z6s/qD9zI1qX3N215O9rXm9N5DasKDNHgP04+wwoETz0i98lP4oz5inN/
zcWJ2OSWxWXIWnGafliSkCubQy+wyKOG8reZgSfaHXEq5/WD+yiXsm3PIZs13tPz
1veo/NxatgyEkvfHeuR8PHtgaT7A3KIDAYYR/A/gx+VjBjlrp8O0BD1rk7tJnuBM
0ehnCXHS+9jK4A4hrCYnU1oP1F/eoAMyn3q86X7nTQcsjktKOxrXQsJkM/IU3vf9
j8BNt+x27ungz87l0G4ilyCg+gOpVkdgtgBgd0sj4mYZ7WLIVZErWBegEgG+NUIm
bB/Ln8mCFxr9OZO31WQxzedsRureNUtKlhITjlNu43HwAz1dAJvydVshgRLN11Fj
3EvmpuH+E9R6vknSQFZPzT9KCwQun4CwnKCXYlhN3N/mJj43ntcBsq2te5j2qv2b
pnmT2mbu/2YOftTAvLV9HWn3pkswOiuguAFZE+w73e/d0KsMv/cge4XuPhpfzo3v
exj09jd5pNSOeGDUTNNUHBR67lFs4VV8eo0GIL07x8KjGfxLvUtp73UFBTSmGqwt
dETFlBagZNZ4j7ruaCbuoCOZu7SVXhvIUPOG/0ictAIQvhqEij8O/iN3IovHhrRu
2KLo8zyw1+kAphHR0svqvSgDQrg0ymWD+yrnF26IiqZxDgzRqyLztsExVxul8Oy7
ph3fc3s370fX1KQRVn+v7fEiQ2hfw8ddxgdWQgmH28fx2i40b8yrZPXSQjhBcSKf
XvOrvXdyCIcFF1d1EkrL9b8jLVOT1SSM49ykiPlBd1OYOmRZuvTXtV8Y5BDGQneA
RRiqOxUdVFGEvVm5UXaawAlq5f+QTWc1RFodcm3ssSM2j4KRFhTZMNaoSRBHmDrb
fq8cWzJPpyN9WBKI0RIJsdHYkDy8fSXypulqnbufFcLgf/IvV7/kw3u27ZYDL7kx
h/ykoo1k6GC/aKhXHxbJTeI8G9BoRUgn62++Sp/FfyLxCPrjYK0Eg3f3FLb9zgIW
4Ut/VZ0lGAQOZP7To626yygeS/DdwHwUqva8oeIfdrVzm+EjEfcevaOxagXyu98k
nlnxwPviEJD7WnZ3LJVk8dExFXNGQ0swqZE0egqqzqxFQ0lkeqpcedqZFNjsQF+Y
xDzpElCeo1SwQD8JWrck5rB0FjAa3xpRU/+dlfQX13QiCGBkQ+5jsY+qij5co4sX
nvwuf6VSfnXXQjhyqzwWpbSm+egYhLp7TS6pgxHndVS3BF8hOeJyX9M0jqrGxN+o
Q0JepkNNBjkVNIYIHHKQN5nlAd9eI+ZZkbXrOaicTIPh+ps33pSqt6M5or5+2iiP
amknBpqIXaZxHWVbZTQcaNhmM2fk4GozsrrddngCjkN6ATUGJdXgUed7UE3GQVgG
/jpw0EpLOlohFmhEhAm1oMT1Ot/c4AKZLni8rdi9MDjuG6KtpdFEpChY+b7BOFlP
EQewZ5TSp8l5vRmT69tOZAN+cc9SXlhB5jo47ruMhGY+k80ZxMop1wR7zYbRU9ZO
n04o8pZzjIUU0aq/MXaiUriyXO8v4KCHNKEEGX2CQ2Hi6zSEO8u4CSPrHQpxV7Bo
7YJ1ZGcW1ZCOHaQPisWBHzsTzlREYqGjtYYKZ+S43KrKSk/NIeOhpKUefgUFRScp
AdaS6Kp+Qv6/Y7D5zG17yXo3Do4WcRA/U94oyIB8pGFOMVC8xoXkl4oIEi38/fVs
AYnsMDhz8rwV0eHL6hlg8uFUbg5ysBdm5xOuLYlUPlxmDBpiW9StLBdpZY9TttuE
vbPKN7W44mfCmx1mPKy33Sq4bJLglLaBfCezjeUO0Ar+p2nTRgUtYZRDMFbXkkkq
lINuMkWIUuCmBIBIe0jPNDgbj1Vuw7Yo8TnNocz54MPW1/l8rcwIL1TJrQxyJuIX
I/5f5cMB6NQQGcIqSxPZxVkyOuwF0XMOx9MhepyndX9cEP1qra685xso7NEkKECa
UkbZW7rwqKpjRStJnJ8zaRkyICfY1k02MDtOgf+RwjHDX3KAGMcUGVYYdJsTu6OY
mDHh5+b0jHAZz0QkAVGtF4IqYnEH9f2GvbBzznIYSX4+NbTFIbkz7GqYnnqxOdcN
1NOaq+GPqF+0eSjj5Xngll8DAL9apOeKo1cFbgq/1ZPjduXEX501bDGTdtIQdZ64
in8yyHAsD/agw3LKwmtsVFAb2b35yMfMhx6PulrACnGChQouBsH21Qn6a5Rc2PPk
I4YZd8Y2hb/MToEhKipOnkJ87iNXpOXedsrcvvQpH4Ey7nYExiWC1fI+QxFNI3W2
FmpR6XZxUds5q3KyB9bRKoeXDANVWbWdyrdhUC0tcqFrnO/8slBchAq9nxd9smNF
Va4+eyrq9lKpgh1IquNYguz5bn0TGE4H031RlVYI53K+hWcUWo3XMOshgpvXCYBy
33Tqye1gjuI9FViW2V6vq1zAIUk0ctExxW1onUtvZkXSbDonJ8SFu7so1I4TKzGe
x2WDBqB3CAR5FvOM7m4F4tUugc84b10Oh8UeAzYXzP7J5F85PW15Wh5uErgFRQ3Z
ZGVoAfYgkbYUSgZVtswBx2A+q/KGFnDjtP34B7O9+/7eVYdUndi/f8ycVIJMNvxW
7Qe3mOzqjFaCTxjoX+N2j+sdsUHWavTdquaS6bfXJ5g/1vg73K2435Jy6zN9m7Mr
SjuKKAQ3fCC46aY3l27VvsHNkMVGn+h/u+Z2Blb7NR1D90bPV5moysMmik5MvqLJ
ANj/nKIJbdOhdDWW7z0bS+Z33QEM+le0DYhG1KzhJ/tJrWygVcxvqQIMAwNhsqNU
VhSBbVImnLvoiIWf2LD8V3d0oncEhI6HL8oK6T1q7TULBBysXRypODUF8qezJj7J
POe8J5LUTGMXdQWOSKUEz19LLT4eswTpvtR3CFklTQkyk6YNmDxvmVKzIMNvM+mz
g06sZmOIdxT7qxzng34Sop2MmrRPQTioNueQmfP8qqxBdRmKLTxVOQncCIOUIEHu
FS/B53DPHuQWt6ypWj2z8tx/89eBNuP2C0fvdaVsSJ0sHStOosnxO8DQ8rLKYH6P
H0123D9Z9l2NxLJxXWOPR1vC8X99Rjxytytavo/l9uW/Ez6/1SA05k4O/EQfyCu5
PaFHQTfU0Gk0l6MU+I1MlFz2p1thuwrUb1BavNuB20TkXROxiuDeSMSk+BEzQljy
ilntBdBYAd37Wfz06tUVvq/fO+GXSMi7whiYIGu1CSsj7WW37WxIAr1jiCgch/s3
3OsIHg01YPqlYedPmVEDYY8yYGBtecL6PnxPfTv3CzYxDIbCwBNMCZV3WZRhP50K
dCo425jMb3X+zEMbA2Iixck1niPmNcLSePdx9KnLV3K4fJOcJ9wM+4klvTpeIsb8
hviJGw41bXOFl5x8IidtrThwp9D9V3z/wMynRx87W1bYFqIWZY/V/UKR0Bk8u/hc
Anqy1X8rF4di79r7+r2MgGIOc6zX38COQBAO4PtopkilVc2ibR3qtP/ro8Up9gyu
MaehITZrxgsX/Y2g2Zje0CZpcWqNY/4+2r7fwj7kXC1gpHf5NCJK/OvDoziclxbk
ku+pKQgxWsjP6fvOBIHITcLDxisF/Qk2dZL3hj/8CaFsVtwLN6vNbGg1WRJagxUB
Y6h7QsIaiBb4r6IsK1ejiCGFH2UWJ9NGmiDcX5uybNodNCQBgxtWEQosIlRp6EWh
nvbv+btmJ9tjl4HZjapC1LRziV8RArbb/GI2wR4RP7SFtCOXLG3+iwlzqZi+LGez
mG9GeVMDs4R18Ixsq9yLXe4ka84FVHQtev/9RTznB9rPVDVXRZTrYxPpnPzS8oHn
TM4LKVOPm4aghMLAeUhzNyJaiaxIFWJ27Ab29HoVCG1sHOM3SO73Rcb35mqueBdG
ZXf1wkHlebeACrz15d77Cz/sayjO5Voz5xK97OtiBQfILwt+h2p7qnPEU9fq1r46
dVc/W4clTFVDo3Vc9qJD+ew5ljutTNqu+WZRGOgcUy1ta1k77xvCOqNtruFiadFb
NRMj4pASuS1WuYul1uuvm6i1rDezftBN+ft4Wu2uEBUj9kmFT90B/VuGIk4lwgdb
uwhVCXvrjAhR7mHRVGNOd0d5OUI/nOH2Q6H/+EriiczrZWCAvgAdICUXLX/W7rpM
ESGDQjhoq8J6g/jDxALKWyRE7Iy6Yh89HJQCR0fO+q0oqhtdNvWGaDvJlH4mK/DF
mTqRygSG71IdFckjhz2PhztW+xzlUnwG0+XIpjhSD9OthV15g4uVRYpVY1TIQCdI
n1IWUK3uL+89A03Q2SfQf4EOjsfJkvGhZ+DRcD4n869z8axYNUtSIrWWeMBtn7u3
GB/hzKxDIe6OLGUqMM1yKk8vYcyu8ssYG8qcD53sLUvopxnaG9AMDRp0lJt7n2Ms
NrQDdBLgyJGGsgzRrM+ZkTU02eRxRZmVhUtLIV03OxxeRkp3/9eXaGgUCXxk+tnC
rLJ7Y5RaeT3mNPvNghg/3eUJ1t+YRdDwvDgkoQ5A2t/N6qp59I1Wk6D2QW+jnHQw
5lMl/w7Bj6Wqhr9kJYv05AGEARob0N1LXKW+YuRdQi6Lm9D73jU4CalA2D0k1ado
PKl+2HbgPgH8SeSD994b90H3fv0kmkXHxhX1y+kVsRNvfOWGk+5Xm+jgzxC1v7lz
X8BJHeVDyAqfO0tfCzLRfsPgd77IW0WblzrnCXmq5pdXqow+IvtkeVZ1Mzirscss
5/3LBBNIbMxQRx4hygramTqNXEanrN7Qi0GfE8G0QTx3iuWvgf3jvc2PE60jrWEb
3j0yUF95aVge/t4/igN6odbc54hImRpj2zgYYgGOhEIWgnC9TOAkNvu+J1VQoj8T
+ONhcfk6ap91oDBxPrq7Sg6aCG69Z7QzIiOUTsChKfb5G2lduWJtKxpVKbo2J9Ds
Zd+aBkjtKnze4Ol7WUh85X6Zxt/WCtVIOK+OT36BJrkMX+cGViLydfa1w8O2Yy0/
CdW1zjuOixrSJwUm0bA0l7lbh/6mY1RJxBy8fmO6LdshcDIADr8yBfnVb2y2IDIX
ZihnGaIot86kXifldR6neUZOTuIB2oto64gaSij7MIPZGQd/mer0acKxru+D8e6W
ZHJ2aA9DJISZeiol0+VOWu/O0Y5n6AARJk6ArF5QozEdYqpS0eOXj5UytyBbWTAi
bg3wONToQd9cVq8wffFyUsynxhH3MI7SrbDIvf8ekzvllwh7nZjXb/yRb0q7SpKI
qQEJqgqk9JPvxtrg/6JENwSoLlSecB/+d6WbvDD8gNOmz1oM9sL/I3JVqNN/jw44
hrWfRFoBlh6zhB3Nn9J+WuBVjVTYLFPQDG3v0C1DxIC4N2uMEzmHOFByzRt64vwH
sVm1aXFywOqELJGIpRfpyxgx/YOFaYXQ8ML1edPomASa3tJbY5SMMu7aWe9y8bdo
czUl76G6LlSq8yz/pbo37OFrRrGRvslgsYdXl7hbswIG7j4XghESJM23l/c4HTuo
JbHcOGeF1VAUG1yXtQDP/volFCy9+ZVHtVnnDMQWwujPmwGa7n3A7XctzuMY0VrY
pNTVDMD26NiUhC3Rf3sjJMcNNsy35cpQZv1qgepnFvYf8FdtuNqjMkLzvdng2MgF
5mH7saisHn06s/vYzfBXgPQezdUrBn3e1zjTSc7EOI6Fm7JK3+fTHwN2x6lY8ilI
rz5ZYqQhQHA+Qxs4hZULkKWf40RgNCQpl4WOnAierukEJW7wdpZFRn7WwtUO4CyR
QIKCmQZsDdv/FEArJWLVmq7raXuv+tT8nfXQOhGoRl3TKdZQgsMnORhtvpIk5Fry
SqG6x2WOuy3rbrZXZuyH4UBqKxBNYX7kjKliCtsbe1i0Mk7fP66Qar9jbj/lcwdn
/3wUD5AJB/iLgI7484g+RN8zhY71gNpBQJnGOS43JSLIDkrO9WLj6VPQrQ+YO2z7
3DZqq2Kw0Sx5jPYW1qUt0leTgkCtDFJCEtdmzhhu6Z/lIcPhoeMYMzSQr44EE3zy
Y8cQD5JLN55moNSnaXX95VtUoCc+2Ho44gyozaZmIqX6OAwC3xAfyTih4v7aM4cy
u9vQ0a171M7i/U4qB5nwksqCWeGBurAx6QodusW78c71DH6WgZQhYStdQY6s0WcV
bcO0tRZ9OrJVuRRuXsrg7mbnNjdVNQmqFeV3neZbli9ucRyWpSPszV5abQIIys36
AS7oH3xRheM7sNg+Z+RKg9HsloXzPSIQcen3Wi6UCdzkTCJZBAXXEZS1w+90zk/o
qud7mCOCVUpg8dLa5e4ow5JqS+tS+rgBJS79osLIMj+ORSQ2oZPIFkssIdL4gyRa
pM+3uWr2iGcF27FrIjvhhsHFN69upZsBZHZjXdFcvVT8oHmhDxCtyCzqH9/MsUmq
C92JovtIE99pHVeziu5i2hgZoUjq7wxd4sQTrrCRchsFFARuVqIBAf9TvuaNVQ/z
1ciuM/DB2eD/39+HdhO5hMioMJYIjSYUQzLCOyhKImXQuZp8mq2TUjm+Q6eNkUlh
4k3if69EKP8wN9uVVLEA9/dI9RDRAWSv0HSy95iqb0p0E7AFFj3RNJFaUTzIBWNI
A1S2SdTJtgU16JTPn7kv32crWdBYTR0UyVsi20JxP7ySUs9vO2JOCpi8oOwT1M6R
c9ERJa0m7yWdjb3WKPSBMZLmFTD1y81zh8CXd7+GODtA6lZVzshrRIaMZ+8blSJk
3tFUoY7ydXmJ8KGzlx0rK1REjDnJcuBWyMEH4IKPBy4GeF8XKxTCRMRL+u/v4w1j
xXbc8zBpCKxZsUtUHjW9BF6mGxKOeB9eYx3GtHf44i5N0hniuZSOnilTiYfdRuOB
WZvi4eJ5Zd+xMEoEWN6Vs/c4RPRIcvTAoza6eqe0JxheHDCrkxcpb/PBQ//OoXiM
ZgnEBoWP2Iwk8VcmrGg0hJ4ID1y51LZ2c1AaZQXzwFfh6JFuRXVXvB4J0mfW4+s4
19Wx1c8isYDJG/LU5paRQL+98mNJUgs0KupSh6sWksleHi3mtJH6oow7RreOPoyY
3iGkGyTTBgeYa8WpnywaDcH1KQYilb4o6t1KyqzLTD57bhF8Tmvvmvs4hK+lCaSZ
vTVjPfSjhPz0mbp91CHcRBUGU47Ld8ivF6wgzbocJ6+UQXOH3prqJpFtCpvcVbnt
hMWpZVwR4t24Ccc7iIs29SB3iDaz1Q5138HeHeaGzTeyShrqnpuqbLyt88OHnB5Q
SV3uI+tdE2ed/YfvXOflYyN5GbtazzTBQvyJtmdwKoxvGrSFglkZp2XqrloqSnZ9
pTVJzMvs5Ipc0kn/JZCUw9cPi2ybiCKQlDUS78HjHPizrTXDyj/Vb3Hqcec2SQhh
m4LRGDif+DxQft4355UnFSlBhSlOHMNNxO6ijBrJDkXOdXL4FLuI6RS8OWR+6R7l
KwZsQpQ54jC4XVK5sVIwBqL3BHPG7dvzTK8WLatlaFulfr6YJ9N9tsx+ibgQz1X/
Pz+xeAYkfkjsYwcx3NH4Jlb50S/7qseTv8vV+YeK/MH2/o/TTPTlqCFU0EiU6cEL
CsF12/0uUZyr68eZoUSL3w+Jd+6tN/RjwajygUVi55JNV6xt4bi6REg0Uz30A765
2rK3WccSD3Z3wDzq9rLIejy12Ih7oY7j7Ka2cZSg0nnY4WdOrepamZ7NgW1Q+Ryy
C3M778Dl4pMBqNKYEizRtftp2+6VIeIbR46w6qFC68eeTiLsb+XufILu2Ujj5fY+
aXBP7yCqrVP8RJt5326xZw8/PYb4+wWRJdVwK7BkVAjLScV8QXwEnXWhSFsSjlg9
ZfOhYxIqBYekb0os00SZSd7OCeLpmOOZY5Wk9LfpJZDQbtJfID78EBKyyN///JjU
evMft7xoeVp9sH4oROtgRZcYNrJdYEeRDi3Wyd56oACvXdASnF9flOsds0QZ+5MZ
iTYncRuDh/j/5hIlzhFJrTroQVHRYXgMi3n0mI3MjTra0Ks7O/FlQMS4pNMjgGlk
qeCnMczlalyaN65vNlWr4LwchVAauOo1rHI+JoiL1TA+ZARY0YFdMtwFYKNsrYfn
E8wWGkzQvt9y3CvNLrcz572Sd7x1IbHXKZ/c7OsZ5rC86X3Yj1Jfci/eVRR9Lzs9
kssdJqJNMMs0gwQgDix1qtckK6w0FGpc9hKe1m7cpjGAWZH8aGMFdsSXabTZCpa4
aQx4AInyL9aec/1J7eCLyYJx69pe89JE24kbp7c5uJ841evG59Qj58lDAfIeLgCR
55t+A27bI8+wNDEQY7u9ULHCGvZBA5aYJ9rWdveRD0kzmqK4B/v98+Bu5S/q0E8x
FgaLtfq4gY4djHeK4LR64Du9HVpfb411l+SPd8odXMQuIlvFznNkpZfpkj5RP5jl
JLMuqlRZps6BDh/yCWqOadUxknQQujAxiZzTnleARi2bzgsx7ejV1XcrKZ8NWN0+
PVPXsDyLq1ALZbn0NjGECGSGD17s9/vP9G5sRD7uR+l/ECRS4Oh5IyLYXGPr1u4/
rDxzIORcMStLA5t40lSI4nRggEcsUFn620thjifeW2OFqSZzsZv3FU2GcJG5UTLU
AMPs/adfqQcXGhBWOCQ+c0pGELxPJDyXjlWASkfG3Ut3n5PonNahdL7/6TtgaiOh
VEyM/BFau3ROqlPUctHBcdlc9QCEmikxGNagoxt7KIfRUbV9Lmq8zNSP+dE+ZEZg
iNjBXy/7eg9X35PrLncHBNKmqnX6kz9GGRXX/dnYxc1RINGP+vc86wxiTHXSNi/+
br2OrBzA9F73/C2ch4z9ikGfVkXYUBNkkWJ+4AF+4P1KwHvs8zTmBxGazhr+Qb8X
q/iBzNvZsauXNi2zzVRuicOd5i+ZaNo6rhI9qzY/qqYiBg6un6LFvzFIUiYl3uUd
MGIyZvGtXXlCTyHz4Xk1K86bbVTxJP6wHRphJn+W16vfLt7iR168V+0VeMI4ndLs
ZqKUvpwhq+JAU9uLRd+Lu6OzQQY7f2C4TfOZW/Z4aYxiIcJGjkh9sGnCDapkfVS0
p0r/srgkNJaX5uZM08QCwjICg1cU5Sb9HtaI3P7aTFFp1dL4/xc/v916XDAPaLSb
D/aCivfrzxeVI+SvB3/wlceN2Wprcag3sntsAmaWyU2JMIXPvlsF4Tr9SCbaHD5T
KNeiGvAqKwcmgVX03vgxncoGAV7QKDzF7jSMs+4B16qSUh1BN6z2CGXKcj9Qnuhi
bEx2pswbvDLMRET95DpUPnnLrTwCRtGG+8FgpwKuZDrAywPfWHP8RDNZGNmcAnvS
s8m9wI7tKxXXiKvSy6nAkX2/8KOIaZlhLxbcLsfJrAOjhRPKHuduujrxTA2nwEZh
qM1SzDpovy34shVLVHgitPtWR4HUpya6kS37lexQ/uNx1HXEYTWRSJfsu+oq24Yx
prHiWfnyGQ13ZiuxN2EaaUQIYqIPwRvAcxAmvQbUDohOo/Xb1HFrVAEa8z34PLCp
Tcj4dPoaeCrSPZSZTCZF3chukJuL+ae87BzSzGpWq1IKPVxTNa7IUYvTMkzkA3Z9
n0BTWDS6ElD8RBlzDWnGjKbTCuL3FuyFD8h5Jt3v9sA5f3nuPKyU0SA5w93PVMYR
QlsuXqtmim/33VOSpTCdSM+f4+Uk/ueGPi5JNXTYsfoyK6Oa2zJGHtPMMWNvPhWX
aAWL/cdmcrRgOjpXdxE5DVs0iOe3ya9DjheRGU7AWhkM4IsJepdRNwhjVf+YM5zV
L5R5nF40EQ7KdId/uv8u1j6BYcbcCYODtVX/AA0TRWL0pi+OcjLUQTHi3+MD3/pW
RsmE1ca20s+4ymmMzyfEA79/JcL1OpVMhTKITBWHiXtvnmePkJ9EAPgk53pW1TRz
LV2m2w+/bGZjigaLtXlh6jLbf7Jr1c5aPvTIgpd4ix4=
`pragma protect end_protected
