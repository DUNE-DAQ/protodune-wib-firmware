// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TLe0f6PX1av9+HT2kGwfTAx4w57X0GDDtEWbyH4jAueyMmNWwppE30zUjz3k3ziA
n5LX52i5fR4olW987ZJcRey9Rs4HRoF7pQdLpG2wXcv8aQcvLHal6fiQURtfEqKF
5byvW0uAufFPkp0+T++iO2QEVWAeeTxRx04K7kgwqOg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 174144)
gaATEWtq67SLBemz/MWD+z36u/uSaAJ+vo2ugtQXZfiNlYPcptsK25ZyBsVaCWTN
IfEwFch3qgb/1mEpR0kSFbTxkNWj67iEoEVu8n1k8Ti2IbDwbBSThtXJ4PxF5Dls
37GEP7eMf2EW8Y2mdVye54XavFRM3hWQ/ELwHE5OR9hJCd8wvFBamO1rNWPNldd/
MkgzWVRM2rYv3gu9cxdIaf5r7XXIvSPokNfIF29vxBfwiVIiBIIzk9TeWquItzdG
BoAza4JS2AWGlEihtiMZ89mG3l4Wed5muxQlKOQaPId8cXHMJj9NDlWUj4bRI6mL
xLcIgBLzTHdchlqJvqb9aWlSrVFb2GD9AC2zyNjMuAa9PFsSrGTbtvCOGFN0Q6Bv
JTa7gE2grRdKHHghAZCzIQ0QQRLDpRKadTlFzKOGwRqtuCi/Jjwrl8dYuo/0QrXC
PsTVCSILW36PgiM99NNhoZHIO929fd69C5MH0RrNANhWp111lc7CX5w8V2Lp+Mr2
xM8DWOxRf/wLtp6u5czddwp976sGg7i8W78G1kzqZ/3X/IJ1Zemvbx5OgbGGYlPA
smr5WNA85VY+tTOTUY5HE4g6mCmCI4FGWdi6IstTV4lpTwkMs4lBHehLy3cg7x/y
O3dQRkLIhQuNGT3NvqlZeNowvjXjtO1tb7f69ZH1FjVW1XuKrgE+CVIqdQUCDqo9
EIWw5GxjwuOxW6GphMRycbXibfxsv6cgPf/mrcJWG3mDg4JsndvMAuhscnV1pG4n
nqEDiQkvvmz2iRJisvwskjrxcOu+KNOUbS1PN+GnWk0W9en94gZT49lHXdqhIRxP
xNEWkPqsS1PdSHDyOw5pM8RH9c93wc5Zjf5zCoS8myFm0CAUsjp12HqlmCD3/cZW
YSMMkcppOjyYwbrNbt6uwScvel8uTKIwOYoCugWHGMWOYtPPX+tEk/X728Tt1/5D
ZtLECHt7VIhFu3yLSl9jlhMOcvPaRiP6vhQ87gKG5ybcy1zJ4eB1+EJJ8DbQ8uZ7
vIm4ltutI7M0UyjRxCZtDIEkR3GKNg9VLc/JwRa9QOn8M/jPM96UJnXBdj/NPw++
7FMh85OAFFX0QPXXuwN8eQorB44sSVfgubIR25WewGsXfw+KXYnrduTuj6POZDvC
QH5Cr9w60arG47jWG4JE+l3Z6W4n4wZ/s6YDs0TfKRntyMeok1GKKlssbEQuh+z6
BK5GlluZgP4ESbddfWuw89BZhR7kwOGkxuJJzygGKqaUuQvO6PBEHll6JOy/uWIF
uXrjkWk/4BPR1YI7Ups9G3Ape/ToCf7sKs8YY3YvsnQ37LjkXVWy2SQ5LXzvfrID
LRLuK9Fxz+AAeNxCwDmrWiLGWemFYhoxrbx9gnrnfP/aNUvpB8fyqPXH+EOJsK59
fjue8Umz2Ot5Aihodbvlty8ilwE9Yx0F9AHHbHYiL2b8QEZ44QumK3HbJ2gdXxly
vM3UZERravf9FXANvbCx+VewvIi16Ii0/53BSTkct1hGN/3Qba6+DeOB7U0yNCe6
EmuOrW8HNdlVkgE2rJqzqK4nZRuPx7mvBLw/WO/oDaX123iXUERKXNM9v4L2HZ2l
IDRCnenl6ADLexR1yp3szmoqTrJ8NZW8TPTurSTwR0PgmuXkBwiBJxL1+2Mf5xQt
EKFku6wxOnRjgGLYCMph/8aJNUT9ixVwEnwleiL6Hlg5bwY/SPEgCRRSYofaTZRq
ieKjSUZyG9/rq2L65Uv+PsIKTrz5k41BsL0LgDXctXrIW/V8BfDtsktX7uGOJk+T
48eg4GOh6TzxolE2/MpDl4jsvUi9YymXhUK9A7vU4VVikS8yGoVSmXqbQVtzFkrv
nz3ZzdXForT5lrEk4oAe6hWQ1LfO0Ab7dngCyUPbVeWdhr2SXao3Nd1qbcURCX/o
T4IBhOVsOgXyOrrFi/V1q2ZRFVSQp8ABx/NOEEQdGAOw4P6N9Ez6UxJw+scGaRQ7
ujcZDdSMAeWQ1hhWa8Rqn5JYVCVrD0UqP7NW7j4Cgt0iXqkyYFswV09hi7UGJgUI
Ems7UY5lE6owpYr9CFJRopqdEGnXApE/MlzQWyToukuGa4DnGf4NsDHjlu2PqKKS
Kfa5c2FVmbdhX4N5aYv7fw334o45VAP/Yj1a9xBRmUzL82y5uRnpQEQL8yH6S+ox
oQ2IakSCSIQirq9tjbl2GpwyQwK4zFC8ZI9HLuvC93dBoTAWwUkwvZ7SlGcwNb3J
9beIs3kNHCFLAnUMULS4Th+Mcgl0gfNShrgSzAcDa8gpIY9jvb84blaOFBRgUf5L
bI/J6bdvIwb83ZdP22SgYKNnVLD4blvcYCea7d41wqoYEo74eLNcutqPb5jwN6p2
tH2yLSYpfLa/t8q5zHud6vAKddLC45bA+4YrcQHvteNw6wNckxPD6+XLT+dwSJqd
9JSRjunogeLdXuucto/WZ/wyB/KHYxl/0O+xzVM9wNbHAHx071iit+Nv6CMBuv4K
DOoJ5RnPF9vxCnLLWSD1rdCDizXG/+m4j7CD3PsaZb1Bo7xlDcUTASSHgTlGCJ65
IxOH4uhpslGPMrS6EjlgJRL2s1kC+JTewUls1zrFzPVM6OnBep/yhmNPb2BGjkjY
AcHArLWvXJn4w3tUpmDxeJS2OcC0B6cYQ2V326q8jqncnoE9KMz3JgpcgK/ndDwo
GrQ++KZnLCw86Vr27Ufgui7ERqnX6Lvo6GcNKJEa3+PcY0gvMOWZpbt5DHhxu5x2
yd6mYTibz47RlC8S3PogtDHwEvw76eJ1aL6MzIUp2Wv2DlViuvUOivdiWx6ZKpCl
0JFNSvg+1zf/6BjXOxRTOxkh3UCq2m5J1mv2UfWQiQfWSRShkL8XWgm60TAi9fTM
VTSd2tVEpUVWofdKEtoJ0BStbL5l/MD/rBHrIUrKYeJiLT31BjYoEMWIdKCnetd7
uaIEgHC/6ciuhvFoAY7TmfReWPuziMwa2qphGlvv1PwpEIAG4jwR0hgZptBpxCV1
D9w4JF5xP2UYNM7iOqLb65qB79LZCJHfoGfk310w0hT7giDnvz3alKa1T64/cX4Q
o5RnAbcmsaWnBz7n+wnGRQEfAb+ZdfG3OLwmoEe5ulJmxBWkZ8G2NB6KTLwfD1S3
+NqUDd/x5vGT1NMQxJMSEbdfqAEUqs+iUtKznJXslXQqau32iMc4EWa8rEEbqB9y
p0sn95KtFQIaMK7F/8VR7wgcHVp443b7ANJsKlmSSgVjQjUialqXwJJmn946M6Jc
lUPmg43hdN7yooTVHfTwGzxDKUjZ/L+hgTMoahMJUvFDegh7M7URKs/SK8X4koO5
HKMJJ4jDW/yjL+VmlSOQkzXCXZKYDJUTH/+b4iFgM1KTI4Jo7GPLxvb6gQohQ6t8
Jt8VzPmzP4fUa06/Mb/RN/fqpr42n9/VS1SVabOdYUFhH0HDeMLmwn3a9V+Dwamx
Fz5E4dQHt5Gc+FO9hQJJKJHfOc4HYFnB+9Oo8yN9xdcpyGgYjvDYJ4Jp8HPVZ2QT
/05N59t0TsbkA59VEQgHvabEGMDjYravEsNEyzu3vEIrlXnfSEVuVJ6yVM6tVLJ5
pV9z0QUW/Ao0Xyp3KB6jz5PGSlghWDfyc5+tN89K90BtnIk4GNl8VX/Eyv21W5LA
9lr9cBPonvZnNa+EMDo+aJ3F5Fw8UXMMyoG9oOR7U5uLFhDCA6nMCyq0dIM0Ok6f
Sjud7OWiFYFzB5d3VintfLaK0RmAlJhY4ubLOyPXyR3d85Y8wv8SlCVcBQB5MzOp
Pz/osHDzsF5HSiDNJNna8eYBWzBmLP4Cq6zhN6ZX6JR5eKSysu3g3r0audg19nui
bHrkPYmPlN5H5yTinqzE4JkmLO/SVs88LsVIACNjFvCnEYyzPdDc3JpC/w00UeD3
FYeavuRSheEFH6roZHyyFwyZPWyY5v/KPFTyKTmwo+cW4PGNdQvj9T51WTml3XTf
562oV4fmUvFVM+B3XH6fsSlqBNbqkDfcCfKo8ppFZ7bwepGj+WFFrbDfeUkDsbSo
iWKQGGgmN6eGAdXpxKRyZKUdbZKlHyI3gjtOhBO0qpqyHHxQCRAqn1cch8V86nrG
mzLxC/vZATuknPQIaPByQXjJLlQYja4bqx2QbrdRu0/CwVdUMIOOf4R7a0Dnx816
srHfSL0gIN/hLUdqPmuj+j/fdnccIaXU9JPxUeQWCC1uupE6CMLWYq9ZKF5gsSfc
zLUaxIDuMO/qC2z24SxDOs3p7aqC3aQtfoIBlUX7MaA47IMTvVCWc4gkohG/MDVA
+63GH1isb7FU3nVBIJ1ObhuN4b31mSzSa7CbBVgegKDIWpEep3chtRmIJMvyTcdv
vE8bIVGCZVAC/jYruyjdSK24PgMENBj5JeHW4e7kidh4sKN+xdTV+z43pD1Rcihu
fQ4fKCJ7bmUSiJfBHIdn7erwJ87ZipMjoKqbyymRV4gJs49YwrOsosk2dALPMFqE
p2i4ym8jbWFsE7fOOG81xRB8ZmYqYQqBLDjlWiN1A1AlJBUtcjMuv0URTOSih3YO
bS36eil4ZZ08HkdZSnjfMbMz2EbD4jcq/DG77Dwppb+/4EAn++BXMw5EtBj+bwpc
pRMCAymthvFXF+hSzy5PmQ5j2oB2fIAksuj7Sa5Rr75x6GP3ScsQ5PhrzKTfO/yo
SbtH3XQ0xqLlvu1kPmvIK+GQVAB1XZnB11jC6cdkOVaawTVbWVTzj3whJ7XmNej8
JMopWCq/LLGv/SUawXmz9KCf6IxI1r1YokJbE6ICiQ+7qIFAJmH7iu0l6OHmC/r9
ICdzRvEIsXS8TtLROqhGvXjqOCBTDNuKPHg/O6JCj+TLI4UtEg4YgbcSBIt7Vhp6
zeUA1jhVjyjrVvtcU8LPf1GLJCbqmnnq2KfwUwIhxv6neUkfZy8JobkPwPCntb8k
S5eVznBEo5PSDPEAq/X6ARcM79uu098KorMRxxDyKHwTfhBrEklf1x1lh1yBYOZd
xyPHWCs1RDQKHEzX2nIOWOBCAWykxycrV58YNLRRoT+2Kat891F63aJRa2vEg4hM
0imVvuCuqg3YoZ3LIBq+/enN1/vCrujsyMpC202J49guYqSGqUVK5qc03dNAS0TC
/IoZoSoLmGTmJpUiYekDQ5vCkOZPzHWari/tHM4MvUfSO0ZL/w85LaJhYp7craOH
NOsjcZ9sVfiwB+5nm//YcTY20JjlHfoB6x6zkg4W1mhjMnG7DZoNFnWw/8D8dSQ8
cSGKcBGaC60DjH7IMD7Wn9XuBPgwanrIhfZLyyG1VoRhxVM1ebYyQYU9dbK3sFDK
53lRxIKe79R7Q+jzh0yQX5zJBowhscMbHtFd55UE6UgD94TZXDc457KVtev6Qrzd
tKClkge15eLDxWFS+XzxCItQYKDSQrS3NTMbxQNo01DsrRpadhFfnTTnuI43nQoX
X+pxG71yY7N9plovm6cGvry5VOyjoBEbveuLp0giPXhMkdcKw0UiCeA2VIXEBoXx
kYmymc/IXJ7c5mJQyf2AwOdhft83OEC2a9riopsrVHmeQbhKGk84CcgtIFqVKZU5
FIuKvb8zIvvzDOPYiEU3KEbYJXfkS2fRVpI4XDxBxdnU5yDb+XQDI+HC9njEbI82
AC1z03e7zcng5Rj6oxCkXeygOLonSSOtq7KwgvhdypmLci+aUAvoaq6kdXonFmBd
TkgpyfPW1bKEIpmlx6HLIYeeiCB7XPssrdsVXBDs3jUDrNbZ6bC3Z9cgLNr1hx8v
YfBwugFa4NqnJoCl2z5mQOsQGzcpcmU0eo0SpU3esW+evYxZCoreHC70L0QQ+T9i
av1LWKpU6/ZVOt84cwIpRn2EGjYnIgkRi1/UcSFyAwRQazBAa8K3t+6nf+uFOdbX
vE2heF6GL/RYyKiCCUIBv1u7+lw2hABI7gUC1Y9TR7xMAxXeO1bLp05S5kGWdVrW
l1LaQ7T75dwe5e1a4COPClgZP+svp+b6xNnvy4uCQkJp8AtKCVey5G7WpfEFmkCp
VFIqv+TtANIEC/BLe94GvHSwTmcXW3mgRQKhFJ0YbqBBKBR0f7BYvybJ6lUKWrD7
AlB7SisFrnDWt2Djl9K3gBOZV8ORI8+rjBo/YvV1IoiePIfOl1ZO4G6i8O4uBgsZ
fnO8OpzA7nJ8zgLL4M/ljo3U/EXMcne7dBsnlc9Cu5DUGTmjBeSTN2wwC+Ixweri
vDxcxeMjrVQq09upZNlvrBymtp3Wma/f0khUUEBtfl8M4Olnm+i0GV9Gp1E02BDy
+KA/5Q4f3Yb4ludUmRbSzV6VNHFYsqrYphsqsgd6QsrNT7jNHht2HFc6k9v10NO2
Nyni2EDqXcwLC0HvffxsxvtOMPswRzeRQFHo24rSJj0Iz4OG3LF/F1JwF5uvUSHc
KoWX8tZ2Sm5n4BwggPurSemL60YinsLWe+rBE6dkbcQstl27IVDI8cFY0WhMpd4f
BrGSc0YbrPR6J5cs3W96IPNrd24SUIfbyJCApemt0CNlP3Fo/FkXvAolluiVFS0m
E5+Ri/bJgzFX9sHmHz8TZWhWnkrolSfw0T0VrRUdchW7ZFU0gUoyVheJd0hd4Roi
L6QRzgBH1CH+l0QOOf2zdajMkMX5zClJl643ZXC3khv8Hbb4ZRfEIeewIyGn0hgW
5dCHVegFaH7FAtCBajDKjgFBQa/7skvWsT3pcBIKkyNlLl9ZNvgDjjWY7/AowQjn
pvQ5OW/GrZXYrzdMFHzbRgcUJObkZl+9Zoxw8C5BIJ78JAP5Rey+faBuovOqrA91
4xw4KqpokdL7b3gIO/PkCAfN4MovuCjCg14aBGHnVlLl7Co3pBArgFzbdtWFnuZa
l+c725Z0YmYRF07zsLUj+Q9ZfvQjlLP66v5SmJHMndbwQsinknbmYKK/PBXL7HSb
4vr+/TfqeXqlgEzD1aGIPDU6WIKoc5hlE106BzDwyRz7lGSFDIeYCWChNkkS1ZVu
zD1uzUVwnTyqlIB9wbHz6r/O/Zaq8vOwMG0/KO7+jQj9mekYQ/jxCvd0KVMbrM4c
SyG+9SRwrJDZu0hFnQfglIPBoHaTsGAVNQYHbWyMPFWCNaYzbsJ2mgOTDMQsIQOS
GnlA3PadY/Bn4E8zuG9C2iyJp6/TLhR/ARiKpKL+/7hNUqq4fr6eA8ho2KFA/Ib7
yKzMtlT0eNviAOKfNTZGNGu2m1su6uyGtU2PGSGg9XEAKuip064B07N9GFGAfi8C
UjoBViyV8waUK/TLY2S0UuPuDU1qGnNbTokHsZ7f6thQq18N2fVVbJqgMHlfu95T
FC6yLliMDvMeLGz4OvZ4t956JD9cNeKWddh87u2DKzw8IfB9WCHfcVjt3flCDeDP
4FU9GLsVTkaMqbmeKPf9w8r1Qz2v9c/EkHV01oVuiGjjG+VaxjQDEC0V1m7zybA4
h+MqaARp3MsGoeyML/i5FYIf9eLhoDSSlPO+mnfwxPWhoQuuByAX4IxLGbYF0dVW
vANeJ+LICZhpUY/TjxzJ/YfYRPKROUs4PXjURat7H/MlLHALB/PZpsR6xi3Y2UkX
hwtLIsyExec6b6pZlr+GIDGgArSZa7U8UZ2TDDcuIuw3jXpFP3QxY1Yfy+5ztMbi
/Hc/4TGv923g97y8F/e5u75cgsck1wjTm/oj+qGjfOkcgWIB++YT5ZoXb8Hs1Dya
m/3iSQQTK/mauzXHNvKhcsQdb0GLyfUcsLuwdR98jpZpQejQICb36mIEmsoyCYMD
90g2aHfNiiJzhN/UXvJpYxbD5ocSrmXucYyxXwdHqyI24SUjsvVjPuw80oyLpTgx
IkGo4F7RXwlmhnBAX/8jMVOw/5uVLy8cb0toEEj7NeCXrY6+DwR0ApS6wRmaT+VP
uuO4a+MQU8bN6Lh5NyzgYI255HnO6U7fAAgPk+SuVOfRRK2g5Y1C071epjTr74hC
G4LWmcAYvWjSlkLeo5mKhQuQvjn4x7FMIwiOfxYqOYxgIM7MCBIqAfVDvmK66Q4E
qu5/P5sayL58a3Oevn1qv4C/DeA41LLjWxppfZiZNv0H05vdmGS0WiForFrfdZEf
HXOW22XwlDeyCaxNnRTpt6DYvV+S24Tx4y1EwQnYkoC5RTtyGTO/zXS1JC9EOxUf
sQfZlHj9sbakoo+yxquHEyi5tmgReOlfW7WZ20sAuMiLeoSFESb98iYLxfNjA7p9
Cmq5sX6rfvvXo0eim8qIBHuK4pkYmw20jARU//w4X6CN1V2qbwG8/MzbfOYN/zHx
dn6qWRGk1wuGokHUMhtbuZ9ZiO3tuw40fG3RXYUKIeKbQ1sQeHrXOtez6Qj5SF/x
jg7x8RS3otQsDtwwPoVdlGXyRFoDb1SkijUlzasmCJ/Pjd6J+jv674p+hr1zAVvX
tUI+LKF2CPwZsN7gPZkqjphUU6CY4dYqpIJ5fWOjSQfX/PA8E4wz47elKqPnHG+A
t2GABT8i7EPXhSjpF4N8/ELojE9E4FDEUs2mswqH/eavTLbhV/pugCRxZQK1g/dx
g2KR3DRoSuu2Cpq+DwXZflubAUF8pnXJm+6ZKwEZogzSJvmPFLLXTEajJ+q2r2cn
YE1ajKDzP51MJOERU27IctWdgkJOZKiZ7zAHhZVcloW2HjUCGWqJU2nXt7ft3eoh
EDxtvuj4Olw8HpaWQmIt//m1oWypnAaWPVoz+xT4wyKHpk6cHh281tKBSecsfyPB
/gKb3iAzqeJoBszG2f88hpAbQYuYorg/NEC8QTNMRPSPdMcb8RSHMBqX+HZ9sRmN
hKZ2+W4dcMkOoVs22/qTKFrjBfVYudyGg2xdrlYTlc5iqrKNgsjds59u0B7U5mqZ
eM56x6OTmMwgQcNujOcOU+17XdJJJiKIEh1FnKCGjaFT2ZY4f8+HQ+NRFMp+UKGc
VIUsYRGss3/4HsUoIaDEXVvJ+V4dVipeKoFylHbiMLgIcHnGNw3QYm0vLkVGuTDc
bb4m+lL4S8++7kuNOns0Om6vZtvySRf1Njo76j9cSq74JHI4PGHkfuE/SRHa9E+D
ssukdLww9a+jGKfGX5nXYShc9TSK/mLwEVQ/v4Sy85rNgeZdYqYpEZAzDWdbrGOe
kEGjy9+XJJoQ2+DlWtwYB82Lkvy00aezsIDuyZ04NCZgZw+gxTHAW9swa2jqreai
XOvyqXB15Hh8tADEpM2VQ8dlWN6xfU5R/6hOGRZdzhi7YNoAkPg+I+ul5GHfKA/r
evapSaweeygEuktyiMCWfgQk8v/96tnQdbdUTme1SrwZmlz71A++Ci6e1s/rs7yc
6Kdq8NrrD1IeLuBL4SnNmO/FGpFlIWoam+LurGpjAWbucujDk0DoFvUCjkQJT80K
bRXiJ/KB7RVEMP9+CBNU0SkpuqSfJNyalEFKhcE4I2ocWdKcV4wJicfVRbkG1fGF
+DZe6JwCqvSdHyxzHBqEHOW5XEQUwhy/gXLHjwobkJorTAXiYDNej1AiomeAfnjj
ZWnBuuT1VSR2TPWQbfhFBTqjNsdUOD66T+u8hbpdXJ7Bwg1Ndc35om8iSADCBhVy
qj+Gj2LFuR9whe9RjVX7BiDmzVGMoR8P93KN0H2mi60n92c783Xcn8UT5CiYP8Uf
T7GN7PQnTBYmLDeLPG1pAyPFdHmcXgGFf37Jpkd05BN9D/DDOeqYUaEsQTjz1khL
LcHZQV7qy8bG5+z12v1xRJVCpIXaDaXJXqhR8c6PF70Q+eVJxTZPkXPISh1xApqY
DFmaiALoIcA/qYF9l39c506pSSl8CWTgJXQTTHTHNeohqafnW6Ij1Xfatzs/c6Ae
CPDfeB4h6qYURhoewuA0v4c/Mz2yhH/TG1peT7uYbdk3uRKbltKiddDMSbFYqZ16
C1jh+TOqTot4iiUIG12vf4ZkRXEJXaoSNhBDi+xofupkjzS5Ykz1UNMWChfXP2qI
tnHgVv6Xw+VMlQTcGIirA81/wCFU4VvU24rzf5G2cLCy/n2rbvs35yNNyibBdB/T
S9kb+dAN1G996sxpbsmYG8co0y3TqgU4HurUedDVjB/exY4WJO1eyJm5Jm+Mf4m4
RWZByleaS+xu6mEy/H9E6/D0lT28zwCut4nYZciM4fbVNE3fQuEn2OznB7SMZqZM
ZrE1QOXbkPY3L5oxyl6xgmGXz+NcIuYyzwtvTWCGZItDrmKWQamrW5yAt7139jHv
Ckl3lPD9ErJmZO/zEnM9rGYTE90VfmzSPVsttovBQRF7PoeDfk3H9yd+3PpHRXrj
WhdwyO8l8rsG6uKTMp+taWZC/ndba9ccr7rwdu2oN4f46mVInWJdfw6fniLnH6WC
FDCcEAda3Fi8vnkg+H5Gv9mS71FhSsyyJ3KjUBUbjbiMagj6srr9GBDuF0jt9RcO
KIkaAckRkQSvMVBbWhMNRDYyVYfo8lHcA4NkkPZydwaRoglVWo/oEW4UZK9AxCVH
LqbL78rnrcv5upvh7078ea7onkee6w2xxlUFcvjBLnONZbMXHQRrYlOJ12z2lD5F
2bbCP3qhGz7TXyWeNpbto/hZ0mttIJU3XGOzajk7XTIlWPNz0vOcWKmsSXSoGo7L
NVNpbIO9BkHHjOYTpi5HS077F1mI6cnSmY792B2MZIbDXtCY45F1pR27ZpfO6lPd
3/oiVCI+RSF0ob4b9e6hle3Et+kWWVT+6+C80kAp5mo3uOGgpPfx+YzQI7xykhDc
ztFa7aL2mLZ/pLlquxD4bulVIPzksXsUQGtYgR8oLE/AXHz4iE+wSx7++4Ld6b0m
3oxnWbpccZm8sWbGcXhw7GOmj0d2+stygh4nrSx7lckaFdcxQeDg9IKL7VacZ4Vp
u6LT+6zyuELx3jjKNFuosHA8ySyZHz4dv2mDRUusoJEO8b2adJt15hvcGfNSpZIh
bSctNYK3yqoTG/3wz8Ezy0i30K8+JLnhL6umVKOp0WzXmj5gC3E0KkG+aEn1IsPS
QfPXTmNX/Flalc3Jo4k48JZGj1qeTCc4z+XLCOY07O6J7+VcH8eGS+IFVr+TQ02U
vvqd4wAeNPoc6oVWs5673wMNhntDvjHpKzqPwh4Dq8HaKXzJ30wyj5W3ctf5dTn/
L7b+gcfE26JKnoRDe2+qToPTuGdI2rTeYjMhvjDPQYt+yeGBlf5r9LE3biv4qje3
iwUIt1pkRR5sYKtj6NdpT36fP9m/w0YCbPvEdsabYZ1pKYp+oxNWdEW73o8ZdCNL
cLAY+oszvMb/j/qlAa0mOFUeLH1PFXQRNuR2cvI04x3/ZE80bHACU5bBhvw3iIg8
fsM2rnrIJ+teDGngva+IhMMoTLlfenlxMD6qqGrQpTgP2QBJ16J5QFOcqQxtCmSH
fQwXoDEYBsYeFXMVK0xaOv4USWRhsTu/qjcE5qvMla10ubOwPRpa7lfcUNSCj2qB
5bgOGEbAxaQnFGULiYh2BMTtzUQQldZ/Xi7JQzIn3Bc3u5MesBLNE5zay3hzo1Ut
Lg7x2R7dsaGuZztfNttGPo8pd0t7r9BI/uqdZo8vmCQ3NmbUNUr/+7AVuYLVJTnF
hdnCJY+yvm+eBWV0dNR7p7yARgU1avbOtPN3Eun2pHTmCezHvK6DgVix06OBMCu5
+IcJmjVz0rkjcvNSP+QRouoGBK/aNEqggoDbCxaaZe38R0FEui0W39wmO0yh2KOY
0sY4aFXWSCtAHoJIj4SbTbgEFkqLCLQkvBaWb844KmsCbIzc5CCFytzAY/4LJdL7
nzNrPgoXKsSgEqXTNa/VsDhV7r+YkCcTGGCkodLNkh53TCn9rAh+E3yeWQL/2mO7
J8F1UgRM+mO6LCiyvgmd8gw9642PH5m/TQ1HuEyUsJakIrI7h6o0oFcymFh11GRk
2VtNbNaHCIjfJwvRwusyrCppit6swKB2yKu0774aGK9MdJuPYQTEEfz6o84f2lYD
LiyWGwpVqV03NsXy+U5MB204TPa/iK4meTu3H2kIT292PhDYNCr9s5ut8VGXYxvE
pXZCOam84vghofJutyh5hsDlreqzEb0rxaoCFbdNlZFCbSD/7ZTYC7/JsjsP1/iy
3NWrlwlGHIsjR6u42j2PP2SV+KfXqhY5M1qrn1zlyS99NU9Lb/eoh3Ng6hFXj/Bi
Hu+ToDxFy8K5uRExXvtQ2Ha4Avr249Z4q5ETCZRlsgYfiVBh9LUeY5TNTowwWsyW
gUxjXS4RrUFopwEEI7ggNp9wVEMz9hukyE8Ah+JVduRmbx2eUSddDIyx+MSFvxlv
iqQz6a1NflYZpHEOZwOngWg2Bd/ROapgocKCiIk35JUUqo64cuoL+JTXAYSJqshH
p35LSwUf2uZYNHXgNqXOrLbWsCkNPS//6vhlKXOHtaqoIO4Xbm4J8xR8FkYEDqIw
L6mBfa+w1Gv9EFKu9M+tr+Iul4HDeCv2uoHAqVAqUzdNMNJ8+EvFvrv8QIEvS4kD
XR5F2LFOYVjNeKs982boz3JKFaQxRm/rm1bM/GXk008Go0pLmzsWeX4W0R38DQVP
AQZj38tIftkcuOFnSTZZJRina+vztY4JuhRMsTx9+mltQpxqaId8HgINI3j2uUiT
OIgG7flyy1v5fRsF+OWdovZatMiJxveqSiqc3K6hw2s4yUhXQHHLzEMxdKmP4nnm
SGVaI2knAC/oI+lCjmbpuwRsxx6nO3JOejgikIpZ5OuFduuAwe2c4uVw0kImSEbo
xJoaMacu/VqpjiRI1mjxScWJIH846OqZ9We93RNtzGEbAgQsk3j9Sy4sKvlTofdw
1wlHH4ax6bpRe/JxebEMMrDD09CjLgzHmGqc+ior5fkKaTx2D8GDRIQYN2digTui
HHib29VgUAWr2gMnwyQhgZCnkhbuPhF+ZLkJuI39VxGhkAqI+9GUQQ+JM7Lcocts
Um0fla0HKt0CUvFl8575ANP+kuVUQQIEsIZnrmowiSk/LqhV3P1qqMFI2qnZ8lAZ
8/3udxz0SAZzuFfLqi3NZQTk6nKh1G6TVmD7Flcg9A7YE1r1S5z0MHHMPjen0Qgx
Nh0ZcM9art6Qv4gPj41YCqpt5eqpaXfyYt3rQ5fCsLi8FzHnOXc1GhHw4Eq6ha3R
X8SOzv41hHwPGoLSvjnh3Jyw7IHlVWlLV+e3s2KivjzQBGGUVv3N6yaOnO4oyetm
0HR+Z5sUHrxaEZZSPWUS6faers4Cr/yIx/p05kpfQJezlNvt921WGaOnKoEDMEe9
T7L+FmQ0clP9VcfdNI8yseLZXOXK4AEcvWkfJcPFJXJmdsn8pdcdYnGyG3BPGFxp
Q2UC8/RR5oaYzhY6NRF1M5AaCwGJZyy55dPGNMiPlijPab2OQ/BLoqY1rX3acCn4
WLx1iWZLSTGr/VpiT+AGv+ZenhfdztNDOGQRxFcGsF5Ifzl8djqWLvgtZp8ihsWV
CjXLbpJc+Q8dthMSd1Te2hszlJVZ6ajw/XMKdtq7rN7TJDnv873jf3DzC9nC3iyc
/dCXxGlKEy/hTWSMV34SSTYrhZj02bE2tBShx0d+LZRu6V3WExdV12y6Aig+TQA5
HFIG9yytKM5vuCRO3M3VV6ddsHxKIaE9qIrYDFZfx93BOqy/3yrBlBgdOHqZE5vP
gGKawXQ8VmovR3rBamNuogT/lINEuteQGLp8ZBIoayPmGyegJowcyBgiXig+U8YZ
DN3TDheq0dq+MLjuXtGYu6fst/KEZ4ZxIyZbCTX9TM4T7CpdvVAB3V0GmG9DT9pX
RyqaexbNIKpwSVXqYY9rA5qska6OmdEY4wMYPgkq/HT7/q+0GAvWpwZvbHfVm8ty
Ia+CRONcU4KuJE1z84ju/8QHAF0eeTvLLJvXn2JPCiugci/91GuKr+sS0GE8btf3
Pmex3XIldkQa1I6LZ+byB5RLty1wQWKA5ovh42Ll94ykMUaw4KKFaLGN+PCHdDvN
G2Oc6SmgvvbcTucVhJsW0VVMdU31JWErdYZ0DwmahzvjdU3Jo7TYh4uDe/4PBGfE
aIyY21hvy53xITeRHedyBA/NvsVAmcb52Ehl0LmtFH2TE+UipOBUw5TYzrsfQwSp
KSiZ02kxwoUOKJuvk1TH0DaXp2QL6BrKtVCJCh7Qvxl7zEoVN2sABZK7g5g2Ee/I
xdRy5o1wWcY4Bv+CHvdejEeWxXOp39WDLnPtvf4WcgldSzVAdPm4WOwtcdbdR8y0
iHjIdDgcQphV7JKNACxYi44ozXurusLwg3gKJUboto5qWVUrkUxw8j7bPwpGaFvL
4RTFnuecO7us1d1f+KSaKRb0ZawLreZEmifRISfgRQy4wgc3M/kP4rlDnGJjGujL
jAGhTah4DOLS2SqSUxU01c2J5iXsWQXg/AOEHuRtn5WirR8n23U/IDHavzpw1gXq
ITE0BVrtoIt1zX8S0g+Zx2MK8ljuH21hJXJwSkrOxNucxMcEbubIbBSm+bojKB4D
N1yuTFzB18nLFcDp+TdE5onnw+nQJAYKIZqkJpZmB4+gn4xIMEji5o6nRRRHAbC0
aZVb/Ybb4orSeG+LJS2vm0mw0LjlTP/Ha/Ti1wFu2j5+R6w2ZXCNpYxjh/TfQJ1L
Mbde2Rw7DbRL66FaIhqFwD2e8dr8AOHBlFKozWSobS8loDKCrKMn0PGDoivbYxcQ
mfAcRUe39oyWKlTjKQsqFXn3RiqMj9Ay+/wn6r3GMitHqljK/Jtx1iKYApqOi/sf
HU9Byyt9pSm/O8z7qTpECTUV0OEqLcZHx1q6WoS17zuVL5/aJ6WG10ub1M8n7JAA
+qwtc1147+FfS3jMPX+AyvIHmtcFbE5Q8jSxPdARhvDg5r1XoB/MStAUgWy7sGKH
SzFBJDnvY3lQ09x7DvSYT152m5X88ff/iLmQKwAIxkoWKKmUAQQtop/+CCuxIWfF
2oSGy5kJMKK8VREb3io6ucX5Sn1EiF1YkmTgM6Yj3Oivi6XlX17RInFAM7clY1wL
hspAoC3eqZ95MvG1HwqtV2VSu/iBqyjqbpLbiG9rqRrWperN82urbWDsakCLbM4e
GtRS/CucGzchuCHxWt6DonZrAalGvRBCKlQtK24+8NUCJ8yzKrj+Ave60nQlhqtj
wHDZikys8Ep3YvwnA98128qt2wnpUQRkRX6Qo1ww1ASomZazmncCrqN9ikfLOh5I
w5YB/la4SX/g9jV6+SzoOxt+XWjhDf+BYEt4dHXMzfsg3zxfdAXosalGA1SrGmOx
WL5k7FCx0DcrjAFklrTwgE7DJ3ZF/HY+48IIHbtDaMcInxWVUln+NEzUljVawjr0
FJTGOZy9zTPqDxoGUg1CpgACtXwo8LQUsyNpVComfWChZq1J1MKQ2+T4SjK27pAf
FxWWBwOmfR4wlORt/8KUEiWI6ijmNxaiq5M8dkgFogfgMFavdVlEZvi9GpqkSH2n
Bbq6EhiM7w3/lsfuPg+6nOMN9zDwW2fNBE6N4/SnsZJ3lf/C884fgq3jNNnHAoV9
HhNyl92reqckGF2U6KK/JA9adz7W39jixudBcxFhCrmPdGOVRr6/om0fSR07wWD+
067KoENd1xJFOQ5bLDHzDR5+nmNN2F4Rk/F5P7+iMtF1QjSWdWSZPQw8K+rDiMeW
cpfOocjFxNpfoFNR1isS+8HoyNK5KM8ESVzG2rTwD+TyU+ML1eKUAuQFFKZKcJ3T
pSC88vlm/YaRPg64CS+SUz5//XOb8vI4OF/gnej2f1Aja+NyOUurLEbWIMrDhj6t
5gnpEcYYr5xateVq+C2nuv/3ygZC09ybN4j7O0jCYHeUs4EgpurtOzsragRKf1iO
9sr3IOwaCtoekqYi3mycBiG/WilVU4bN7A2lju8nKV0vUZrt3I32nHCTr+iYUk9c
fxiDnAJdzIdopHVcEYHvlJstmagVpmFoK7zwAnOvuD091s0HvlDG4/vRhS9CN6ME
+T6I7QdjReynoaMN6/UTvpyfb4dXvkfMp0dvAAtDUE6Iop+3Kh/GaaMk6xI/byZ/
ad+O8k6zCE774hLhs4pIqBid6AOgYZ+M5B1DcOfpiBrThEC/rpgbXcUeFjwp4+28
f1wLDy6D8f8PO9HNNcpsm/eBKLjvCvsU4A6G7bx7uxiG92IBqfYxdZtXLNiwtbwy
y7uT+pLtlvl5EOHXixWgfrRMCMZRHqXjEesgFItPonyBg2PxMLuN6Mnfg5P9tYq+
5qhYuRJDfYUYvSpbTN68KZ8JnZV1VIujHpvy7yuKl3EoWRx5RZAgtyfT5oN2H6Ya
EZP2v3ftu5rv8KaKs4jcrdpqCP/Sl435Q7GLCN6CHAv6P8oKQ8qyUBHkXWOSNikd
Lu0BsnyZNNTIXcMDBbNzLZAwOSQmPH7Xg6FnxscdBJI/STxEsIUbAuLDtW9G94a+
KoJhxmSXje232kl5i817LAoXuW2te8gtitzO5wThsuq65vCFIg+2lbO6LWrTAZUE
SeoUvSgoS6IcA4/ZTZnquyg5Z0M7uMSYYsZvO4RSjYK8mkSO090xjZNzAtKSbuMn
yIXfSkP0KbAf4JDArdnRdLtMr+iPvgR9vf+ddySsSSgrHQjBEtrngOWCb+Gbev8u
Iy+DeRHcS4xz6EEiD50s94V47+0ffs96RkRq1lCpAcgpmTzAm6wFkvpP2xGRIf9B
IYhTWboNF2gSEXQxsJ44wl2z9G6mSBoV9FN34PxIiKiOXEKvlFI5r2/G1ksWs4SF
0ZE2SCpjzFB9wYD5h4vUazMm5Hn6aFwZVF2r4bIUmHHBLDu6Q+DSPC2VNEo5NQhd
mjxx21q5zFAkgGqzvX/Bn1cBMlj1TD7h4X7y/aS8AMzKmxwZJDzhQ8ntt7t1pLqX
pu+9qM4rvNINukyO9qf/Gfflu1ePPYIlnjyMTPL8OPtAZyn7ULYcaRmtcpt39J+O
ctK6XpwxfhLQnqXsXiI1jijHZJsNppB15F8f/VBzH2az9MmegSKOVMB+Wd1GXLiw
/n2RdoduRec7Q5KflzMBpmQ20WFhvj/JpoYZyZxp8heTSXTu+/RJFwTtxHaZoAAM
xG7GYNwajKVbtGRlksSxLalrDVGsLCq439iV3k5inCl9njlkovptx8o2IYAuf91I
r7WvoD6jOLW4eRc43FXzMFK2V2Q1f6UYt5nBW2Vpud/VTJmEQwhLDmAEOopSVIlS
JHa4urhxacEWHwVKcDQDmaCDe6oiWmaLii8MXbnS6mCv/WQaALwMDFeePQQhzE+G
m2kNV+FKDLtAC2S+t9g29Bpdw02qP/Gh7IBJ0tk1tC7DYmO0p99OLFQVIo6alzU5
Kh3B3H6YnQwc/AWFg5MCxLnESfLgJF72Sdmqo/s09Mf31bI8OI7TL1yLq4FKwxjc
UHPktB3BK1sAZlfaUnfKEGcfLZ+XLwSfoacwpFaRCEyNZLJ1NhY7pX1GhtFVNlDA
l1II+reuavg7tutgNY7HoboDWzbPTe+pblGaWMwPDdVsRYugqQXodu15b3g9TRD2
zLT42tFEf0ZiZurUFeb9FDpmWhl0D5eXcBxwMEhAfi+G0LqOynohYDaGluErDPR+
0efFgPbtF3EmnnZRNpSKSbizCxNVwSuleef3ChUdo6mOCWQrkibwK2rT5ba0omeK
rfZnLNOvzJXIIH8r4/g6gP3tuOFnY6uplS4ROx19oBvcIIVEIfqDaEXpxOOt98eu
2XlZv1s91CFuA0XvWBvBqagJ2QPkQNjB+/YJT+ppFBSveb9D+NwKqmv/IViXBmAp
gWX4oBQqrv5fgcSlZu9FB3CeoiHOb8yMK3ojFDw0g/dz06EycDaK3SfBHQaKi1hg
ZBRC+ewXT+rpRVFlD/bxiqcuQy3NaNfLf68kyS7RXM7iY6vdB6g71G8EJHJoM43A
cgJtyXX7zXMr/XBA2j5b+PCdwErx37riluP8cHq16/9EJUXxUQ6h7PkSoSr1jQsH
bNI1uT+Jxk8d5UA5bq5UhEodc0LNk9/t+i/DsA9I2+8q9HQq9AxnPes4ETU1LkbN
MpK7zVWhryrccreJyE4l1mvqyZWWWXrulAy36faO2CAh+kpzLaeipuNoI4YIdI5S
0I9XFatjrX/hRhx3lffp9DEfMknB+b08gCxQWaRjdeF7SrebEgbVe9R72qlL72RO
AL75dx1R7p847qzSV3OeTr58lR1qQwdTT06btxYhqpBWQDXy4cIwhSm27TEBfxp2
kYwbzzbVBENr3MHvAI8l0Sz5OQQjcqyuo/S6QbxwHeDfq7k0EehFL03sDAvZjtEV
IbHMlYsgVld46mVMAYbJOq3SkWZPOdOM4ZtlaNTHTA2NHXIbAq8wf+eibg8ejaWq
lkikmxUmGMpOoglYlzvhHl3x2H62KIemAqEpT9dqkj305/HPefFpqUBzcK8tpchA
rgJHcva9/hSxDmp4HW2OTaePR6TS6SSdFs6NAZBiS4ZuNRGIe4dmWCVSNHf/cS3M
6uRvQ7LerMFvGbcT20gdsgUeACwNW236M2oHOSeYUsLc9mHivKchm/lcabiozktY
PlPiwdL83iVqX70DJNKZaNaD4Pyr5nGgYhh4Y2MxMDZv6mx7aOCSKv4L1EHktRuV
mSUsqFUmcfSg3ys+9TCdXOTADW+Q8onWyudUtL1NEgi+BWwBPQ8lPGqvS+Px1372
IAK80qTKAjJM/n6qKMw6Le/M+Hpshe6bOu+qtgAgiQtoMW0gSMA/33fn51VcNxdU
+oy1xX7Us6kuNbJfwPYOiQJTV1zkOTSUJdQ1h1rFW6kaJ9afTSduKGBh5rbRdpyd
4fsrdVeAcgV0JGjxngN9T4jHV5z2uIXn8YVW30YcVbYJBWQmR7X+MO766uUXnM5N
fRyiBC4hTCe1iyAEGNaC/XZIb+kXkQlPVNjWfzGHKsaiG4+Dkb8P6rlKYfRnq70o
QQxrX46nq+vEBSs7TdnB60QqxMQcnliTzLdlSGutk/IdeOAsZnFXmPZEPjWMxE5b
PhWCRbnYvlgJx8yopPbBU6VINvZYy31qnw/LfuLL7B4p1ztB0ltUWipRfDwekN5W
K5N7lkzNZe/s/4a4Lk3Y/YAfHrSe9njXPVeHjgxaDiKbCea63SrInqUlbWAidQtm
PV8U91VcL4kQlVSFSCDTvCJqOEJ3IrR5hiofCxnS2zEGwVYNjSE+HFoDO/yd/T9X
Akz205U2dniOocxVPiZbnvevMKjz6xv5lPLmNGCZO8i87aLO0isvlH0rZB86wNPg
C7q8bXLqEaMYwlAetR1HgIg2rioI/k7RhB98Jq10AhHg3rga/BmoEqGVRvDzj2G3
x+qvz6IhVyNNYhIprAB5BSw7JKYgvqpzjPtl//iDj8kijWXcWyQXwgPWgR8a/dJf
UJiNF/7EqkGlZIj3bCbAMoTDsi4laCJM7TQblyJJnrmioZ51kgUHp/HzUXhagef+
6KqGquBqI2Bfk8L+zek3kgpNQ+dSQZDwLQeinosm3NX/Kolhv/Supq0VKNGioprP
/afzPoc0r6kAwwRuGRLJEcIcbbrxNOrLv4T7vbeFwj5rGGJEdoMdJUsmSVm0Cnca
FDEx4FaLXdEptBEiI+cvwXUM4I8kdMZcFHSx6QxBM1BJkIvdgsnNuqOSiSO0+jL7
dlVb4itkyR5VmMHrKuKM4tgcsfNl8AzK3/tPdwGj9rF6gjUc9alTh6F1VCfUjE9j
C0QhSGviWxjdRFPRc1jGI3p4ms5K5YI0IBcCdbkJSzYtCZB6QL8Jyl0xJe1NkO1u
ReCOy2s7s6wNey9uNokKhnUPYM+cdfHBVoQwA++BQwYIaMQ6ND/o172UtM6BXGxK
TcYQiRhy+uAR9o1bXzu7AX4xl0ZnDIpRbGkt4wv11PiQ2kLeOEZsb7VVzczwAENs
O7BJEfc2m+s5xRMJ/+njwAZ6TwlPAhEzgU3WTpiat0GwLiorZTwZ69ImYqHlSvvs
F2L4zarHCC9awmuygD6Vh1mtqo5iWiE6nMdcOZJA62hbXQwVkN+Pz9BU3890ldk/
CrgbM419hilf5rQofCFLh+ZT+MRPqeWYQhb2/noMfhGyFXppltxueyAwfrAaqUBx
CyPGz+szjmEW9IXF680XniqEq2nbuOUITDfkUDZDMBw9DGjcawQyYiMj/3fS8n4z
hCHwSLIg13jhnsHOWQlnXENK2GISCaeGkx49mfkDHOi/sy4r4J2elEN4ynnhSMzw
xsLN0A4o6e0q0oEzUvBfzS23wjsSI6f27TP8SqIsyn0a1EMhopQ1TPg5cXmi2owm
7355ZEv/NcZuErlZfGz/FWxgJf7xLFCTNdJIBfM+oFs+IfsUi0q7bIkmHIrvdH2v
Ct3fK6Bj8EkasTnZ8dQ9FfWdHPefV4CBcqzLTun6kXQMl0oWqtaq14Onr7NAi6F1
urwBO78ND1un3mxcQoMWZeIS7XARvysi78JFyFbkCYzrxmtIWMER753GMXk+ETes
1BS0tSOtPMEwcrym1OIMr71rHjExQUWfvK1RmJpLc+82aK0V5lrwY6iHKK7tthaz
DKkvS64htTaIqHuAgbSs5YWJ29+aLheC3frdhT8Cxw71+7R/4W/LzBdABOgHVMjS
brqdYzM753P9VWAcT3a4fEvnCHnM0IoaFC+HayyIKQV5T7yeuxPamh+dmMWvDMst
JbXCN8QegTZ39F+ExBucQmUBeEVy9cvxQYhQ2P3bCdxJgh+h68bYiptktb5OTIez
9VKkFzsoruwCU9Cg8J+EA5MBn5+hHe6fLw/r92JbzBqNczsBSmYURw1QY28a1lkG
D+Fw8F92W/4euQJzd/+CYwtiWLG3QQ7wTHUObfvWV1t5mC5+h1xbtLAChkobAMfQ
yv6uG4hr3T3r6P6afdLfCCLsWThbvxHQ3Svm+/qg6wE0Is2qo94GSKh6ri+IOuL9
/lHNokaH9RSUKZO7+B2JK+DuR3qvoovRy59L7JJVioZN/W4N326qeXP8OYlqid/b
3lYoEFr41dvLvAaMKqtcYKp0Hevgoi+yYJGdAIQ2JJCmhss6bt0XmaIGGa0CI8J0
ou3iKw3iiTuNdkKl5PbG/y/0fn4FRTqoy8s8uEJDyyjSIy5nI08PjENHfJbqG1cN
EDwCxm4GHDDMAECn0gtQEUtW/6lcf/UhUz8vXHOEC7Oz/nUKAiNs4sNsopa+3XJp
Kl0IS0ARWEMmXJYLeaEHLQJXPCRVe93OnkViMjYiGDu34RKR1uZz1L0h4rlGRDkT
xV/M2Pxn+dip0R0AH1Y/O1YGXyN8JDSYZ7r4ndIkKGAzmkIGfld0kAPXeEyRUiOm
tlpWLxC/nE+21X0MV7wj9uordkRah0r/4vMHwTt4ZOkwESdQiczLUfqQcptsppZ7
EoVAgVmmY3AnKLbkKQ84ZHuVje0Tikx4nAmO0kKqjdgELSyUvxoKApSfHZ8qvTuS
Q+LfsC3qm2l6nznJBZ4/lL5zY15EWaeZBQ+mGInlqEkETcNFdYl+UbVZyThjTpkp
KOzOHuuQLfUyFb3PZOgUkljO+HDbf8kOm1ScisJ3Cqw8zeSsO/w3Cua9/z2eH0KS
A1FgpFAlimshTu+tWLETn9yZK5YwcELxCy270unQFS2uxr0Hrv782lMlPGGRGi9N
L3KUJuK4/4S3DhgYLcPUcn2Fjhop5L0omy5FW1I7mbMmqXwzeQuRpxrc8djchsfg
T6AE6goF3mndZywLmOIf+C6HYlOIh/CcltUMWyMe6X9cA5xXaCF16Ouohs3Bmwx7
2aTN9dPbH2Q6zAAOy90XzMYY3rt65WOK6UraCY0OA6ewA/+bwejNxmT7uQs+7S+T
hHZE9qq7YuCoLBCcFDeRqeXhYo9fAqZZAgzohIiDRa5c12SZ8Zmq6EIDtset4v+L
tnwU5rimg3z+56gh/XEtP1D9ufeAnTzB2u6wtF59lcZ3rCaBka7B9L57tV1XkKwQ
IXXfsVUhneoUdsWrTK7IckHyHuTYPvubP1alPqhhTwdNehlE12ud1Owpi6/jkGji
60D8WNdjBERwo4/pVXzBuuAwWL3BP8/BpKavm92ndoBX198XFdGehGNiTqyvq9GJ
FUV5Ps2xknD/k6Lmo6DozF8MtQqsoH64H1+Glp46h/Wwp4LxjBswsnfM+N83wq99
Zxe/qEh0ktKWBTEPks/eFl9h+tRyf6lYmgjBNsWrmqilwj5Wb2Luxj1RDB7ePPaf
XMZFa5oB2TZ+4/HaMVAtMIhxJaBpEqcLSORouegyoayUtG5wS/A4IUWLi7DTltQz
kAqK8hQG7zBdM8D2o3ophlfYMwHbmlBK78Xkt1LkgazZq6f1CkwH892+qnDsz+M4
AisQRGY5Ubthe/WRtSdXlzM81tYuOU3Vq4bZFP4PMOIoLh6Tva+mSYcyyVsUQ+Zy
Drs9ttbp2x/kBzgh8r6McoSGltEM1Rk8XfK89wGcUNMOGdEqjIVRobvf2f/O0Zgf
UM5mIQrXpD4tpHx8tSXBtn0xT8SJy2F3lql2EGJqPiptfkb1orwVXux1b2Xp8xhE
wpty1BSNMQwMrkAv5meQ2HQlwQy8NlSPdfg6Hi1QG0A6254EPx+1XLF4GkpBSzsk
1aDm+0SaW+8BPmJKl287JDZrRXLoUugQWckLtLZ+FmW5ql87etlOVe9Ms1xBCQ6N
ku21EMzLXMEc76J9clKBNhPNjqx84O9oxOP9/qfdUM+ZInnvxoCnQZlYdYktOxFm
LL/BQU40yVuOfVnjYshZcA6nkLoBGPPh6pp0+xazppPEZoYvU2WwZUxULXtUsR9O
6k//QEEQIR8QlcWhHs/zMLRHTDnckrW9hgCbkfd2nBjd4K00x7U4zFurUxMOqpD3
O3R4HGijEcT3md6gtjyWcxdvs7uM88WgPGcfCILKV9HLVgcTYPndHDmAF2o8aIsk
jdDzKNqgWauzD4RG0Qt7wFSjjfkwBGdv2zcynDpClv2cVlpoOKz4ozcNZnIPs0y5
sCyTzmLbChOmmhCC0RqPBthm3kREeflytWV5BhS/MgdPZjUYkYlP8ZLmaiu00f3O
o6TyUgm+4i++fy2ql6oUijQZUJXpQNwfhFYUIzmsz9aKZ7mFdI0+1NEHXVZSjy9W
nWVINo7asfZmU6Q8b8NXjxH8j+FQberexKe3epI0rrJSzjI2e5vevx0ES/e9MnXS
ifDgpEcfCaEewf80ab64b15t6GsqTzU+BR1iYxAkgkbezJeFQYPDDajb9/QTp9qK
zKhSxw/uYtqV1pMiASkQNfnsP9vahUfnuYc6JRFOvUcHZ7dM6osROH6bqIQ+D0E0
uZ/mw1Zt/Loq1xCZ3ebSb36NbkZtLNRFFQJECoorrb2WzoHk8U5A52Ih8VazJ6DG
Ka6Ae3rP5+u49bh+dMOZJjpJAEfJ8+NRw1hsh1aLlc5mG/EEw0MRPPz8bb249W+w
Bwieq46yVomn4APd8AJwCbrIMZBxKZC3ke/f8sEjxIzxhEZ/fA8kxJiPlij/rYnj
zXjQzlKnarQee76oJYzMXina+u9LVu5r3YE3//QZoL28cMGwjcE+MEo1osaMBKIy
wz6r16YvRMl+k5ZU4fwjcuxT2rRZ6iE1NBV5zJMXAWSlY11A96B/5TPm6xc6AVDY
D0mE/zhDBpO6XvVApUxfe0I5FvF5B+2mgq4Ck0QJCCixkj1i03w8H4AcgxZTcdzO
WG/ZSXPi1htgFgQ2DeG26gNJe0sm0C10I7q+wz+G4iEQWNs2Adu772rnG3kq5E67
+LSFPoOg1xR1IXYvcH40qBy0/U5B4kexavtio3H4ck0SI/wj28uP3xtWIpsjMaMn
qrNp4QGZtkexuzYBFuXQ4wdDW3AZ5A2JVUStNfftvtzZymMFgZvnq7GQqk8x+G7D
Y8TOwHRSMrTXJiFAut0ZuZKvUHEXDxFegBKQYkrW5O4MS9GONjIXtSHjSNXuY/nz
dBs7tF1fHMyCP8ZK1NSIea3wSeJSVy/GRMhoFCGBJVRB77guSRuHK2yHMJdYDf8p
KkpfJuE9f6Os5U0HI7an5LN9Gc8M79WUU/NN+ZSOLhRjS2rKEG7joJCguz86Ivhw
gM4OdHryq4sunlf811uma3LhI5zQ/pM/4sBs71MVabD2xEVvtlWXndXxelMKB29R
7BLxAXVAgmtixkNBCVaExVMTUTKoojaZ7liSLkoZkSUEndl7JNbdlBDa60NkAKnp
ntm6+Jtsa7fJulHRcjoGNAKBh1wPmygcDBZHIIA2ZeHzVhJlRy04fTYr/ZyJWnVU
wlFUe3aau++5q6aYZD8pfIrw3z+pYzitgSrMp2WLNPM98ROnM2kvatSyYDOkyWo2
O2F5v0fgPaLO7rHmp1vaWgJ6QChNk9o23GuXPyNlcEDyqLzfjlv0oN4pglousXPp
SZ5zxiBSaQeuia4QJ0ceLQum3MklTy5d5/TB46yW/bRW4gLtYYSadCi3qSZQ6WVz
Qv7vDw6DD+6ErsX1M/t6K/tETITHuRSi8W/Cw2lMjS5Td3PhEGpMNk0ERd+wLy/0
4917hvMg1PxvYBQVYnIuX1cIAnqTh5BZeuBAePwcpxGQk6gSA0vEWu1/L1lBF5N/
9cJddwI4SOx1nOXevEFvPWV4coalopYr9/f2bbi4yuWOJq5lYYs1vKC8BxWt0yKL
HZGXxdagi6UsPZ0GCZ9Unma9xUWjCRdmDQZEXwdH3QqvfOMu+SJkhlH3HP6/gqmB
NR2q5V24bXE7FsTyuekpsoqJizwc9dLwmogMXlqFAjfy1/xOlYvnJXUwYyDU5OvJ
GmgPkzDUKfGgMoAyU2XOaWMbEbt9j8m5sYJqbPpALUF6RsMIxtgJRcVy2m8nQni6
QEEZx7iup7E1Li41/xsMO7KUwBLa8ZWIHFYJxLv0ulz33dvuaXbIW+WuGOwbIBSE
bdaFB+6qDckUhMrhuG6k5et2dxUiZUsyC+QAEFQJsKHReENOZfF9ClKZLPpM+BWO
rdx4UQsE6WCgxqbyCmTvAMFfsgDAF6iGJwehxNFRs9Wjg6QPm60GsXQ832yO57s+
NXXNOAqt0TWfg2tct9vLyuu2ae0LfLyG62qigw2BroHqf6rqWbYcRo8iAngCUFA1
4T3hdqLJwnYYjrhmVuttfGIcbIT6z0z1Kna/Hqe8oiELtytHA0B2leSK4uxeAtBy
0CPhWC+HcoSCdJwHCyqT18SMru2yYnc6pnPU8waaCpeBTIY0CDW9Fh9DULbheTmC
RMoKsncW/SlP7Z3pFqQNMX+jQf2o1srp2v4EMsj3SQFm5otQqvw18MjvMGrlrqq1
4+ATpzRlBb4qnXvm2/3lRM7wsKIuhKhxkPR/UaXBerBQb7S6k8+G+usgGDBYDdqP
140EO0XkDASbZemxIHXLZojyE4dZ9e8U5qmDpRfy06tDNBg7E4/vJ1c3057ukKG7
rmGzTKkphMp40ICP5t9gYD+h296oc/VUOyGCynexgVOz4ZgjjqwHPVnGj2g8SUKc
F1ZsqSm3YHIWk4UHq45OlnEs8zZmhooxQ1qtmuO1al8R/xSdQ8gACLUizwYU+pjx
8L+ogEVGRbV1ZPhKrz8JsgAdFlc0ERssfXr1C85P2m+vgFPhe87WPsisYhHXbkbg
el0/5PkVmJeC8ugcX2MdhQ+JFl5A59Tue+J4RIsr3g47jzZzmHzU2qPBKd5bRx1S
JTzyyiUxUJ0F70GRUDqez8Xzfshn5Qx+U511cqd18c8UdTlDr1f7UZWiRpPWUuuZ
EfLbaQwMHdxqlzYLb5GVGfruBpdWbNKXD89iyQdnYHcEVv9PO2Fq2AmNNL9Qpxu9
QxW4zmA07TA0g4dxP68nuzwz+r0bCfwJxrHAmb9xFcukyWpcr+Tp3K2DhW6r0JBo
zZ8dHoLUrmoxIKtwm6tLz2HIRt+xweoSx7O3nJnEbGNE04sITs8DdEDkAvIpO4h9
19S+ge6REjzbxeVjcq3pOHpRqOtRJURDP2d1OBucLATCyBhByFexkZryg/APG+vm
jnQA0zAGopF3nGbcgZ/v2XEY96t8pN2YsDEBuIkvEVvssJx+zy5Av4qPojcWGeVO
NAAaXVRXVjvheG1q3MgJYkMfun+H5K07D60IBOsp7+CEV+s7IqUyVCPlHL8drLqj
SzTPJQm2vSuJdI0UTvqEV/qdy3jYhj/o438vZ1ph/00FvZRvyDfrEZC15jfepP/X
ZrBKNUJoGlm3Oghc7bxHm3Fi23tGeq/e2fVctW65T3KZnVzzyHYyZ8hz1eZpFnDg
vqV88LtXJ5IO+BJZIGEqPCHI4IfBTBORoNwY3M2aweoAty/FMOc4u5GYs1Lj4CLp
qUC+WLjb3nRIYqAD57IDVwDpLA4tMHg+odlRbE3Id4oMa83WgDpDUQ71EMMM4gAZ
oVj4LoTFvKAptxUS0UrkWczFkstqZhfpfV5YV9M0a1Z2xpMp/gBuaRhUE4aoXh3+
thnWkoEuYbKfjwBeMfI4UIg+6oR+xckJJeDc4KODMi3m1IIaJMJJubh6OzDO3lAh
0Rz6+vOflaVwqDIkhGqmQvsJZw9BaYhnQACasxEVR0Bo9mIXbsY714aNbHJDTMjH
AM2rkyug011zUotnjxETFHwZ6eZy8IXVEtnhwmMWYvzZJpZagDMlpe7cx29QagFy
aOJvyy/2dWN7bvI2OysWgSv+7PgTqw+bzx5bKcHyB/UrGb2bTAJZ38L0hyto58ss
Zr/mpKObpTnyp/7PTmj+xeOuZ9mNIO5MhGvdx4Ud7soTaia+slfwG339yKzsM+fH
QHPMv0Om/H4g8prgBDXMC2ORRFCtxp9adz6Zqya4J6NISqurfJ5fPI+eEHQ0vqQj
kdAAVYix37mp/64MBHYV+BhStlfvQTAQvNwi9fhPEUpH2kom4pGo2qVysE/f/phj
/r8zjJBCJdAhY/aeFELp9yELGgOf11RRMApFyTlANi4JI6ApnqmwdAXYamI6YW6X
FhLtJXTEQsEvCHmxQ6E8/OTIl2Ql/XDyB8b05E1L3VLtF0WaGLYlROQ3BQ8r+P6Q
f7xX9DeDC6hfg3WJi+0pmnz7VRseJYmHqN0abUUfo+wfotqI196i075gXPK1lzN/
YlYocTPXOBqCzGpRnffFDlgJZYGYDF8XQRRe4Xs2cZnh6sr6pWGk8OJHwYp+g9HW
qrl392XMw8JYcbl9N2iDlMmMyfVdxiPUAFva+vTqvKCWRB2xubn1R42EA8gQJvsJ
ht1NY37uJewjqydpLabnoqEtWa0WXK+9yP3OQsurnqTXSI+RrjMMnp8wRAPqfhMU
RxvMEzWQRFnjcY4pasbnKKyM9j0vYjniTsLSntUlxHworZITNxWfxqLcyD6UGzdI
YYDkJuE/Os+NQ2QWy+02F+AnGgvxLKokODTEORH/l3OUdukaM+WkwcjyAdDaxfSv
Mcb/M3lHcy+6JncdNFvJH6EHkYF4sJrgpLGm0MS6/olfGGI2DwNIFhn84slBrEXW
OxJjIe5ih5go2vXQH27Ll6o01od0Y/hUPMsY4EtoA1FGmY7lERbd/ykfwZZbNH5l
v+ql0XE/Qg5gJW4+ndzDJPZkd5HsEEo88BWAjUNFjF0rsWwFWipRN+P2TCv2XXLD
3wJUkjmVOB5+F6uuCmJctugI64vVQMSMPFnCO9bBy8Cyy/oF90RJrLnjB3LJ3nho
pHBp6jSOvjESIDh9I1S3WHc/ZdT+G1rLwvsnrKPTsCZCnHsZRuqiyhKuyOuaqCxt
3pa//JlFxPH2fxJ4MZh6+FA7UqxIX22l29kw+JTEliaGPHjGBEzSXLwJn6gHl6wz
tVdsy4Doxfa1clmMi1sF17U+JbDsUxI2Z0K4ZMkN10D2leU5xOQJi5109UxLmYQB
SiMGNGZ+pXzRtzuBooHCUcWJW1iS8UCq31sQ8oPL3rcGJffeftSye2SJ7ykLxkVN
ZP8QLiUPANddS9uiopf9uVFX0VFWQ557ss0eIS2XZNY+zMKH/+XCpZ02ELS77NvJ
2RAbrzgLc6uI35yB9Va4+EysNpC1zTdnU7JEqOcrwzjCfjAl0fiAqf3F6gPcmzzb
7af8bhxWxrzoh//LC8TRJ2P1MDvfEMT9P2ruQch8/qzHlOBZeY/jklAW6BmuLBi7
hXpC4O0/vz1dr8ixQX9tLIPhWP7QKtJuEjNUwTCWTD/CcBU7gFl2t9BXijbFh4b7
YA/pzKZdD1t/RwBsDIRJC7jUercX2ro65qcvpLN3jlXNtEh7S9XQWy29VEoKt3pD
Nm2ZmYcBHElanvPi6GIonpYGf7ntnZAjVHKMYjvFLuIT8MUTy7kkOl+59lHFcCFV
XWBglFAOtolyP/BwEKvRIyZksBjE/yRLnlsU8LzBarHErofZP7S8ZQjsEyRE2UO3
pIjGEpSbtUoOWn2Ao0RqwRBwRVyBNUE9d5SwlWBo16CQQAzbQLCF5WwyMYA/h31W
o7/qUxxaorexTnv/cTmTrnzw+XqtJBo+a2ZeKqwSwgR3po/rPM4+4BUSZ+uQnxzH
muSsdzxXv31Uvra56z65novKJxSeayNT0nznL4ls+cb8mz9c3ABk4FtKVEQIr+75
sSutN4cZmb048E7wdrs8yHNDqaIEysKGNTInDdte4J0uEFQ3jzEhwTl8OGEb1C0a
ZVTasWeGJELYqytm04LfoTh7IEd+7eTxcPVFLINuI/6RU3ab/t0W/MsbirawSKUU
+Y8trFeA1gzpWJulLuCIjeP2J+ladFG3Us49/8MzbyFkOjXul+2m0xsV81jxJfy2
p7orGphjNTaU5fl45ghhUkmGvJA+65D2bjr4tuNJZ+NGTFMlNNuieJPvHiNzAe+A
aUHVH0JuLgIavL2nMuVO0Xt84BZObDqrR451994DvgewnqjtHcJ4fO8RbHkHAfD8
KnhH424+o0gsrD+ErdOzAN3ORE/482nY7PrfjZ4roRB8kj5EaU7KuVmJN3t61jxS
XRipkxam/TtStuOot8DBuKXjluA10K7/edYxa7yeIQ27AyHOeUWOODISfiCDF/1N
UhL1sTmFSl8YaLz5lPrVibgbPAi/SxT4a7VsvrWr/KPtahP1bdubdNXiIbczHfvl
VLSPD/WWQC1W+woa/R94UC59PWG/JdzeLrt7Z46rtlKTnYg77IkPH3yIio6LoDvO
F146QVOGP4wXnjbinkxO+Lztomugw4gEVG8N+AyX4zNbT3An2mNU3mqmHzp/auSe
HOpi3AjKz8FRZEVcKcRAoD+/y9R9RY8HaCgwTQrVsvSelebcTUb3fNiSPD9qHJsi
6aOOoqzaoJO4GQCCyHAX80WjyD/FqORaPWB/0IBew7+X0U4tc+NBWPtLSh+6MFHX
IvJEzCbMq9QZBZURzOajzVzaAkPOxxip6P8pXVjk1OOuXqCvNncwZc9nR60x6W9Q
DyAgepwTMJURlwreDeggYb6i8BaiP+rUexql70+w1bpMW8kMX6eQ8fXmfuOQ44Ob
qFyYo63m72iHp+yexXfycRtBgQZKAZf1UY7h0NcHrLtmD3l2+GniyXA0/VCIGGnS
AuwaeFz/iU5b0/Eo5F1uCTAZqo6YBqvqC7icMqNpE2QCoIMVXFD6KzuYt3UZhrKU
XBvrdHLpqUPORrQ5S7pd6fuXuEiV6olX22HDE2cKB6rHZHGeoPNPs0+QHDzoqJqB
VidFUaZmjmEPx2aO+LglGvLS8ZBS9avHBQbDG5xRYbuG2HOdp8OO6qver1W2fyBZ
5aQzfaykRv+W/8kENRi/g+Dlskr6hu96+qEXkbtuhbS+K1BBOHYsXlIcal++iA/J
kS2aJijHPgJH0wyclAWJzmdtRiy5C24wAtQZSutkZnKGSWBX2xqgi8AJ6G/L9e25
ilwrV5Pe+hWOjBDJvvVwdOpifBOHRRzj6q/s2Uorhtz6uL8f2nsUv+VBZ+PFutxL
ACkcS/hZkI11srl7lLUQW8yxReLf5S7kmDk3J53OKrxS5FZI7F1QzEGJYm5GaKgt
kNs5jsBUT2L+hTxWbHy3WFJr5YnW+q5D/DIBKcuuPlEDIAWNNqv14brvDJug6N/n
3EoJADiWc7a9K7eUGJzXQTuASwJ0uxrfACjVSOirTgYHzd4iidT5Mc9vbqYbWZLa
8TQGZl8pJvz6xCT/TprhbgZey2r7Bl2DhyjUgyqW4ZhirEUnZ1IKu59Alljy3fi5
oiLcg9kB3A38obS8zfbSU9DIoX4YGS0mKaYePQ5cu9j55S9HLh85M57GS4xM+8Uz
XtlyZSbDGWx9rG1Jc3uSJS80IUxOAS44Fj9EGcLEXJoGg4Gv8VXkuawJo4xftz6n
oEqgmIYChPnemy9kpX5pcxHEEzX/m1dR38szJqhQV9/kYYIbX50mxsZetNLRdLK1
UthyHoolWzfSMCl42Z6cWZ7c5JObjOs0EhXIDpFvaMc2LoeQGxOHV/uao17LVVHI
YNFPA1qJKW6EXzPg1F8eRXDsSjEXNlAN8vK/fqZLHdznoHM+CMZwQoXFoWbA4TnR
hHSuPFQPrE0cRzjtauBs5EVAznIXJv0sqzJqtX3G3ILGcTLh6CU+uqgI6mayhV3X
QB5VVlgBRJ4P/UscwZ+z91u3XvddUoQWfcm+ule7aIIBKW1r71p0jmX5ePDAkIC8
sR/4QRKJFPreUrkznwXCkaTUci2g07nIIs3l4n7QY4zoRxNFg22HtgMtKmj4k96+
6vOlhH+Y840CJVyaHDDft8xJb9GzYmmwiOYwEP4aEvWIaQwCGlkDM4AZaJVAVhSd
4nkIC2iwIe7q6X5pUDSko1Yn1AIWL4MqkWlGvKTXVPjHMxIlUos0hMEbw2T9nsTX
AUBVYIq13+fnlbuD5rhL0wr4RE1gU+1B6YaXpnNYjF9JNfY/14PNjy4hnDr/45iS
XJVVrgM8eJIjtkYRYQIWYwFIT/tu0jICTFJ8PhkZxgobyg4IVlHokxx3v0on5Ih/
w7ZegVGl9innUMX2MUez9qqcgekky4T1+ddBkkn5SLI/IBkLzsZq9OqewzuIYm9w
nLau5djC1apCrE3ptzff/YZruqdD4euyJoHo3/MeeJPzOor3SD0qFpXFn3E430aA
vSNJVJmLvefdbhak5XhfA75M4iBMxqa5H5pzu5yZjKHc12CsAJQLCSm6Xq0MStt6
z8XFUbFxK8VUDJXxlTM3dUyYsWT58Rn2MPgJsSMLkIgAUJYnK3BLF4QTdi/UjLop
q13exC5tioBYRz1mL9Q8R4H9r1YQtFvOIBaH+tmS98iShIiJ9fx8sdEDTax6Uxz1
3GDZOW9o05jDLlA3lFWvDmAkFd60MY3+VaNFwVTrg6tgrV4myZfKlS8zAXeBKKuE
ngMHSOt2t1mOLOIFU2Aq/Okc4zOnVBU0eLMOJCSRfNkSTpNBVFFRxuo7rm3UO68c
jXpZZpgjySMOtXaj6F/l4dTtp6yYtJPNDV3UjOQ/QVG2DMnyZ1JShqMMN5QaBsPG
MZ8B5ZudtSDjqBlPwbiK0FKm1IiJurTNqwp+qg4jsm7sR/aM9XnF1SlhnsUXLViJ
0kPXFMgBQsTvVM/liqlJ1dk4wsQzfs3Jux38bNVMnNWAzFPf1Z7jFIx7LhUWOsMK
tIC4j3U0rF2D7ToyDGns3oKFX+809HM0EKbpkHe/izexfEi33vOWPLbtqWXc0adx
L5muD2UCV/IajbBSr6Q8UUjsdLgQjKpraNFGh+Sy9RxOqrYi/LxQhOhbweCx6Rof
EQzgMz5OOuENHwCdd2W98tqh+U8qYaVFvoM7MsNi5xCKP6Rh0S9xf0YnIZKkxlk3
oaTIy0V4WdTEJtav2uJacC6F+OfXbtlJjYKE3mY7PGTfyHf9PO1EZTvCEZfIPsy/
xh/7RjU5QT13vZzjRMJ2M6VBFPI8OIJK/5+YfxXvJtoh/yo0E9orTgsSYI/ZoQ09
s+tei+MMesJhB8XMG3LMtWOb/pmS7hUMjty8Z31E0j3zoreNUMJmd4ZvdbpONNB6
hzRMS0WU5xrwxdtAOQf08+6hu4NQv6AKIwuYW1FOzmRb9MoL65Ryt9jDrehK1xco
EVqzdt7ced8izvyzFbAdY4bp64zFpQ+kfNqy5ORSxoXDm5R9nBCuA+nBXhyNNXi8
Y1eXUx/5QQMNKV7IvK7ugiLseQoZnHmCR7UenqX1fQHMPK88PvV9yYygbggYDwTN
nDncpxARldRXZk4K2CWSpn4uq/r5b/sobp6Lc3o+0wXzwu5xSK5EmySNXinDOehq
4KlUfBSjdknSEwCCT1meynhxMpoXTfHkW594WR56HmwTO/Gy82kA8G2egB+Mx1Wh
ifDDzQ7+vGYAbPoha2g4RyIkkqPNQlQ7r3ziomuXByynhYadW45I/Omzm2AixagQ
nx7nRdsIaTtaegdRWomne7mejaNsLRfzGHTm7DHi/dPKel/Cok/dktMvTMVj9vcO
pxNl9ykGOUH19mV2RalwfDQOwXdJtcvNELiHBY99Sv1lwEYTOQjWWFxUDCXqTB/e
iQndqtICV1kFsF18hRY0mUqjkVAFjarRnYNbvKH4/gca2uqMOHNh2hZlimE4aINH
iU+7KGRiH3e13vtYjmmte97+MYg9j0Hpq3h5XcYnnqbjQz5UUrd8WgirbL6xha7o
YSLQawxAFNMsdk3YdBbGm2RD8NzKiR84c+DA1x64oVjnANgSwYzOgC5rsu0F/WoS
j00AGBQmpmwxVdTAkXh+ojYpi8GkjOsxPOXP7jfzc/VCvTrZr0b7d2f0H17f5JaT
aEjQnVuKunMhogw5B3c2HPklzCZdkG1ySpQPW5viDo7fAFn6p5p9XR/HhWATWr8a
lNV5X38eea0xGw4ACodRP1b4uTQfwi9vipxq5nn3WoDGWxAS5OMLJM9EqYgVZ5Ar
T+TDegh02e2qqsDgWFMGyRaQ90K7+zARUlzr06jy0jaMTGNnXrgnM5EYDE+zvWYq
mqrCcuF09/UCmq20nozdKiHOAwJS/jhSJotIw9WIW52N7TT18vf/Pg2efl4g9Yvu
L2vezTD7aVmYFpzi99F3asFQyajB53aaKMWND5VLrNnMwbLlFwZhtZL9L8Mat6gt
mWt/Nf21+Ccus1/3rOyHhvFHe5lhsq+fSRcjaLVP5m1xGHqzasC2W2hutI9HHJIm
lwcnru0FL8oK7AROl4dXmzavujEdxiwxs9dGyOhoG6sGxzMFc4TcVV94rMg1R1ff
pLBHAoTj5HOt08AncaG4DXQ1YDbRSYJoUa8QKPRQ4m/wGGC0u3gah1jg+9yNFCzN
6kwRi2kY1X9A0LXniozQ4q48kLv3Nl135Cnk8if24tJYnzE9loRATBrPlYbeEToY
qNY63dZLgRoWbx7C+2y1GSf00MdbLMhwoxEBcztwnIHf3QkprXENL0kkFyUOGLX2
u9Ppc8J2xqPzjuHgiz1NhHygxLzBn+jRiiIfsu86nmF/cPHxbxaSpvTt2SG5I9bo
zig3W+ynJWpFmKij42N4UH/CZnraJbupaU2H9HTQ+JtekHQDu+FyADgQPOu+TClA
SZAvj7YRn4tcSe2TaqFNxFZ8jc3HzKdxo4AGJw1v3vqlGlxuq+zOwr1u73pP7UMK
Eu3dzzPizdmsMzW1ye+u26PnGwTjwJZesdP4XeFjScSRMsa2TQ68B2HnD/3b9lzL
O6k87stZnmZLkoyND21aI3Q9rOrgFr8QPQrr/n5km8vBvN0nVLlo3JubPjPiAqJ1
2j4yeLhTuqfYCFcC3u7TLTIsSGLgSc4xa9SapKL6xlz4brxWTLGuWH2Dd28uIddq
L2qZoH2lor38N6/8EsgY3WGnBO+9YT5mZiiaVzIAONkAfObO9phV6IktYupmCXRK
cgblxtVsUN7B/8EXwK1/HhgM5gcL1lxrmKweufVvV/GKUhzPmXzqq5uEwWolVej2
34QJYN45avr7t/KkxuwBpZXwxkVDsjRVESWwCp+ioP488SyDn2JMrhIZo/Hc04f+
wRR6zO6cZFvL1lpqLI9+mVZI8lLLufUKAv6ClFmyPALfPz6RSyXra6NQU9n6ARpD
iP9nx4LnPSB684+oS+3C1wf116hIGKXOHu8k8fVm1rbcWArwAnu7vuoQZp78MRaX
yFZHUq+R2/XD6OW1UFbrydT1fsHPItdWqX7RZZGANQRaO39gpaqWprLpYzEssw4j
5lv6B4fuXBfIBNHpJ2PxY8y3Vkb1QJrU22F0NxhZF+Q+RHwEYj08NmhyUkqWK6gc
L7Gb880naHAh1Frj14dAya4c9LpoJ9Cr81kChPkUa8ERP4m8PjvE8a6pfBe8E+uu
7d6oWx2gqwIxJeaEY4IGszldfKLeGrRshqjMsiK8lzcOvUuPD02qwH52KwnTE9Pw
pgMUdVlATS1UtTp5TC2NrWH5LcsaDgqAuny27nLWAvTNW7qhvh/J4EzZypj6LlDo
nhRVJ34iGlHOWmRAvtveVKxSPBhcQQLul+Xb5S/ZTst/777OlyipXUW+I01ewcrr
IocXt/qZFJcfNFxqg3849dHj6OJ5R33ReDwALhjWblM7CEGglfRSDytpcf8hbSpZ
LAIyUEdt+M1YSNkSQI6+Qp5F3ZfhB8VdSdj0xRWjH+SP/D6YBUe/CodO2nL2zD1P
vaZEqmScphYbNIyALKcY5LB1mh3wYHxxF/PUM2lTG5M+kxuTwx3gbMKrJ7uRgKC0
keXayMThNFkPnyr+lBm83DJzqBGJx21MAtMKeMI4QQMH3lWwAXB3nieBNngO3Y/n
YumtgVyt5nUSTbZQaA6lL6pxWp08OGmJHfpazf9ouX7PbiivIhUdT+zhyf3gGA9G
JMOzLINPoYtpnaGrx6xTSHWzDjikbPNFTBSPZ+bn9DZ8uyE/jZ9vRm1g8OqRdGK1
H5vOGHHyDOuGs0nf+i0zTOY6R/QzUCm/bx23a+Q0cCkzX/SnhDPc2D7IB9cxk6jV
IGz0DPnQk8J2FOZsNa718D8QzizQbur+hLMYpzEueGW+0NLeqC6U4zsU8jsnPL/k
CtUmyFcs37CmB9f1EkV+lB0Tdx3ZepFHivhgH1MroCjCB1j5wd37XmUhK+L8mw5o
KmgYh1litLaq465BTSqdBnrqBVuvp0JgHraEL7Q9CwGCegrsq+Sphuy9BpCwbele
tID1XgrZwIgJJmGgHWgFD4GWIo/UayIMhutfv/qc4wdYHB8Hb6qZzqnXw4d3C8MZ
dAF7g8E+dqzilRZmqMbt0zE8AqmKrzmtZHvIDzIvGe1Q0xNgDBQfvY9TuY4CHWhG
EiSVLui64V1cKHvol3hUd8JL3YI+tBRtOEuEb6cI9a/3JP2KR2LXyWPBa6AR6XfQ
JIKzC4T+hENEJFTPCOrX+0/xnglIYrPeBPF/AAHPzlI9gK35W4J14QzY1ygpfWHj
jht2KX+WETKxY3QLG7bykBobTNoGjwJsiKlbz/O6n0m8oIZvzJRI/PNH7GOqfJz6
JxN2h5lEq1t+ukTTarguThQivYk1FrFjbXgnjlFxqSQjRaDg6vgZU7DbVzafN7d+
3hwJX3gLnXEHZnuO5HTHLTPsCYEl6q3bMhtSRtUjoyfRdrNmsiQzgFJIqJ4TxCHe
1i0Jat6MQacN2m/hItSEW4KjsJl2GKp5umpV8AaTFrk7vAHDoDlUa7FtYwl+Ip8t
VER87SvzQieC9Q9n9B2PlPBqYF538XwgzhiX5NW5xj4UMXDqFlLyElNd9O9zVOKs
d7kWlWXQvFTkSXQDnACfN7ex9D+xDDq4YpGlf6wgnM3pPlTFitZmdCM42xFpwb/8
2m4MRtCas/H68ZmHjP/EZ/HRQLOBEKAQ+34xjIsH0+M6/D17mzuXc4osRzbfM61u
4a0rB0O2kClo98u/2ge3VPrr6RaGMigouf/lgOpAxn9U7Nyo7g3tqbwobN81j1tN
/Kf2AcVEe+JaQ8M4YSBpZVzSQX6Z7DM13xQp+berYGjCuZR8jyMPrCyVDkecfsGi
nmqYHBxpxlmEfQnzXGGozpcvI50iEo0zHfunUTyfsYwR1uxImmjhmGBvyLYQsoXG
r+yPj6jOecVGkoOhz/odpd+WVqKwouWrZSeeNflc0rSxsqeZA4Xl2Q44j9JN3VlQ
K4g7Yu/YM+JJIS8NoAyBw+iCzNh4tEGlVGzJi4SSede2y/fcXiB0a5mXGT3RwKo1
42wejh/EDg2hM2mCcbHW07k04D1c71pjAXMBnZ2FvL9fbdw0KiDjBp53Yxtzdsms
Zi889j8lckwR/CkDwdYZzIJQ9pUnKPYbCGpBsCscgEn50b1wTvEG1KCc3eU5xDaJ
QvJbp9Dfc46i1hl3++043u/fcj9HaQjqDfNWgrZyKygbiIl9DbpTH3UpYSueUv5W
TArfPM2qJGRarWlHOfRTjVJryuNTYz7jlQ30jXsb5cw+RZIP3ArQ3xtko4/pQfHe
Xe+rYuyYd2K72VxTSbX8JBETf/e1AwqfgqcA9uBDkrM1Q2nZEbJFNLX/jFypYN1J
b6XL9UgRl7Yk5rsgoMKzr+o9iQcaLA/JKQFLJXzTzwn1+DSKYrhESB4KCmiR2rmo
MX76ZbA+oNIrzr2Jm24pCWAbTg4IRb5432bXTmWQ0hCg0glw4Oz1mElMyRJRQNWC
lIsLo68xU8Au3TZFLybcHfbTnCEyD/aUZUGNfsFBYsTgCukkWhDHPGJcRmAPtkWz
pYRqysSBrH6FqQPlsSQTebQ8/76/of4Fh+523dZ2fzw+Ao7J5F6hyQDOX6LriFvW
4YXPqkJ7gjG2zFG1MXjRXyzlrX3roYysBOAVMIaMqKUWK+gfwkYC2+EbPnzBJ6ES
eom6fT10SKgpq4cx8jbDkeqgACuxgO5oKIp+X8GsqkbUcYuvEJhx2QE5+TYYoKze
CqXrtqR3eYeg4a38XClZQLOqw7BOV1bTsnDwkPbfRmPsqjapzBFmzFtF57wxViSS
HssuOL2GI4EjYIvVFWGj60nO0f3jzSnRXLYRhARha3Rog7Hqk2Xi9uL3HIGsjUjD
kEACck5F8rE6+E71Cabw09kqA9IH0LNrqs2HEj9KdRm8213Gb6RvAOClqWqjtDxb
KYHnPhAOUjsKjcnKqiiCZFbYVEWxdJvSBC/sNNOPdd6vi30XOH4h7koNhppAfTK7
v926UJ1YnXFRv8XiLTRs+dvzgY1imIO74sgeL7fH5ov70xiJdFEpTvPP36HcHD4Q
CgNVgu7gpBT5Hybqcmpt15ibQkSJNeTYmyFTolB1z9C2pCjkz4WBziplzn3gejBx
7Drj+xLW5Pbq1Oq/qVaYgc+fofT1Y3CRjV6W9cJu5cSNcR1rGZuCWQAUOjVhwP9Z
Z+c1qDQz7wUYBl/Qkw7Cn4NXllfB+JVDDSMfo1PPY00ki6u3vKQ2XxyYLzTyNy/M
DEnAUu/FGMAWsBrSGdn00sh43939Lkx3hSHoz55yCbabKR2pwnxx/Q7yzLPgpPLb
Dk42uQnPPYeIhKKRas9DE2ZD/T8jYnYfhoWEi3Wc0hVwUlMHJSoEr2NrCug5HmSv
Fo4beVCyY8krO/DyrOW+YyWVkRZpeTLW330nzvwGrBeL8VtucFAcsBwbbpCvMlbE
j9cg80Vz6+9Xiue7YcnNQb7E7kuAQWfxgEb/G6k6nY6c5zySgecr2Kmsu/DcIeNp
PPnVIpLFuqV26BglZwtV6vGlIoqhl5skacQo4yuTUmpcoSkfYyc84FKdbOe7floN
Z1yy/QaWzrhTmVThSFOFv6hNeOmpDuqeCionv/smOiKA29YNI5dX+L3I30TCCJWQ
YHL4Xbb86+EjeSZqRovvTzdqtPgWUucTxoR4HOxffw+6ln+d0R+FuAMigoyZ2xkZ
YoHn4NHiqbJc5i5RK8RBieUnZVLPHLe4Pbcj64Mofy0UI1NX5jY3Vwp0d0wezG7/
H5AIVZEseVpPIvEkzyZHRPeHbseX9CgyHpM3h89DCYBSr4N11n0bO+LLRwBw90Wg
2WUf/9F9sjmgvULsUFfktU3jNT7t8LDqa0oYkuNa//VEp2RHnEX++RU2VL1eU7dz
RwDF2A5XsceQC8d2vtuHZtb3AngkP2IccdRMGaLebfsoOcNpe0flUtT60jEaQw6K
N2QmVQuS0hX/BffY6XSxiftataEePErcY5426bXbNvGz/Dau8zeWmUOaeLPebtSS
JzUZEFfT/3uwDddKyZ6KZhj4k+75hI/iqdg639L+f5X9KjNzv3am4iWOa8uc3uUo
Pr7wEf4wUnCi0uffiFZUY49Jmi7Cod/eO/FvwIFJCDnVfP0UKck1/L5H95r663no
JRR0m4ArzssFir/njW97G9HTxBbuq1WzCimL2PE0dwCymLFTsHpmHPzbM5KdoczV
zV9DebmdBP/Fi+8K8j5Rw4pDj6M9UV7ERbjJUbEYQeyMudbHme6zWqOEcwgqk/uu
q0xnAai7ov/iDJLje35Se2pUjr5SrWfJ4MFE4Cz7pWGY7azPHu3c6/c4p2ZrBCWO
mYpacvI/NsdKD2zgpswkTYkHSXXBYcgfMixjrPXwppvIsHb+HuSHlNAvDEAH1ftY
aes9he8F04Wwdenqs8bqKelmlTQ69w4W52c327pQhKDfRUOs2RifJSROC3Mz7aKe
X7hCCJDp/2xHAx2wMA3QzXg39bzijHwa6srlprKwx4IMkTZ3xx6Xug9dsxGOW5Cy
R3niP0obUXxD07hXVIYSmoGuEGbH6cyCOpBDZ13pWwzzTN+rOGtgyTbJ5898Nl4O
QyW3ChEvoUcokw9KKDecdBqSPjxW8BTiuqPRTwd+o7utMG9QxrEo6YKOnaQZ1hbX
yMMR643XSvhd6JWvTVenHVwFMIrSuCtsuLdMsIwjdRv7+8k2k+VH+xOeRi0gL9e0
RZf1pJrHXlJ22dlwpBGfkWZe2n0PNpYVOHh3CR74XFME/1LZD1+gPiO1fkt9oTaf
c9v9ovXZhc+NbTdxoxK8Td5kIuxQg3CMgwTrcYS52+VDHJsgT/CV5MP0GWRohZN6
XOwAkIM6GbKkXyJFmp2O4I5vQywAeZTEi1XcDiz3po3B/ZwrwrApYZfilPp7669d
Oy//pUos1xwl3GUdYVKEQwoHei0wDt6uDQ3mBkRvXGZZnqp6t32HRx0BbTex/1rH
BG3zty4aA3uud6bYe/wFyI15bQoS2bRg/X9kFJYoFrq/NEkiQimvMwFFCjICjzF3
nuZccm3+EeZgmQfI7L58s2Amfbsb4qRRfm0YNJlGrG25m3wuiVzkGPVAhxjZFJVW
VJvFEjR0JnVgNg1/xzThVMBAIz/oBh9Uc+uZI4Cq7U3oAHueGuEchbjPOkqaFXDA
DxyYT/kN8pYj8ncdCAb+HhNPjj0Io/p8F4e7Bqkb2U6lMQHdm2D7dQzARQy1ou+1
3kSGKQwafESRzVXU+iwWnaH6LxFI1KNpuJb9i2qr4W/iMAwTG02lwowygVf/IB94
Ic9U9FOOBeWcjzXVYBm/GubALke0BZqqD7PzghaqThbD1HaA/8OhD8eN3iZ+Rsr5
vP9qEIX3xlZBOkFyLl8mJa+FfTQ3+Gt1bblQ2iq/sYsBlekETpqFYLMi5TOMBRmo
8CvBFyFV7ph6hWJhfhE5WO5lQl7IV85oc4wbls0RF/7XFFFSWavzaKharY0j+Yza
l98G82tfey5xhqa1vjfkMWl/FHsg3YOTzeCvaii27h6Vz2404dzW3gjgbahG+X+s
PRHz91+UTgGPHB+q58fZbFzmOeYkJK780qT1vJY4IZARlqxOrAD4FplDY3akShNu
/9ED3b1edFtO3GeUuf0g1KTOHCdIsYYg5iyi6uJ+2Gxo4IGEZtxSIVL4pqjMv/+a
rKiivFNEDn3pCgN/ozfUzGL68vwLsjkY4RaEn5KrE3aFXKR0X9bFNpBbVndbzk60
6CG7RiSvwuI3It4f2MFH3jtnC0cf3yIDEzbspk9vdlA8vhmM+Pn4hhzQS8dZbln2
UADIRIQDVSJDcBCarIelrCgGOoK4dtfEwBro2axK7vkvT26MSnJjHyGqA9iE/APr
nZIIsb+fOmf+Hb0KT9antLv9PjEsZxA76KXqj7Z3XFFIPykYszsP4gwdlqfTcAqH
5nNoPOGFIotohfmwHmVrQUPqPdu2NSslzk8Yi967w0IDA3JhyL+fn5fOhqYr10Uo
A1Som5UTTIaRwljtq+A7pn6NydxgZjNBO9PTyGCR20QDyNrygBhMxnDxvYi1fCVB
wRzax1n9lcugvIX0XJ+vIP/qDW92k34VAAZcP65HcN/hCH1HvwoNXYZ5tHRJPj+X
t4/rMfyp/mEvL92w7WYuW8HhYeaIzjO1aF9pRLt/jA1Ct5luQbfhf47FOCchqZzT
18cWkgHRFTZqlMsY0af76RcFHPxGqG/PMFZBo5y5VfSEfF7fLLydvwK0Vzd5JX0k
YHadHUkeYV9eE37H2bdPTYSO1jCUyl5xQRgWzKENCTJwK1Jds6FtZnw/yrKrpT1Q
2nLnPlC6Ene8CL/OXFMo3E4AEzDjJ7rlU//ADBok5aR+7cjYeZGxhA7XKbwNW3Er
RttrBclgwBgT0nS6O+bGVy7kP8kVlBOgHHfnWRocr1QAjfPNn53lQrDJAWjyvxsV
YRXdjc3sxCiNV/TKQI4N0SKI2xCQJP44OZ751ttGVfhf6dGMwsPKbKt+D48I8hCU
6C5VGI4CUf6l5FBKEn2xLTJeMEKjAg1ZzZtDQ2atUlL/Ubax/1hs0FZ6LVwfdYyx
/2Kb06ohVFhiChUc95Ljui5WTfs36F3VN5MibqQfxfQZexEyK16DD/zR4LQwILCE
WX3x7hVqUThw3P8r78SsZf4A58TcBiYQ7TdOIycn7aOZeQR8l49Lk67c/CsIBk4i
UcwTKr8ubBl3XT5bZ0NkOM/mqVBAe3e6vq2OVNe4KkE8IQ928D0f6Gl2RDaYdmEt
z9afQU+ZkUK3diE3GTmaxMTsJ1bikAEj+QztjQAvwuujUjytsiQliCbD40utG87y
Ltwah59K40Z96oVOnyXOmHUtBvIzwdp9uB+/mgNjqNFjPP0242Z7hbxZS21yNyDQ
UMopS0HQ7xZk8Ifu7zJMfR8Q5wI0976TlbVx6it5Aj5xudqmmXDPPd+Dlx9U4dJJ
v+rmUjMd+0hJ70Cuv7SruW/EsQ1HImDYZNDd6D3AgU+G+fy7VgtVPRg3J/yLsaMN
RhF77AYv5L+3nA8XzOUEUVnJXnWImmjLoLF451Z/PoRTXNoEA50Db3cjEDBakdEK
JJHr8zjBMPE526ki5dgEtDJv0EmqZUtlq2Swjbq5PRhLhbUv8doafYwyp+WHKQxI
vI/fpApmEKbGOkb9QT5cEY7Ug9pPKQ540RvGWrYxQG0Kq25gso9Pt460fEVkXRFf
y8wtsOvUFqfcgVJ0W8ItSopqw9siAx6enV4/YCF4ko+3IfjvPG4T3+GmLeVmQ/49
XYzja7Cx5YczI0L2xGcPu85rZpfh7Lv3lE/uXODDUYyNpDaxwXxEMaNi2XC5EEAv
QcyLYey4Ws3VUtMOjQpQSPvawTOPJyKEdAjMF3fJlT/ZmXO43jrX/qjNEFtZFYxr
uExYxTuQPST9XXBsp0878KGkpMXiFspZuNT/PNUD70D2fz8FyKPTJMLfPIN8Iq7W
NHsrHMArQjZs/Vn3b2WUSB3DdyYEhEVoPoo6YnfI+DItxyUQqbUWttsaaniru0EL
7CpkmWJqmq7p2U1PVlHI4RCcvL62mS+a/Rjzqlx/LVOiBoDIHmHmvYNakqrBqmQ5
OXaLgNgTqUBm2R8Mk1u5apQ9jRKkPJ1tl7Lk+l46oDTZmoXFbY+t3KCQy/EYpvta
7vN6ItPwYbcm/q0JcgrR5fdkOFcQ9our1UPaEmzTy3mASMnuGvZBlfUEGFz1iefX
RBG0oaCuEVHUe1LXxoVVb1jYkUPukSSyAK0GRIF6KcYSWhQJlfjk/suAKYAomYi0
mkrwT8cv46f/8F0cAbrMgxb0Gi+kWZKcfca1Ks7NoHlbnGBpFeiqTIBpaMM2yraf
omy9goadwz2Vx9X3xXl+7U5uzcMPgACZfDITFmIR5Lsi8lhsppwB1qfmJgG80i42
QqGwgC22ZMtq8hY3tKocinF4g4KSlkK0t5hJAeB2aZCAhVXtM92gIdFJfTCsWOkM
ecQTypckNQfB9sq8fajoYnbYbAMrAiEZ46gIrD/Ymr+TCE9EhEZr//myiO1QPx2l
YeJTmA4pgLfXIGvZDU/IBV5UKSj2ccDaPj7GjcxlgiQqiTazAVR9wN1b4kcjF9tE
jR97k1wcNUskPJU/qtbO150kkwryFO5zZi22rIxxoUKrTyMGLdhXxxFxAkkfHQ/E
hdiKP2aHjqQDrSH5XgeVX53mqaYduM4mHHV0hwUaJMI8x40gByD9sort2kp0BxTv
NW3qDwK2QQmSvRsng8OV5+DsX5S6L/eAWoURpGCWJr77JqKH69P6uKOIBWoT+g8a
alWdi/komlbs4XaacUG6DBKeX7mhD9ufuRNEe+uWPovfRaErRINQFy6cA2glfJDM
VBLirUZprdu2Q92TI0W1mSHt+C9vj/rGqNR7lccibe239Vy7Wp8cqdF+3O7GVTmk
a2KSRe/6REqnPKhz8aYtLpFX+ZZ1vLph31l9z6lW0qQHGCvIp7k4V5NXuy63aEgd
7+NPhPTZQ8I6x6cjbAxpfncmXN82aSlQtERvO66SUX1tu/vj9Or1zJdDf7SwRW/X
0SjLwSSCLnH3kiYoKMNWW6hFGt5mAmb+Pny4dmYs9p1vKN0ZparMN3syBVi4Uhdc
EwXIA6UTF4aQnzO8iURmhRglzi5Z70o7/9ZyRZnAwkAakux/8CMLzVnjWA3ktduT
91buAi8UU947+iWIkNMh3sleDb2O6v4NCSAqhZzdIBnbteNGcbW0UyewH0JxaqyO
auNzarjeqMvu5TKdyj6xhxhTCY2Au+WQuVT6Yjlednht3hHsomkIFXv0XjOnqLAK
B4OlK/TUnyVGemIfNMpP2K2TgpvkKxyVXczmNAzCHAVJlDZejvHdSKk1kMf9b0jw
SqkzLq+8kQ34RRCfzHd2V3tk9GLUSSX5dZHy2j90pUljhhBCrV6+m9+ji3J1zKSp
mBDUroHfLNEavZReDv1Y3kY979CIunjjGddR9ypm/PbDTSKxv/Gnc9xjimhJ/9J6
nAObPGTbk4NTUbBvnwYd7m6hCEAI+DTVtZO7bHHe1dybqI0MvJFQciSomTEoo/i8
ta3Ht7HOBbXH2c3NzCAAdN/C9lnRBXzHwBDVBHvEwM+UIMA1DONO3CNztDGChwyM
b6JggL6hkCGVfo7PIhtRdX8E/vBy0Usm6gKHJr8Wi8jWMZthTZCJB6+492jm0pbn
UyjcrIQjLdA3nGO0k0DQiRD17q0Vw1E3TjqEV94ihhmRp4c5x/GisBP7N5u0gXxs
iYGRgxFO+SgTL03HyXJ5zUkhOlwuxwjcCPyNkB3746pCMhLQ9AZv2/5zp6AowsAK
6Gh4jrT87XngDlexQ7X46fvHcGhFOBl7HuwzH1sfJDjGIfnQpnXgBawiBT8WMZsL
RWojre4z00gXp1p9E5LkGu3IGrAwqr6SMSvKUgsJhMwZ11xBZCUCF19UDc7JKy6O
1P08fSJXe2EGPZVqPcflEJHltfxPQfSUpoRlj1brNg2qq5ZiQDfCY9Fw55f8OWvR
a5Gp86zgtBpeRTx3ayV7VK5JCZBse3ZuKowC5AQ4GYltnMieWXvIAGMDApzcK9jG
DtW5qvr9t5LBi0K2Sgqq711B163S9Zm8MhH5dPxdhmcw9rKjca+w1zgZSTpxkBxZ
Ckm5BcjhasERhmXS/6Mxz/6AXDZgRiMKAGljRho00Wkec/J5lC2JSEwETcKNqFf2
x3bqjPtc9Sg4MTHpg5w+BAoq7Mr4HR5JvfPGRBBPO/9YoCVBPYeHPhQeYlASfmLV
InIZpsnoH+9sR5eQbnLDwgEZjDjoR0jo/syx45yOLpMygDeJKU8pVviGhGDkVTtV
+OKS5pAJ9K+NlKH87jDFyr2jCLwYUAoP++pjCcmJ+svxstEWh2f5H14Th/j/4gBm
HLgW3k2JXiKHAH4hm9FFXacoS0s13iCj6mszkz+Cqcvz1Vl03WXdKLQf+X/zah1H
+3fRzi0ZR+KBCCDko2+FOVYSFj/E9yQbEkXQUWr1gHcnjGgTyYcHaTMTLmqYwl1E
YxnOBffCwWcA4T0GTQa1aGoFMUXZygVJyFWwQpiyv5XQqQFSHWzwRfp/MNzCQIjn
UMCgypjBoFGl16rBamswy7DvnhqfYnfRe89U7LOy+RISc+NAgnP+wyEYnHT0mn0C
mDYdXRrZkrzE6eCCwapjQGfAunWUw5kNC4H8Q3R3DqE1bWm3KHOtMcevzWDup5/9
VP/sv1ESBJM798ZETLV17XNOcR+C86eqI9OKIas9QlgC+uYneb2bx6LzVEppriTQ
T3461vMjTtdwRrckg94/cY7ezKscbG0w0McgpJD+jrW4xsiwiv/kdIKDb6o7aEPe
c8r38NNwsnzKIkpz9FvVpg7eGgh5OOKfRcLfPZOCANj6h1Pw4PpboOB+Xyj/x6+I
v3BoiTgkLD1LyI22trrHsf8SIf7OmwhAGu8YwJxbY0a39vR6Q+p59ExibksQu8Vq
oXHZPLPTqpKXNK2QwQhnpeUpxp345/ubALUSKyXOgfKTmkYiwdUa+zptytv86//x
xY0ZzO0uub/MqDe+uq9Av8AAD+lnwLYTsO1PiJfVOAryo1kMHS94xYLjP4/i6SvK
h8fjaZpw+QK4HdQyTIFXsreguSSXBsg/5JXvFpiX610WBYlkvkq7j7fU9B9rwXPO
tUY+OwC3ty1BNWx5y5P+NI42px64waNfaaN1MUpQgSMl+FCx6s1phyx9Fziy1kg9
EblH847BLI3LGtR7XMjg/0Cie8igxzLScmpdPvpNmYF4D0/TR5RtmrC1SmgU+Gys
mCCZOzh6QemIBit91j2ayJfKXa9hOe6rA8BBBy0EL6k2UxoYIC1U5fghvypzwYg8
1pO3LzvHhqL4bM0RL/r+UiMh+QiAbrxlv5grgom4+/EDYH1I7AJ7LMsvm1nCwnV+
hb9+2hVFfnKErtrXlyzapK83u3XVFf55DfT6J5oaQOhOPherYfdAJOLjII5gViiT
3e2/DgcOepFF1vuufHjQGMLwXPfUq/WW2Sy6rpZljurJbHlD4Ty+QLcTqA/YyBHu
UhuvxcCe5rVYKZ6P52kTJ86SOPJVpJozs6uVd8q2YP3tI9bIr5uUbD2ln7FNP3Nn
afh9SjBJeNmXgO48PwHcxWSg/5tOEemSVRm6QvxaP77DUE6tIjo/3SmmPjF91vb1
JN8hWR+ezLfk3tMlxKn+7rtiX+UmWYMqDP+XPT6/KF/LP388xgFVP9B+aenRMAcf
nVLZ5Po6tCHMVY+xnThmlRBXmTUOdaogv/U0yMJq4CPweowOXXKlU6vX8svpVOjK
P/oVbDEqRBVmYha6D72nTb23Itaeuh/vrYfJZRFGW3U4cKdhusc3qnhMFUSsamxd
uH4FdasbWQfcnjLh1thvsKa8Ve2XkQ7GWpTPZZZYUqfvGYmwVDKqwkIKd06dM/G4
QyMja3nmm6WUiorogeje0LAG7D6fQFLcA5s7PbDS4GOK/zTwhH0DgUzIKSOGlf6J
H25viEygZ+RTU86xgWO2mLZj0tGSaHnG6ni5nObfekJ5yCQeygGz1j7qNoGS7fth
kZXUmri5f779NFyWl4XqU2/XYYmPYv9uq1p3lYzb45FwbtCt+kQDiZqNDCCbLLGe
SBdJ5gxGrF0oqABZGfRatP2b4/AOvm87OwtQ64H9AtEmAdjJ+cNSTFtCw9/ZD43V
bHPFKdhfVifJB3X5zACrkAy8Zpy3fIGlF6gQoDH5W49eIEw/RKZ0Ugog/feLA10v
m+l7meG9yxIzSoLt0cf8Wwy5OinVVRZ+l9lDnRCgpVW3yzWe6X8y+/hpcdAzE/Gt
gnA7BQWylmYMQfKnnuMjQRpGTQdQ3qEXuOImQZ4FJeCo1R4Okr5a1cmYQYGyC1tv
OgwJME3kygH0wFmiTO6ZpmATK64no3YhndmvbgR+T9/WHfhcH6ZCQJn3ETEQVho7
1bMYs0qNUjNz2xlAtAMkWlCVcSUffQZIFa5KA+CaX+vbIFOfLzLY1tjO1UXwk8ac
MFR3qsOHNVo45wKKAA0XSSCxHXts95RRhxiYVYZtLz2lPb7lPpOJA3174b8uI+01
lTnseEiPj1/JO5v/Ds9tdoqVoPATpsNR3VRKzPmnBKCGrDEZQUQNbp5ZlL0OM5Nb
N3e66Nm3T26ur1cKwApB7QNXopL2LBHms1QYPX3x0Byhq869Ol4IbPmIC3GwfwJt
SqqaI8Bi9vlZ2TLpxUa2u3XEP+awwmenH/3i9BU5ckEfzoucw+pEf/sF0ydpJMQA
mG232f6OO8f+qFPaxYNNQh2nXuYzSYhWtJpsjtw8ht5H2kZ3erGIci5nfqV3F/4e
sBkiVeLHOi0duYHrE2ODe9CADzccHfs+TpkvB6C0GnbNSV2kPRYTws7GAJQfaXI0
1Ba9caAJaVnDRGHerLNuSfH/wEY9hWmJbi58CLHOMp5y0wcnUWEDaTbKm4Zt1WtJ
2gTL4nS5N3zO+8II8+BBZj6wMGewj9HvqhgCa3NgwnhvkD6qPnAp2jNnB3iSCUNC
MYS3+JKh9uAXgcrBMSaTZoE25JVcPrct+4nMC5rZVpjgOSZQsa+3W0ixW06YtEEN
Fjj+fKAI3zv7uhIyLo4WfHLVS3lWNrSoBntgZRFeZFfya0rzcWfNbat7D2ZH5wTf
uT9mou3ADKUFcok65XjrWI3RNEL7pEq5OvYoaedtDBwR6IiIsIhqobnvdJCyOyJz
8cdmphnGaAYRNlkQq0EVGgUM+QI5+QdanOVHD++4Oz9BBluselHaoLY/mzOxEQ3N
6a3fWSdQzKl0+lXCLyMmg2OiGxo+GgTAHXuwNMx6mssYNd0XszkEB4ToX6cJPFCx
ODiF1suklS7rNBsKZkPBc+q+g8vO8gifuaZ4fgwcRsuAKMPcQ2cRaWMWc+lscxGJ
Pp0Rkfu/vwkLjnjm4gND+fcBcXj9Pnmxk9XAKRzESneKlitDL8oXVL+tYGqypsQb
SQ6F1ZlqMzNPscY1oZkDrQCbcfg39e9qDuqJbK3SMOiIxoWjaTcicMUoszQE0HmY
vxH/MTFsdwan3pkI2fcVh4ulXqfoO/ERATIcbNp1KS7ff4b8rBBQIPswLeCvZU1l
DOBntPEU/PaLwJSJjfrN3GcuR8X1S96ri09XqR3Wu5pbNI1jKYHMNyfFRDYqR1DH
BzdeuAPb/Hjl/9I3ttnv9FrL4GYTK9zswwvazNv+Dt3n7TA5zeiLMAd1AASb9rFJ
mAbtN3/+EWSJFmJ1Wmi5b6Ys3jF/NSXN0jGRkw9LGq9OBhw2/hB8yvDK4wqYbr+/
MjTpjKp5XkVehhCBIzr1nj7uhB8IVnxK4J38hC3hmePTzKSVPI9zst5n2UzuMVs4
hkxaW6HrbkYQw+MblrghKzHuYM/W158Z9oqX0y0okStEU2lkWwnQsmRYSsg2dsUQ
644ncfInru/m93a62A/2GK2Wc4BlRRgwFjg+KXmKL0vjYtH0VlHvSk7Vr96qDPCB
C1GmkKr8RzWcObb9ipyrXMM/Yuxf/cjc+Y702UgGhfI5yoU8lmwMRAE4EVP+NOA6
rRELy0YFVLlmm/47duyQ493JXCWFevSrHaNIWf3Ybj+rkLNQ3ZwmJSqTIObhWcUZ
nYEUN9NvT1STIWqMYSFsh3UhaGk7eL6jzuFrBcxLDMAI1By/I6Faob+1GcnQ9XMZ
jHcZZPcB+SxlEB/FQm+4vfn1Et0pHXgNJb2eCGB+hctm6/7ZCKZHDqvsG2PcoaKP
VWq+gjMgp7bzFvzL866wDp8c5DRXVDc7oX/l5lYim5XTUn534gX2pQQ7PjiDHDSf
7iN2ekUaY/YaEWMkqZ4DgXvXJaT/L+e4GyyIHB6xYT+CaRPtyEko2ff35Y3J+c4D
1xcXhK+/FCPz6IlmM9ONotTnRtr8+U8dgn0CVGb2tsffFRaAPByW0D3og31hB13W
lqoE8EFzvrQCNgBzR6w1bqN1NMMg+S/5foWw4b2DH4aMy5BnQxUPdD9Uhhu/mwr1
0X7wB77e/aWXnqKvo14Xk5PXeCtwHm2IvTFQcT2kP8dNCvnyJM4v05YErMEN7XlR
m0QEbMth4815wX/nWcFn2bSmqNsYc7UE444tdAxOGwCdL2kuqLGyVMkvYIh6Oe/x
8X8WhedIJH2kFv5M95LT/UshELrILNwYY5C5koi6spIw5ELvPPOWD+EiA2KDhcg3
OTqnr4tWLb8CVpMmfQfJkgPkCdc2wPVHCFu/aE20SzueINwUdJWthFmJxZGT8N0y
VmNI6lhxY7p4VaxC7/S31d1klcFObP8CRxBoB7wF4OmQFyLcR7Vvqey7ZTvjw0EG
amdMw+nYIhph2b0Eo4nW+z8AZJh9QgQ0glTQyznsMHwhRQqka20VZsTYb90wXvPJ
exIhV3ehg/mJnVnx7FaRGgEZQwmFR7t+/gBX2ZGJcS+V1MDp5AcWzyDEwNkuRa/w
YX9eTMKYxHJzibtF2etU16bYuULQGxu+qCrdtcQQpITbOCQE7uXZ3KUgypcVkk/k
AVs8tFo4T6UTGY1T0wqKgHRkfkQC3BsJpe1tUHe1Lc2b5LbXoD5fF09xp13xTAEK
SbI9if/Ig1K35Cg8DCEBe05VG7L6N5H021pTr0zXBMckyzNl/XqUGJqNNwB/U2sV
oef0y21MKSE01o2Ni1ZmBL06A6k2xAoSQj+1/FP56DUwXXmGTfY0P68wjQTqVJZJ
p9x8Fnm+fUUCQK9JhNVoDrrgCUPbM6p03/XyaNA6FotcCDiVjTypJwqu1RaA6iCl
ugnAWvBQ2gu1GSaRZbXCzvzPZ0uL3ZBGzw7txxj8FcMuPZd1h2sjWewjLTK2vTzi
MYZgzQLl+qvlzbrxUq/FeM5zl7DXdsM4V0ZjX502afY6dyQH7I6Hnd2WTwAtPNVS
gtuczDwkSkfDOa63yWWk50YsYAlvwp6r0fwO24N62629slaJ+jr6oexqSXOZJ9l3
MGJQt4J8lX6Z9ZqDzASAr/SisOYr8Yryi4zmmrYV1vbrgRaGjpSX0ZKrRo4l41BK
cV5PNMNEHtmO8e76ujkYyE6QW0Q8dWXb8Pf5O2wybxw5ICycM061LZ6l9GCRdo+q
4qsBrs390l+QjqC69+qMPaotD7+wchftkCzIox03jSUGoPlqlgaK0w/Uzmgk2V+J
A8mZ8eUMbFr+aaUw+KVMwaxW2XFEtX+shbWg0bGgyFSOnp3J0ftLnWJs3NYn4tiI
7nRd4hUFTSgD3m5VXJySap46DqPSdcsftp6mPxaZjiw55WsSXBwN0gBbH5jFknjB
1sa/bjIKPYtK+hEMQP2HDiKm3I1iSF+pcQVVKpMfRC6fAlcQOuHstn70nw9YVVYj
UBh4WE2cSu99kgV1FJPE0g9FT6orhAKdK+gSFAdfygSX7lB3HCOYsHbgdVwkWej0
qOQQXsHJ2kQrl6Y9cYS70sj3e00oowyX1kjuE+g4gwogPI0Gs0kVGZ0sLnoDxS5w
BP/ph+N29Q8VyP/wNccmJlBylbbYFOGcjbn/7NXGuWTPEeMSSuPnLrLiFi0OCQlF
QX36Mkc//w2ZbIWHppd4jqedT1Uv8KU++tV8khy063A9j9cwCxDv30Apg+dZjqii
4Sh574yabc5piTvtIGayfpIchQ4rhJ5mCqdO6Hr1OG3DeNVzv82R60KPaxcUEzH1
EPP/QeoZU5KpAsJ5j7pnKuLb6TvCkI0OOYLHlfkktwR26NwjdJDd8l4Rg1A0j32Q
JVdk9MIWXHOqcaH7LacOs4DKmayQYOYaEXWMz6JpuBZRf5NMtHCVxZsOVouAUm/I
CYz9r/N5Awk3lWpIJOKPoI+fwchiaSHHT+Oesy8rNuJ+Km/Qs0OtS061/o23d4XQ
jBNPeMgq48923o6pAT6SxF+Rm5kuaS4KLb/S8FNO9DTMnbM5uDwI1HECMkgKrRGO
tLvpZi0f/WaXzVF6j6KGrOK5rWKTpLhbiqwpZXaNO9RExUUtwTaGUYX/z+iTDRxH
mjgMjQwbIe3r10PS4yLzt6t/JAYg06R4YaE9BKkRAO5VODIDQZp6fAiNpaNOmUjg
JWIsaXGH00g0y9Nwppa7y7a1+cj7QVNihOg9wpzoXed61XDCQUUGahyX3SInLXy0
8bftR+4uGAsKAlBM7shR7GD6xYZMy/2UzBzitkHhv1wtAle7gz/mZXnPM9pSX/um
gZ7hzWTduaLLjXa4M5Tu8AJ5qdsCkbEhPtFzIL3ylYSZflDPZMAsKIvBB8TrCzUQ
RdHCQdPTHXO0BPEmQzc3Z52sxPWLXRzsF6GxjPTEAlr8EbbBQoR2MlQ5j13u6wFw
+gDXPIL8JAlx/L9MVhu1GMLyK8j+xf9u//z+HurX58Zdxe2t/N8ZVFkLT77Xt0C1
G08+v9hJaPdYGXLwgo7XOnkwLFeJHexejdunVvousBpFehVeiWNAxbJHUXSdc4N5
67xtotvHWGyG8fsFgex8/CjrgAjyccNoIxEakQZ4QozRAZykSuF51u/6dcTLaNn+
HZHkk5cehhylvP0ENEasVe3gaSzto6KmoO/gljWuyjgb6ataZplm0rK85mtda7/J
59uxmF2e8/fKaB8GgPvLATEvqknqJYkx+tbECyc02AWURYr6pyZIyCdCgHsscTEX
+ZjCfEN1yL0flolf0DYJ+7cuwjRVvWV4LjaOjywawqU1K7iSV/PUxfyI7xfLeQfn
qd/JZn8o7q9hLQ9i8i5ih/QaH+PMB0ZIB0HpKYrt4RpKuaK7U2blf1crU6+FBdhA
gTASEBbpvmkp0ubN0wBxsasbRwku6DB/xc3pMSCMUiJwl3rTiwL7cd2aAjV1XSxV
JMHNoyKrnsyCFtq60DEv0T43eyJI0Dz8Tzb6Z6VicL53jTeTM5hNE/8XFE8eiV8N
2oOAW90gFTuD5s/KCi97H/FArkbQJUtpc66qgEA0YAPy9kV+Q60iMgqZIQ1JYi9J
8c9S1MwqRMhAgx18+ZckaoYm6qorfDZvAABJEHIe5cKu1JbcAnk9yaq6GXICq8tb
wSqHz1eUkYSXyBYPxL/D9RK1WU8SWrm6TRwL+MfnCUpGta+fPtnKEphmumNW8r4A
h/tx51bI5OgZdiuxdY3kLknQQlFpr40/JGg6cbOAaNGScwEyyXtS/ZAkM3h8v1x1
tD0fR1xgxPJW8eF+evsk4iEyP19ml3hYaz/3SezDPsK7RgN0FtpmCcK/IKujOKqy
GZqKn14yqYUSLgaDoTshgrIuUuAUrpElBbeQiWeEKl/+nKSHKcQvdMt7lRb/VjGR
Ys7+Gw1a7vsPXnAivxh8n9jOgQUftgMBSIUv7+CEuepuXyJVWvWmnNJe4Ahc4aAd
QpnbYk2i4HlwWJlmRAKzkxN7cKcj43q8KVL9I7xqW6dmxxPW4CnkYjSe9U8sha74
sDspGgqxnQeSTqu51PdhtPvVoNKEG/fagRYUj6JjNVR2dqu66fhLxPepti3zX4i7
8ASfDQEGcpJQmqriQUmL8QsHJ11fgrCuHxzN/t8hlkjEpw2CWTzQDj3GqdTyQw4h
yVzwYVzu+wAhjpy2auTxwrgv40+zDpAh+8hnOuMSBXhCsWpQ60zPnnuP6owtHIRu
UYPmr1MgvN87YxMvQTyve2xyRLtIRZ9D8RYAcdpUpQxmfutdygL4s/aKmgD4p9kZ
jR7AONn69MDXxco/VkeSulWecNl2tHcvewyJQrIh27rKsZl8fM+C6VStuY4CAMqu
4WXdAzyAWLl8pILerGvGKdGQxYWe1b/NSKdrtsyeJb35v21yHtIrGmgWVbl5wz1O
AJcPtm47Ey4pOquOze0tr4sP+NwbQNClKBMpetV/7Fucxq/q+zMfa5IE0QNrePcR
2V2OsxUR2jIqHjJx00qPV/VCwYd1gkT8H7DzdURo5j3TvQNvgqp/3Mk+j/EtDi0j
e9jigWMQNEFX1fA0wz0TSoFK1kQ6yDACe8qFjuZ4ocl5SBVdbXfBBiDm/EAbMDu0
3CTmov6ZYYEbGfcmH5frsdh5izV7qWDq/I8zoQLIwzIBjG2CNsqpR8fc0CHoy9N8
MoHX0qXA96AUbw+/IoyWPRNfdQeCyBhUIm22g8zkyCq3rQ8N/OCqGN0Bj6Z8ia5f
WH539iFicgpXVQhxwnd8kpBy97pW8fhD/no+OjRhNc6is7SzFgfmETSDmymIaZj0
A1a05CvOzQv8mKlCHXSZ+Go4kDazc0ca2kSMd1nRM7XYazRsYooXXn0lidqpFP5U
lJIUFfVW9XJ2PWiYbVHNtkXkhcQbt6aG/dWoK2E449a50xRXACJSRvasZGxphr/n
T4OnFSNGo5HGvKMSgmTiAmZRKxNapXi5MaeK/87ngvAxKTrrbJGn0d0d7h96w40l
fjq0Pk5xgGuRl6QBQiE3YRoAu1Nxhe9DlNEcAi4cW1/4gKCAjwvuiIee/7QXq1wK
vxmoPOwyErD9qn54gWw4EY2Ckx4LRm7Dmfsb+HWrJBPkKU90mp8ojkRcKQcz0yGE
V2BeLFjULFb3n5pK6BFE71lmEQ1lW34TLl82MDhkh8s4df6Y8+TwKbCkth5Qxxx2
pKW/0X2oTNXpFQsxWyinW/dCs0QISzFTKj/6C/wwHvv6+TpArxmEReOXNPxlzVlh
n3zwHAQofyPzRjVAqHVVWKgB1DzQfPuYAaPW+M3vEJ3STIEwuhKvyEq703yEmloD
OqK7AsA93pnHoO8WXZpeXrgJlyqDbhLx3jxNpR5tH033hkqrPe2g8o059E12rh2C
XGk+1TfBSSSEjTWT7xRbLO65+kPtXvdiiDve6oxDNrSv63RLaLgbOgUaB/6qYnB4
oH6wBmAV6q2I7bOd2Ez0+oBuMc9hT6U4J5/ZmCfNQQ/nvK/XUmqfxEEujgvL4Z7H
rGvMW+DCSzhsQ4hDCxFAiCgSQ+5biymQXrL3n72sRvuRHpAac1ZHSF+xzvUG7LBx
fp2x3/kKcn7qiEqX9Y6aLOAgEhxT5dxszMS6vtGGGFlfzVc2ZvRMifAB6W9F1Qg8
729LY7ZJ9T6E+cpoHeViS9Or3/q5ru4HWqnNPU4JyqfYsxmmRhB8YqtsdnfvJRTA
dklcpEf4/g37gw3FJAUkHk4ZNibHWsQqi/36InnBzKXi/jNovtYvtPyrY15BmAmo
13r8XR5ImZ48wNR6BAKZOvFPd5tLFPbqkgHIRZkXyUDzMWQD0hcbdl8kjbhDgCmb
CUeSnBe9EnXu+cDwhmkjTFpQyQdS3skFkoTUIS7OPSbD4Cb0Ulh6GT8VJoagM/xs
794dfPb4ZSm9KlbC/HA8FckfoUcNgL8eDsZ84DNHV4kmYmbb7qcShUUZ2hLcbaXA
sBpjNoPzQn8IKw7iuaZ8k/TpIc3Yc9rfDO55yNG4TxXTQsZtNsFOqP+O3Ok6ym5G
+KMyH6rCkOjWx0Fw2Ob0HDEbr73sJMw/kYfL9hFmu+nVxm26OqaAuwbImye9dwnk
PzfPuvRmchmPxE+xsbxL/GQyW7lWI3yvQm5iWTKfisI2YGIaZVcIeokfqL53n52v
aYshPI55ehkyWPbHTnLpJWxdjupJL7XyBhWNMLus48FjhY2D3UvUuNfLoQ/9Y08U
LYmm2JMSGGobA250lkvuLvCaREMjJvHbOmk2wuhIfguzfj5g1iMz/cSs8By4TiJ6
poCW8Ijtp+ngQ+q4Lv/SujKHRIFbVMhjifSYvlEVTnUHleUFcZLd+Unaxq07Q8Jm
61p/6p/+XW00vqzmv7ndtLqRf1GfB9+x83xwCRi3JLuP6xtO42e1piqMS/zxQZz0
Rhe+aGDjNVetCUPT2uPHt8wWvwhUCTXNc63eJf0XDZB/DrieYtgZZ0FjlCHhX3hc
w5UjeOb0CyjF6VotkPbPweTqGfoSgghPXTIeyguO7lgew6H4Oq40gh4NHTni1LHM
zWRBZcyXEHmonxycJ9scfcs2oFuZfbSEDRfePlDwqp50ogrxclOX9kHPCJmRQ/vR
CYavH+Qkc+dvlJ3y+/WDgct8KXtMUL5CtjKuFk56zvGhbrfAa4dhg78Oo6QJ+Elt
Rl3c0+9KxcnYfTztzayb17r54pfmHwxDn1vxHLZmf7/UxhXmEsDE14Wi8Iqa1ors
e799CsgZp62EeqVTquKoEGYYYRGfDnhiLRziI99M9gjLwZCEMgvn6TybXoFsJ8g9
Ya1MOpM+u2T8Upzhj4fd6pZ5lA//GCR+79BWm1GqGfC3Ip2bmwnHQXJRSxiu/JgV
g/lP4f4ZzsA+SOww3VRxnsne7LIs+NoF95EE+lwxffTPcrmYYFpY/WQlUOeEac0T
lS9GtAJuYZOGuKjQos9IiDyF2P2S2vjXCI7ugEmpxEhtMfwtT49XEdD7FSXv3gr8
jQotVtJsX/zcBddhL+KAIK5TPtkwF5mbEoS4dmmprgtflIj2sqXWigk0FSZiBO+8
8mNl//h70Dkdu2Ho6qpEeiRyncXz+SoUG7/D6bkG1l3RpYKHJkSXBNh1X4l60L3O
+1BkzEDIuHHShwd+FV3WGJ3o2T+q2wUj8hmEpw9BdnSkxrOBkUxC5Df1T5Kwk1PY
gQByxG2wHzlKY7/zkjv7EvPcUmC5Ar0/c21QSSq66U9on4bRPBgLu5tIzlx8HKaa
/a66rxNKPTQV/jqPPhSI/srzmQ713fkv3ZV6bA/c6Y0WyUPxgaSJHhSGsJ63dsTA
cA3Zw7lI89NQuHi9EUhNiRcz6JXjf7iW3BcNHjiTEHC3Nxj5psLSu7nMVMZsrvLS
6Rt0V+DVOyRQB1oknEfiHVZHgsI/wIX+SfyjtE3kTFfj/CDI2Poz7N+hXx7jvgco
CMiCZVOP9ILOIoTPbwvjwoFtZQx4IbUINTQU5DQnb476kmCiaYnQvcboIEy07z9i
J6Iz8dEjt5rO0wzEeu0/P3AfEAwGlaTekuFPeUWXTdJpDjrA9iKBkH2eCjHhQxCz
+Fm1Juzf9xFqUVSPwnPDFjLVXqJQRcYr1F3jrQxK20zwRnv6V4DyQNWDWRGLCLmg
scLqG0rx40ITT1lkiAQA6lL1Bj0Pib92hchCNZkKeTguncDuJdKJogv+Dh5i4acd
OnoTFn51+5zXNidoQ40YEJMlHoMjpOupf0cHNaZc7xLIynMns2Fh+Jd+wMATafwC
xQc6UwRKTt3S//Cifvu9Q3Fsag1myQZ3yAUjjnwrJAgaWMGFCDkf/hbtfTy3lXE9
gyeGY/cDTRWlUc6FFUvTjjzdC/PJWrfuYiZQAiNmPoo/wjY/FGtqI/UkzQOw2xGl
A54l9/cswmXf283MzJs/BXPsqUptrWtL5Mc6gGvUUbixLC6Bb4HpLa8ZfAY95tpp
m1slx6cDqEuFqIQkOFlP3/0mscD0i447d1gAcNpxuUP/zqadA0+1QdB6W2lEBnUS
GvwcnlxBXevY7oL1ss7UDtZmoKBvG7QrINoZqdJ/2R8awSDC9gw/HVMVfTfsRbXF
AEKbvpc/255jvbuZt3MqOU2d9xhMm4bWeWABUdSiRWF0PU/fNtU1aHDIC2DoJgVr
Vox/eZF/FfT1/zF1JX7/gLRFSQX9z4bdxq34thPvSPajzW4Sz287DTilP5gcMBuS
U8a9RwKtNtjOmYya4aVaoEcys/hJtptxnJpa0axEDeIAzGEU77MLuJX/FoWudZSW
zAcZHheZdNwNNqY+QJStAGcgVNNkvPwMlTfqWc4UQNnm1MRq2SUSCK/WXdWb1jVV
PQoxDoTBOn2JApDNTfOTsbRrQp1gQptlmZZwuG5peNm8mjnYg5tADSAVrpX9VPTV
2+l6w1p2csf7LPIRqMu8DJ+XJ6J0JY9sH3T/SlKmQ/lbrrkj4jcX3dQenyYx7APh
xLxD8akoXEglKKLRa6lk2P1uC58KBauKYTrkRmcSE9OZtS5VSaTQkfqMyifkSDi/
6YV9wCbz0EVGInOeRBlm+Ee4N55gOwDpoQDZzQlYNK5EbGGI1FrsV38dPFixiMlG
vrwSN3/hWULhzKWnjDd19FBKVwn3ipvi4DZGdH71DkrdInrxwUC0ghFZdWO5+HKk
2NUs9lqWW6YH1DAZLzSMdssmnEMhSbQJTQ2dwbrIX7sVxMmfbWKCb1EIGGwSyBnm
oQa6APMCgysJejPJae4gYhc6JMv8JhISFgq5T9fS6sjKd/uyFpiYOKaoFJOdbW6K
8eqtJYgqforeXsDf21QjfH8Lgm0wDUm07wZUk2jCl5JlCGRaZRzRFdBrZpTMUtQY
K6r/3090w8WFt4vDJTFeljeXjvM3K8yZYMvYdzFBXJy6wQN9I8FmpgJYngq3j4gK
Za3XjFuf197ma29XtzJ0KTfx0j3SZPKdt6U3OBt3Z1yqEntA9HP4PtNKcG6RT7Mo
S5dO8ra9WYmmpIOiTBOh7M3gnwnOWMdqISm6rIKAYi6WMoR3E0OSf9FhbXqdA/Rt
z/C5ky9u6b+yCMifHSRNp8O52o5F8E2bsFEnCbsf0i+IqThYMm+WeAfiIsHZByQb
BMXCwK+08tdxKdGlya0/dr1+sVY3wPRAuqk8pkPODp7gOO0pXXdrOdMhSTuLkiNh
Phe9EwFMHma0F+FW5OM8Z/plmEk36zYha+wP0mZzOHrsDOsoHmxZgBaVNIZcCcKD
ehWI8EqdmGunPbzuyVQkNJzCkqAEevKqSoXRN0g4GG0mBxjG1QxZO4ygp42eht7f
Opf7+fI6HAECCGYcEliyrTV4mgsrv3/0FqVrMc0HtpGDbUNoPyPzuWFCCihjwttW
oJYlsMI/5Gc0cDwAzzYK/O4CSDYvrWx4JcNicYlCVr05MutesFG01Sy3EkR8vaEb
wj0VA7+iDbVkL4vUR4UMVsRqBJMpWRpLNUEdl+IFiyYwx+WCuLtqCk/gP/5Xr+sd
Duu7FTVa8f17HycG6IBnMTdxvt7rDVaKbNQLUwVtHyimBu4Yb1YwGGDOB+orRuEi
1sOxe8tADDD0wDwgtXCryuks76+FUP8s829o5QEZLCUrGz9u4JUc5VJGV3rmrZrQ
94LoRImKtmFPTAariZrvgUssotbkfkn9sFlHJGyl6kzRNke4DqIDGJ474JJUTma+
IVbFowPGBelVCzHQaH7NdVDkZlf2Kn57BtxbrrcQ9PxV193EsTq7lFl0LpObl9js
gdDEFm0fhehEtpNk6BGDRXjtaQOyqAqowvCgkLRmxYNhhrASAp+p4byXP4X4XXVN
Yc86GfA4xqQhUgjoSlDJiFMbOKs+R57WvjtRBxEZA6QzYlpci1+sccxcK25IHWqv
BxryhN6jK8KIOEEPVP7x0MQHOY/NEnIPV5EMTVTw6AoX+TKsXw9ylKYJCyHjB+3D
iaFHDjCTb4fJb0juN+iVqAVngqRg6evH9h6CKj0In8IHN4+Gy83lz1cNVTxdKCzK
U7mVse8jNhVRxX+cE5T3rM60Z2sG3o2rrUJdfJELM3s0rqAJNWQvta5n0UsHF0Yw
zTgdik/wJ4fwc983JTgERC0GJdyjjnrBy5xQGKSEHpjhh57d6Ku0dHW6DuhtCg7m
+z8N+1F2BR5bYQAaBnfp24HJP3ToDKxMLXLSajvoQutM4DEtA+7nbxur+C2lVLf0
npn2cJOXVY1bSFdYLGsf5KVNkVf/5uoVGsr6/SPspoGB3OzDRTR4/FrpFb8YiJ1d
MDgT5+OFiH8ECxd2EwEDy7n3l7u9YwQ1m7im3ZscPM8XSQoXINczqKa0KORpGupT
Or84MYMeleYjbDyWpdeWDbhfUoPVmC3gb/DuvkbbMhD844s8zyRSt9NK8TSmoCbY
1ByWA3iiXBlXcf/hvFu68IJYXaZ40IIV25m94u9xjRcWK4jY95FRxMpbJ27Cfk4D
M/rpW4U6hoNGMeQRnWgwHyOHlYVjQquY3LTj1uKgbcauXVdXPPqQ3DZoeRx0wrRH
w238ApUmap9+6q9m9T05kvedNLkzrd8Jz97NbFfTr0R1bXKMjlU+lmObDxP+fkER
4UhSI/taS+107/T3fHZqhSJorobHJMRjCJ9+BoeBohNUAyrbeg3GbD+kT/vjItKw
t9Q4fU5xewHAQGtcgacgUkXFTNXGC6oeArMhQ/fnXfEwe0DiOkKe4Z1qUprBF3CH
isB8U7LigLGXH1olR5EAr46FHdOz957wrDyuV8lu8lZjClZigXkLuVCo+EdJQ1NZ
WRQyj3yz1jfvIZIxT+0bVu9Z4Pe/1vO90ZZhmL311+T/pn0Aezoq7EO+ZPNLu8ip
crMnYHkjXF3ihT9adMzDCAg5qWAetmiixq/XF+ACPfAtw17N9M4z/CcR+Jht+XWa
h/1pcvz5E/mAqsp+WW7QS1ct9dhxHeZ+xaL0f6Rof3znZT1/b7uo3JoJGr90Sea5
oK5aScijPHXqMZCpARn5bB5VBeeNQoFchquLz11Hec+KsfamfBWmAOEU1Ztcneq6
o0oKQ5Ep0tQSBgJ3/0pwu26pSS36Lq+pIysiX+gRCJBzxCAAnGxSS3ZC5mZNX9v3
WqndGNZC7StqRsKJYKbMofMBP8d/7rI3vSEPwNy0C7aTU8+DWT2Ll8OsF+fEe0SR
sobLVHN6v7WjdZL+kQOCdhV79sOCuyIhE8VJAk9Bx4H8LBFTC0t3j5vxRPak6Hfj
HJsiZft1PDSzjAdyNi2J5PPC4cX8FU0sr5dZ+jb8auy5H3YnKoBdkWDLQ46PqDJI
G65doUfPXvZHDYkLOFg0AvcbIxIU7/OY/NiSf2xKLbLoANWufW+P7tNCKLz9Uo0w
ZL6KfVsynrISR0PM4MjDFBHt+e4Jl3qVX6LMVOdNYBqNMgN2jy8gZEz+Smwqo8sY
GAQAlZKzdIbdYos/T+Mrgw1lizwqisBi6oGF2hX76A51oMdTX8tes6LFffRRaD8Q
zzSkb0S0IT6rT7JCSqIRJ095m1hOHSfWS2USj2ZA9qqANVfxk7VUh0ZMnECJ8/2d
l6fH4F+/Qgv3GWO+JUuUt8qpT+ebBfM31l/nZywvpzHS/j75ygrpY0M6JO3d6ifU
A4pew7WpfwUAmBHydrOYQZrr4ha0gorsNkgNz0FIlrlXNGNMRJeGHUM2K3R4tyLX
xakyy17TV0tJJRSg43rKtby2o8qDGYdIOyvjaMOzs33LR+3qCRGovSVHDMJ/tQkV
44Vr0zTan4ab+R9TVDAkck9W2xMqoUyITWA7QQsyZOXtHK65+edYHI1SEniy9Jr8
Qv3jGZHCEvWFsmsX0FYpuCxVqo4/xcGh0NG8+ZXLAD8wS1Onw8/+GUggSUplHy5+
iBfoyQqiiqdZoZCUrF5/Euhjms7PnF+kMO4pga0qNuNREcuyuGw0ABbXHlbEgVgb
PPVFwH5658Tr/YzjXTzQktmPc++nJpiw8zl4UpQ77KKglX+1aHrqlpU0eaNMJMZz
GHvY2/lT/O6FH+EV2LCqo9FHuU9ETWJvofHCZeIkCFKiX4WRIJYKbQvc+B5gxY81
erwTLxGbHZkwpiOeDy9X8N0XuaLfEM4sA9rF/b2h3w6iMBVpfBYDCiFz1cajUx7T
XuhrPzSCMjI1+HB6pqF4eUEPeP0NXW4knHFSLvGtdpAJIEr3FD6K+qmlL5dvvLJN
rrKxcd+Q9zIK+b6O1v1EPmf3lfCuQ/EefjNbk9x7YklAr1UeJkeV7XfjsK03Idfm
GSQZ2t8s9EOAxyOmWKsLVVe3APpX+MNB6wL8lrGWx0W9PgsFh7NfmTO/CHmEHaK1
XYrYKCgcmly2vZHBNh3SWbqPeyMmYS140d5gRmgeemr4022nsjhAFsjf0gcQwzqT
P4dtXrTU718rjjO2OCfUbyD1Z5zKOTMDdOnx44LUnoegyF8QGNsEP6sVcDSbjnHH
5m+Z4HypRPrccNq7X6m6b+gj+yQgFnucBJwdRgIBYwwtDqZb6nr0y28bPDLDhyUp
IIJladmMdTp0orULrYkdaabXwJoK7iMthmGWNOZT3s/W+oehHQPPApF3T7wEKs7L
nikT/nLWwa2IRURsHL1sJfdQlm6/Cf4Rt9JFHz/rKR7rMQffVb/cs4uALnQWS9NE
0yXuurrqOAsYxNVopuzXea194FE2WYUJpqPVBUwd0WDuaUNGQxfRSmUBnejxETix
tV2dUPR1HCek3LiUgh4w4hnD1exPw7rPzYa1J72doEzhIhc7IdyflNyU983t6kNZ
CRvhqIpu/yZiFJ34suzTgzSKXJJxmF5KsxlvXRAsbWY4i73ZtddQlrjfJ6+jLAc5
bCs8aV3iOu1tP5BsryVrzmKFLKeqY+brtyESnB0CrhN0ZiO0hNKGNZyvQ/y1NYLy
4Z0xruXJq9RdTeEWApV1kd1MMJxzyRodeIRe7oUh8n0S+DwI+rmwOHEj3tSjDXWz
X0RezutlUpqflG3spARfc6fQPzBFmI0zon0sqVy9mf2pEmGPSQpEfqVc9DipQe23
VrwfaO2XzI+z6/JQbbK5IiE0L1qhXeVl4DBprDhuHJBnO4N55m+QkmF/8dsM/kYO
Bk2cPyKhoAve9z5OVsXPmHXabuMh+KUqQ0Wc94jhxx35Lcsdh1bQwGt/E0wtCGtq
2PIYUyYWmRVhfdeS2ETsjrYl0XMgKbGqTE+wDZqtPuq564JkydwdX4B10kRzAgbA
OxHhHWR74ASYRFWQTYjXWU2wTpwNgrZ19mzrX5Obu12E4SIoBS9sprHpnBOjDRos
0NCFduomPgPCFbptYtfzIKJ2X+K9MvUZGLXhpFo2XZqwIEPGEE0PgrdVbteIWRPB
7EldbhVytYvwUnB1OQovfZZeP2weFzb/vb4ATGB24o2Wi8UfaXS1pGNhKqgNtsqD
izLvdN8isId/gA6L1fWxWs2UOSJcuKWGohiMhoNDnV2GAV4/I98aQJXGRIO47jGp
mGY7kzstwwZQiC964UWvK4Lcy71Ei+SGymavQeZGSlaQh5l1EF+IBnr16abAsMe/
nGaxhZP1dr/O5oVgzvSuXqJDLa9tYpXdkBlGzrz+NAqd0pLwd4Wq/4Bmo+mq1RJW
tbEEECEq3zskaYT1vgEFFlXB9xrxmnONs3qP+B/NqtK86f+Qyd5LomtqeW+OsQWL
d2NcXtAdWyb9RUzwOHh78R0NBp3AQhZQ+SKBRJ+YyuMgggDkeEU1gpVk3CuJ0q+2
a+TlGWknWzpsIxbov3JaNEjicqUsy9a2RKGIer+leq4eXaoc764molv934OmwAEh
YIMK7zCOEF+mWc6ED0iJn06iWF4Pcuer1USWo1+CKfC2s7FNAFui2rbgUKN36RF6
VpzPi+VDByfj2HcRvPZw9XzdWHGuEN89YcPdvUcCF5cGyjWh9t9XxuFVM5kxfnvN
FP+jyWXeAf3mnzbFVpKgO+R+xMDGt6UGzmJkggUc/vS4YLoqDtANyeckVJP0Ppl1
wHgFFsZjWBjsKWTNgHtnptA0kkFl7Zyt1DP2happxXi/QvQ8C4ewYuiX4RG2z7gW
i9E7E3w6QWOwxn4PokIsIj/ljOgDhlVQmreEaTkt/A5nsxMR0UunsarOocS16el+
Fq4IUjqEXnGsRlh8ljp4ied2Q1EXbXftWAq3f7ONmIIu+A8X5ZUliCmuw/ThKrVn
Wwgc3VsIbP5ynWhItoBBYhTDltuHimQTahC4EIqTlWJV334YQ3N+K5t/pLhcMNoO
XMs/bWTR6zQ4I/dUpqe4AwT5rt4kY2mGdp1/5qXIeluAyTwpqB1eEPuV3PXsmXPa
6C91/SFG6rDQ3+ATj7vkqD/PQebpCiRq0vTWcdAeTbLSfn/I78U/gobQ8f57XHyr
HeFu/HbJOWm61hyfMbhmhf8ABREfueW7SJy0jTLU4jDIGULvrNmMkGLmgwA0NIxa
vmnuqgh2oUPb5OHQKa8sBNhgOkcR+gkzvRds8X4AeCWNGi/Wb8FR92X66XcH7XeS
bWm9DSGmqCZodU5W+tyqT168rv7ZzWjkh52/hLEjOo9hy8nKMKseQHD5kAdXQzZ5
E6PEq90usLFPW0dmHZFHtob2UKuWDCvbjU8XAiC2K3VWvXUgUirv/Df6ITF6/zO+
lWfsI/CoPOVoxX6as1N/o633GCrOItxGiUhaSlGLyFdu3owioYDcgaCAMq7UHx5o
OiFfouDShfImtiCibVPYyK30ow8rG2xH7ODBVy1jG6LTU51zcIjxWrOZ/vFT3pzx
ClM0ltntLHmQc/Gv+3hkqJHlKfLnk+AZ4RnVAAzbgHuugThRk7Rb+zesqiCxnUCB
IsQNadgxfI2MGEPH1qD3+xKufUuoxQQTxPHUv9S9+JI+fIDvE1nGVjQ7FO0lM/xS
4kKhwwyQKZ06IlRJLMHnuoqxXGLj8TYG8nn9915eeUWabvxwe+N6jrD2G2UMaI7X
e0KpEpbHoTQnYRbFzR4FAH++cVj2OpP2gLLyxULevqkZILrxsnWDePANNGB01RQ1
xmgWR8B23mxc3wOu7VqUHRg9zVOtOdMppuBukAEJ2Bvx+Ox9Dw+EO9xlW2J7AOpx
Gu9xVZKaUost2mQ5an8xDqVW5Sk9S6GHXQ7MR7+I+sv08q/qXAxw2HhAStN4ioWD
yfgm+IK9j7PJVXqJv5dUiJg9FDsJ33re4oy35fN7hBgUgJ3QFBxb0qpQt3K0D6Ei
oXIqjI/+5q46BA8md39UKT9Bwb4d7YsWAq4EEzxuqmkvQ5tUBKvxoid/Uch8nPja
qzRFg4lcgo7PGYM/5kAkHTJ8Ar6LuPaCDN5PJ++4l2dY/Hrp9NiawFvxkjSrIP1u
84FQXD+ZO3WWZQQU+2uD2qRb+BP/P2NJNvYDgKLED75UHkrvueFOKkqqGqap/RL+
8eIhobFHEfh4gIx9/8x7fnQRl6XD6g+BhnKmRfpOGQ0aSHlopNgHmnDZY50FzI2w
wh1uxWr3/gD/Ce3iID+GKLLNx+62r8AJUdvSf6eCP7NJNxG6NIVi+ubwElMP7qww
1CjdoRiJyyitDuMmFOvOvP0mR+SDqo7+UL81ZPgfq23rIYY8YZSykUBJwMRqFd6m
vxVK63EchF4aW15xd+Fseu1blnYGJ9cObN9Zxxpiyh9ZZAtcpOzQp0AVqggh3WKo
y4lZGJbsnG641mCaW1wFiADWZUrEt7rkMPRNHENrRRDh8kCOh9WGH3y1YU+eNT+H
KABDyPU+NwJDZ34t83e2nSat8GDIszu/cCpwItXVkLLAz/AkHD+zrRnoQ5+fJaVc
AhVTndXz1+/cOyvN1QgayWOul5HdPf2svtOJxLfK/Sm8OVEGaMe+EbbC2lQTreDf
2tmIu2oN3gpV6wFrmKQqXyeLYghdIUzD5ssTPGFtmAm0dj3tB2/ODscZaF0SeyIy
nSbt8vE37N6q1nxGhW/mcjTDREbPgUkCFy7Nc2fKYYN8PB0C4D7kKzCQQjsSskIs
ZSHDyiFgDQSBfAMqYeBUADM8wU2MAHj6SdwmUy4mNFswAOudbDZitGRXiL0gUyfP
6TzEIWkJve3VEAbGVGvIrURcOi2Bqy8WUaNkB7bv4HE8rJY+CVORTZutU2VkwV59
UduKkFBsnutb8WaIpA6iQhMseXTMJ+w6qUD8dYt0Y6mpA/AaVBj7MyGyk6HKbQBP
N4cOT48Qj3Ua27h3Dsu81qpTfIhFJedHZFp/ZlMAzZWiXk+i+dY5oRHqVfpW4/kv
mQpsy66YVMlzCIZT0/vjY7m0Ap1i0DnAkduoCjmuNq4VwPfxYbBD3ciW0+7sL0SF
xdfX/UuHdT6g2Xt/c6ah8VrCVMq1lRnN0ttmKIYttOMuy0tzLW8jknu9/5X3H3Nh
HXk/391oml+CfoBAjEMKTRXjDYZfV9cw0/8rdqOKIQPMJuwzyLyUsFhSicm1g/rE
k8UuLTVMd14ItIhpEHuAxqqoXeRPqfz6MuMuIXzP2VREZLdlX3cIEj8HZbhkR42B
mE3mVkCoWlQimktNXVaB83pFrNaUE2S1Ou3/IQQ/ZStIc1Rk6EPGOrAo0z0uBtim
qxYvciQpoGYSbGjhc2EaCR3d7HPoHgDUHcm/Ln9B464WTw4MxVYcGFrmn8xlu1y3
f7fJg0nfL5CBt8Ybc6xKL1ve6fD3FV3wubgwH4OqtkZAtR5A6+3BrMTYO3y6RdUO
4tyM+/v7g0KSHdoh5iDxgzzhbl7rmIXAgWsY9Li5TFe7UfqI9Fz9+kFwh5aiBxhz
PdeMFpuquOb6BQp6D+j0J6gqNDXEksARtO+AojV4F/4xWa+iSV5deJo0vUbai/Sd
KLwg0abt7nxVk7YrE8r2Y6jTT7cPUdf1+HqCLfTkB114zO6vUwTrouxbDQ+qIc5J
CLX17MSvZVNc+0UnW+/rI0zGB3/3IDilOFkzWFlMekIEoS2dUejZRN/R0JMBR9gN
ey7GsPlHEUo1cwaoKogep8zcOKwtkka5yaC/7YGUgf/1cBoEnyjSSJYb6LjzVHWu
8j9mwVz96B6vUS2zuwIwjpFqtX+10+U/HoNwdxO3mC8j1XkTuaCZDZV7sfdLDcjL
S1oKdV0g3JHGQzZAQL4Flfr2Ro0/WB00wDlEit8LHlD5vNgpdZT+v3ndVOu2+Z+E
XGavv3O2kYZas4nftD7Kfw5EcQ+I4UhZmluVQpudfC1l8jr9+scG+Cvf5gMGtaFk
3OU8sGuj7ask51zt4Jr5O5qcSsAW4hBfGQ+DD/XpZjYUxjgDTE7ICEV+K1eZUNoN
6khBDJTkFhgcngwfuCclxJQRM4QBWZUeCOe3hD5dkRGDa6xqT/mStBaqlzR5wdGD
egE3ln1GXTCU0HYJ/Xm5JAqnHzRaiwDS3WyCbMUm7L+zETv6XehMtQZY2sOnJ6JT
e2/RIuDUSsKuFMYVE2hPlf72gAeCAqUPrYH5Yo5zzL98dAOwOApcBvxznHi7qTjw
gUwjfCnakM7WRLdG38mQDva+cruk5zbk1x5D3fnzibXTOaK4X9tLqcnXyFQEYH7c
W6wOrFcZSFHlAn+PAWBqaU6wqWjMAwjIin396EEOK1kWCdsPTzqXi91LBNOF+7ap
dqsCAfG+OOT7Fy9kkxGHAOTVjUdymJS6RCDmeJPE+gqR7jKcCnE9H32sgZoHTZF7
XQreoGDbZsFYXBYJ2NewDr1dCtyDzFMyhRrFe576mCE+bAHJVCSJQ8pxRbx8QNrL
l/2z0CIu9adr/GB7+A9XgoPMrqvcV/aixRIAZulK4pFDp8cZad03Vb0MF1R/OHli
wpOqUlrYC+B7qebe9DLxxg5UrznPt9Zotc+BTxJ7K604o4V3XEjYO1ySrBDoxtVC
magH5q/6R45t6znYtQ4Hf3AalEax9vP3Qte5cfFYDWh4OSutnbD4dmPA5Kwu6CCg
1IFaZXFQtAff6tl5QfKhVGCM+NwbhQryuMC1TjL7mhCtiwOXF0fBPmu5ntQc+qcn
q6Sdbl7+SO2BbG/+93qTCXhU6IqiE43GcNSmfbwUrG9qaFkiL8aIOe1j5W8U+8po
+9cvR7cP97RlouQ3GJYOVJV6/FCzg4AdqkZ/KdlCI14fHv8SU7uNbAJK1KGnx9NQ
R7Y+A+ORbML/oZ/M5HS9Zppv2FAT2XuEcVaWz/mDEWMJCcTuWd57CZeB2+M/lnga
3FGMhtxbyM8NlJjLpJb4jLcfe3m1Xl8/W5+7W9Hz0u+E53SCGymrKNZfC15Vuj5U
3hQmJjPJIO1gujEhUEkfFpveUXk5Lfjp7Kv04OJkbi7KwsatCAKtCOBswFVmL+or
O3yW/4Y1Rz6SrA01gGKjvg+lK2t04OwIaTjgiZKLYh7yp5QuurizzrdfEnkjjK35
9zz435ou+0AQ2rD8C8D9mEXjPdNphtOPFWtrZcATp97hS5C+tDOAcpC93jDWIhEL
ynSphlTFBNZIa9F1oTJF106nXn2OGplTXJWv3ySwDBzX7ejhFKxo7YHegmhUPvpX
7CVzjjSTXdYm6cXF/o9IFy5Y7jBJDqs5OeKBI0287IXyWCjDntqyzDN1+flh5oCB
5KBfrwGvLiAihYG2L2GNtxvDHsPG6M0+ILGl9GuScGOgM/COtNjk6ziuLo7ViLLo
RrElCKBabbJjRHbL68ymBrI1UeRf2P7tg7DG+SrG9Md6StaJnh+jyJPDoo0ysbgj
kMOyAaCZk7RL/uKafUpk+4KzioaQZ+H489JG2IWT+9+QLLmI1vT35oxAurmBB6DK
eUn5AfqbpEpKYpaLVWFwevU2fqDJW6QoK5xmaifxwtyEJpX2tpcYV80bD6SSpb5Q
5//3ftGdFZCkDPdsnQkMZKh7ssHosal1pzAiHZv9+6FFUK/0AoIG3W5q+47wTMlJ
LTBoECCPH9qjSm7jo1FqEUj1sDIVY0pt4DA1SZ/ENvg/JxsZt0+3WtQyERff9thg
pPCexBbI1YuoXQaJ3if6lXeE5MFdJ84FK+sSEq8zXv73ylP2FrI9wdYoN06nvA61
ZnHt4CCYmJzevKpFLfCALshgw1FRup5HqSHnuYBg7Fw7Ne/rz4MYBgNL0+0w02IU
QBCOQdt8A3OBCX+mn4jtV/nAGZhn+J6NCXVFGXG1sXTYb2MoHPtRrrZmJ5hFku/7
zjaI1dZgUe3X3WyONiF68OP4eKNF2x+9CLvsQCMpDhzk0ZmrS/XKJ742pCQtSJkr
nd6fj8WgdIifRzv3WlehDNz/9DRduTPniKTKKdNEBXmKK23SMsgHx+bR0bI2zNX/
0Yzynulw1AHTAuY3hvQA8yHruvFSCmpeGeNgGrXecTqVjIql4XryU1WhQwjBGw6K
OFD5FkE931GIRND01O9wJO2LNKvrAPPBQJPsdIrUaX6Rll61wZALGaRH9wYQYCk4
WzmJDEOd/HdvNLKDfTnNV+nbN1rpDil06CcwIqWSCjilA1gIDSdaEXqaYAB01wCI
a1hMGkUVJgEScO6PL+PnGznYQmoGg6GX9URYO52JUr9VeMigEzgamSbfpFW4mwTF
qY/YRv2SKPlO2YumbJP6ji5Qd5MmLp6A/tpgeWwkyQNfbCJt11dbOzB+0X4plzrk
loSKa8MXT7AywNZfKGKrOH0qQCMyiDrsZJGPmPzhfgTaLrrcf9OmYggt5I46GbLE
W3L7/WQlVRbyQrhE7anfPbeieC3Q0uhVEIrPeuh5WmHtBdW7dqWERxDgb+FxTzLm
Nu+5xtFrSDhA0b7BA6HrDbwpPxPnwc0rgnnOqwNG5PY8R1jHu3JgWekTU+2FguX3
DbinAczI0F+mbA0dxdoo8GZNt1mXWhzz+8A7vX/12qfFHpnjuLp+wXXeiwza9+C4
cz0HTT/wuGAdZafs1yeIvfw4HAlUT0RS1UAAd05eoVnDrjGgUZmg8vkmwlxunsoe
ox8dkCSTAZzKRrgE3TH8Uq5VrHNEcHa7xHew42bddaDd36V5MGEtUUbFVAUGob2w
E1saJuNoXKXpsnb7u/jZqrzCvG8iduN3feSQS68VvHtcioKF01pSFTPK2FRZ0Cu3
gMh11GLb6IqzhCQnt7amXS6/5QladpAzd4x2FdzCF3GTBYLchsKw681ggXtcb2Rr
FQWRRpYcNCoQguYLLX0f321K8CQd+OuAGAZVnANAzmjJrO73wN6+6xJy86x3JAvk
Za6EL0nR0pbc2/JJjFVwTiwwheT6jxDUal6NfOFo2MX+ESj6SQAztBKbDYcnucvo
g6n3m2NUeMr5Nvbur8N2YeyGRB/E79Uu6xZ0BjhYCS7oV1mj/cH88ALgW69OCXk5
pWKf54Hj0PbOdA/FjTJi82VFcBt2c2dJNihFzvoVhjSoq7vgy7GZOZJGD13MPgIR
GtJ6q9rmKN/q/4A2MCBvuhAOnZ4cIUYCCqw3oFO9t8HskokVViQdrBpopFwUjvRp
fGYwY8SvHT0cyAdANYWIc7yRwjiJby6+yOpsTuHIryPbSkB3zV/ywoBfXU8qT4rw
+kcfC0luUAehV805g6cIbP0kTi6TsJpiXzupg3XhdenDSr8Zjpoguwwos00TLPLl
xpUErrL46XzMVhTsbD1KXj6oz95yngJfMB0/NZbkzXQEZ+B+GvuSk7IYUkpwflzQ
F0x/8+9gi6555jEqLvj3VFu4GbxLYOVbCpGFALyin16PV3YbiNyERY0jh20EUZAC
a+z+j04ekih8XWcEFryUhYcJmVPanP4AcYcNwGIWAKIXRmeDrNB0XAWvnt3g1Qj8
/0Ae6kmmYss+EPCriEWe6qR1EExouBSXfI8wFINSSMFi9q/fiFepY4eubHYFJ8Pu
lEvSAEo8KvS8a9zBbMv6Q6cjeLdLhpzCWbzegPMlO4elk+I98QNDzzsiqVQflOZk
nX35iD/yUj191GR2WAMODssD/vOF1yHt8DvXDClgdWJYFrJl5j60ZPWLYbI0rxeZ
Dq0nhLNhNNVBUW5NDEulw7B7gLmtKPSktXOE3BfkTr89UnItH2qfAjQ18DRHhO1k
ThZAmMxqlVGt+Cq/0QFUwtLzr/lKJtt2ylTZ2/1YlV8tZgH3TOA48lwhD8c/8TXa
AB/R2x5rFlcDZlrzQyS0DmyOph+FWFAQCmr/NWn4h5XurNihrYJ+UdHMUTISDDgD
x9OkUwIVIRwP6D8ULUBCFiG9F2izEMBHOqPMB/Cr4CiUVSCVDc7w5gW+bsOqr0la
YBm7q43Rl83yOkOw0jepkLVvvr+knCqc1O5KKe/BhhHzliZsuxCp0CMoluIxguZt
wrMd5Mvqol+qwnPBGHBqsbyCMLxlqomv3huWjfvEgdpyHq6Wa6LNltQVOjMAFYXU
D05EBszuviwHRyP4Azd/KA7YuOik/T5yCvuHm/GIh/mA+/N6Kg7SXTd+5ge/2N1A
ZgAPkdRrnL19nuDz0KhHz/n9w/zDnpjsJ9N+Nzf5yKinzb6GIqwUfBapO8hj5P7M
o4Ony/oVTzzCv7RPycA3NZytkcrpmtxrcFCuiKtjfYk41ei3HcORhvwzB0Mb7Kf9
tNV+VhflQbVZeiMtSUBS1bqISckQDd3YOSwmyb21GdTWUPFehyX4CtTxmFsuU53z
+6fpWtaQH6AmO4wdFbckdxGgARnPGO3s8u61HwBMtTev3eMcJoSI1NhdpGUsYT7L
xOt0Ufx++Tz0sq/9cffoal/S9c9NspNG0I6ST0YnT8MzwlFePcV4JIkB3ttQpYmM
zUoqa8ZXq785gcZ65flmGprchxAaf61KIIinYw+LB612qXC3iLYYvJ5bPVCk1PRL
pjBYTAVJgty5uYQ3U2Kn4PqqxvnUByAT2wG3WDGNnGNz46VqYu53PBmOSOL2ogS+
ZdPCAHvbUwYQ+jXlGxK9AbriyUbcuhfImaYGvYJWPyKzELhGXpgXCAsH0FcPfPJQ
spILd1bn5F8ajIz3B1bDVfSD8evn+v63d+OQvT2/uownvZz9oSTXRK/wre4c6pIn
uvfvQJfwu9QEGL8KtRvv7GzJp4lWvZByesPSoaml3JLz2SvF9er137k7qHTRZY6G
/TvGPkRzXONbkZ4klGGgRhu6n2LeJG47jy7nmfFBspNtCZ0O/VCQYlXQrdAaGUlP
WMOyGkw1calR7eYYy8Hmf8++61Eb9mdqQmkW1FmP+vyRqE/JpivlfELxpjDlZPfi
2+LIsQ4vb6vmcE9anDnJbwzbM8VRsdX4TD9+vSb9C0ZqclSQ17lrMB6SdQHJsEmi
d5ixuyLVdaLVPQ3Wrd/wtuWWBytVamN0nwutHY81B/6cPoxQR3k80jFT3qclMBsG
Mz1+BHvp+BvGtuEayILcg/f8Yq0z6Bb2ws46FPniNmIdRPHhK1hFt/gS6d041EVE
3f5p3TUSCVqUAWnmKeIY3S5N++B6zijVJy7S4rRkjw4Nh9g1iizfhRxiM0HTKxdE
CvYPMDR8Vw8wazia0mFqP/OHm+kLERkJzjoBN4cT5V9WzobOVUElnlGJKmaN6s94
hDwoy5AN60L+MjqyaGTRqlzcoqcXcU3F8yMn4okwDDCH4VMWKMjSqBeq/PuQtUKe
B8qFpUIpKOj3GjFrRYQeZBWJgrD8Ao9jbhU+/zPygJ9xFQT+Eds4bMlXiz9wCmjP
pTvjQbr3NbWjtDA8yyo3x0aPc2oaGqUQRPb30fQfpgzEcqLGW9MYfF1pH3YIxy/A
NvIpiZR1HBQLB4oOfwqNBqEe8Ld20Unnu4uot230WnIf8bIsniLR72hTAi3c/kEg
a4Kn1c3RnG084LtlEapfWaIryu/XAJnRcPrq+K1Iw/o8VNWEu0iH4279HcWsIM2f
2X9+4iNaelwd5BXU5VSY93pMSiNqcEJJwC7hwIKDahxTEXQ5edDJcz6JR9FzoKeo
gSohsW6r9mVMM+md3VNzwGKQadjFiBN3H9WQcxu31hrW/sQlUy4d8gNnqg4+weZT
dV49T7uVyL9xz2dK8JhJHOhB7uWXsyTnH1GrELTtRQ/FhVbX0E/e/2puI7oiU0Ag
nK37fSUbY0g890djppIP8pGOizYwg45MOWhBkXKlWJpJq2nAncC7/ZaYDyoDwyGV
YhR19CvEUNcJXjuB1SmLBK8nnRII/FdAb+RdcEaEFl0iQ9Qgws2LMfEKD8WaqN76
EE4LFdHoyQ5neB6gfsMT0UqOYnADuihpFuzL/xSRcQHf/KbZ1jtPo2pYn8b86GCN
k7gDo+klx9FIsBwKT9+pQxwQdJL66MO42Jm3Uzsl7VBY5Zr7ayKKzIw7ljrsNo6W
zsat1k5p0aXdIBw1Wx4m9PFwHScN1zvr18ovvD7UqeLJNm7URCZ3VuIYOrl6cysu
CSDQ3KQbAO5EiNy0xK7mWxcbvbsKpwv+qtyB17CbyBbCMqglSkIAKGT2TUun/cCh
VoDmi7tPOaZBEZl6Afgm6KrZbSOflPIholoUagczz0TJb6xFqbt+ZSJpohl+njRk
fdhGaPtP2pdvMBqpd0lhGU6EklJ9Y4O2xmmknbixSQzJcF0P6KoxRBGzkE1moHiQ
pgc/OPMWU4cCtLYoIOtKhc8MxxqXG5STgL9ORvFrzBgUQTn/1vmQoWp+Ja+Lp3CR
MyDnLQFbxIT39QWCl2tI8jZ9lqK/eohLtYMQ8FAH5DWF7/aWwAwSpcFbJZ08A3Rf
XJ1zticraMgUMDI+f67f8EJcSNvvHWv6qSdGMWNW0JeQRIHsFpo0R+060TuHWmPk
UMP3sEQtIct43/7mqJxI06aF0St4lqrHKK80wz5WZ4FzOklyYJvnAB6UHMMlMdUI
qDF3epm01Pv31GQV38tpe5Vbt35np1g6Do2qx6G4Aguf//hcOtwmp0uhMLUoM0kS
uMNXk60QRoGiihl34Y9Fpxc57Uae+9VpM+BjNDsFqRyiM0S4YFgiQIyaf/ZU7/tK
CeOfXx5ZUm3Mcs2zGfgrrX7VAW7sVX5Mhw11sY/9EcmrNvVK7MGREVaLoHNWItwu
wxZJWLQRy3z09wGuSmB+65mTacnevsMh+n977OkuCgxu9ybW9HiZy7krex29l6Fl
PA59Lbg/ZmvE9fkTxN+rkwpDJ8vCV29FM7+Y4FGBQCJEe7pbQ8fn6UDSOXehlNdF
G3FADpx0g4ND6Fuo9k9mhrlaXOC0U3cpKR/zC3w25SKjH8a+H1IRNkUvyaU3ogHG
7lUfztuHzEQfIJax4p2hDCamhKflzHxYRCiBj4GIxjhlnOhnMjlSbwKeuxHf37qD
/3h2Mh/ZtwKpznJMhY1auNUyBX973ZJOJnfwbXRm4ASp/Aphz7oMuWV3ce/EA3xI
G6GMjcnsqZYBslBarxRDs3fMGjs2lQ0EGzY7UEzg9f8nq8Q79h02Bbn6++wFZSaj
HFaPVvHTghprQBhFIH6PxNvz9nTc9boF+K0BCprKODGiyrfbUc+PjRwHe5+SUXU2
MDU9HZ7VnDNO5HPqKgTF41DmFkgC3N8VxX7SBetrErwtWaJCy5LUHQxwFdLkCGSX
TC4OceItQpNP0gfuPhnbJrVFqFu6iyDu1jOlo0w7jl/L7VPUB0doElIdVQFRwwOW
z92IWsJoFu2ilCOrePR+OxDAquE/vaG9BWg9uGa7JM71yE/c/ii5kmH5SmJvUYkE
c2ZqS8wz5GGRM4Z6X/v1iKKV2hTv56v28M8eFAQzREf8WY8/R7oFIlBuir2gZ/s8
fFfX4M7hplMYTN3CPIRBo5nQZMqal3dx1vgRPQgLkqSFry0+OA/2T4RKSnObYFnV
pDLhxzjgC1JSF0oPx8gZmMl88qu/I4wnRUYmX4Q8tcborfIwUUI3B+Ea5RnkK5vl
QLQiOt3GY09h5h+72zp+r2ZAatU16zzvKW+UGSW5ShTmrwpt+G0b9rfMicy4i+eV
GaomxvAQ4usGMxANLP86tYjBOteVpMX2Y/Ee669z180vio8oory8Athdtwd6CQCv
SBW2uF4zMC4T//EPYYjlwmEd+i8aIFeDtVNJGBW20g8tRmnotKeb63UW80xgmi8l
pj2uN0pItkEZ0lX6JoNHfHseMNL0NRKG8vkVANq1P1P9pFF3rSGL8NrOI4DfXAO3
3LREOjgyiukr7WsvQe2ceZFxBCn6DVmTyjD1Iq9H17KEuJsLol8e2P8calXXwPu3
08EXOZexH0wwAouGKy+2oLRCUHF+QJx+77giFRKfrina1+Lbre5xcKZxqgeMNo9o
jNC8WeEpxX26jVZqbc2JUTJw8adn4K21dGexcT3pnU/CxgxFOo6CbliN9+InAWji
3Unce00RArVW6Hiq34LG4l5sxsNPdSwtqMPZ1JGhshcCyIhhiCBTFN84etpKxhvq
DatRVS4Oj3T/C2oqf5o3wI5cgIpLv14KajaJcOk9egMXFFVrJ8i7m3/nxPpHxDro
qlkedzW8ZPa7gfBRYdLlhQG9cMHVzyF49y146d6ZuvBSKsnTYr4+s8w77jLMmlnW
hiu39JEQmrWDe0sdpyyeJR8+kkCe4MzhYwdHCHqPNALN7MffudX5Q58p62L+pHwJ
3jVTRsG1ArWDLuFVhd1vFJffrY2AZ1j2VKZ2dV94RSLPRduy6wRTGoOhJrQ24No+
xXwwuFywhoVLC6EHIuoZNd8MHjp0b7wwyOi0dtbdVqYjK8ZuZAgZ/7xUNLOY8+1n
fJlsBJlHkLNtTGYPMZIWbcIXemureo62ZnrSZakDdISQJQIYQXYBix5huWKsTaSC
uHIVXlyOXS8oUmBnzonZTMFZpefOPmFLTp1LxiVt9jmFPl/TgbkbkRVJuUz0iABG
Je4AEr3MgbARsERBT5w88htCToQjod1QSeWxFwvRaUQso8FSV3dScdswY+KEdhgC
5lhUiy97MQb7ivQLC0hrhHPvRF6kuQ4kE1hDruuBXelLDBjP6CzrzIFslGBi6htC
JwU2ghRIE252AT+dJY0g4uQHlmeefZ1++v/QeVPGcZJf5hhLuHb0jCzj+xuOBhi+
t0o6Js4ND4MToLb+DyIB2EdBHlXnzNBjSG1WMRHTfNxJ/hNNW401YWwoaAsQcqgf
cl5G/s/hG5zrbip6GctQR1oSz0b3x3MaltD9nxI8PXsMBcN3FMmFEt5ewGOZT24I
Rsj9zvm1Bgjed5LJWWu3xW49Exh5G3uiKhU4WpheUguu2I+NnNfCUg+WrhrxJv5H
mm3qCfvcqZgi8CD12cwBdrO124z59/S6j5r5UzVyrehPP5XJzDPvRiFDQ1eQ5fGI
ylgB++lCxi38W8fEUjF2oY+N2Kbxzt1xL0U4L0/JBTMHtw3Ni1gY4IaoM8CEFsEL
/yjJm+6HrItguczv0OpgADPOE2iNXo2HtIHXeWv40NzyUc08ukW7wFtWZ0B/fN9W
g6ueOXuO9A58574661KPnwusTUOaUqWueBbGx0WEzq3mEQZP07HxviID6IfiLtmi
oBgQD8jXwJkoLC9WBFg5vywa3tp47hXNQajcaP53nMOknwJwYMiLR4bkJuzIkhVK
szQB0BuPoOzB9I9quLsAjBhmryIe+tXXT2z7GVEBYY92Bmdc1ntiLGfzFrKXqB0U
jQ17sZojmSERIY/StzvYQwllkDdDwS1mS2nz21GHRBjswOz7A9RMF2sOl/H3s9yI
0fASfTg4NSBBOZhKEJA7a/97jqeGVinpERvom6BywGmuAxkUEFl5ZqQcgPpCFcrN
l9uEljZ8hHk/DysQTaGIc4g/A48PkRsly2xdUu8BUr0FJuinep+tVKejUxEkWDAn
cizzxJcdgXv3vap4ron6tQbHbt9kknjZh7QUkVQJNiwAoPYxTDvNz59t9ouQKoMq
pcfnDw084G1soURYmPIEWOiHB5iZxZ/PRCqmqH6o1Fsdh2CHjC5WD9oMlcVUWHw7
l2O7L46SKWFioJ6hD8YC+W9t1YGeEOPROq0DN5TuAriJNX8LWTWtN1rJHijApkl0
4FDrLhIF3BoIlv9NU+3xTAQTuoSujn9cMg2ZYcI3sr0Ekig5sRU0tQSo6D/RLW0p
hv79BO9pceOWw3tjXtfXNA3rwSX2va7YIVkAEj/nDrBgTAcjAKbbjpoB0QZP2hhg
Xm5MkIJOWwh10xfVlaJJMav1VkCAN07mDHofbcHyHHlMagHwKnUpS2a6FeMWDKs5
h2j2QFU2PO3Ja+TY25UC7P8vg/zqi5FTPBZZQTTHD0TPoOPBnvXn9BLmmrg8JRfq
j4RbbZ7gB8qX6TkQ4fOBxuZHriYNXfRdsElQBxSbwClNxBk91FvCP/iVIUAdeTRW
4XEFPVgmuEc2ETT4uvBPXJd7FwWTsPCVGLOtCVcF0pN2HzkDX0CmLNtl3i+preJS
7z+WBEoVqASneaJrgPOUXmevmlSoQzdPG81s4NVoKMrpIGc8ULgS9+5WzMFfsWvp
M+KtneZyPxnZXegKHkyPNVN9skuf60x8Q3RARaKDy3TQ+M6xnk8AguzZwtP++N+u
6vSAGNjrcuDBG/LxHNHDPlxd2JUkS3iP96qbN7ZFbr14dJGl/dVuDn9Mfy933Ela
0CpiQPGEgHj2Zd6UNKWK1q8TJDQYckG4/mgSn4C4R+xXKOD7E3ZuRZhAZm5mo6g7
WedRFyr9oW8wwrjInV0jxjlxz4HqMlV8gjs8pSt+jy+dHOX14o8polRenbVD+CAI
00MPDIxieRL0/BBU5UA4rSennFI7TVYd1YqECj9AxH4v6Pc30vkJtVo9EAlxGwzP
nQ5+KKidz8jLP+vXUCLLZlV64Pai2nuqEyf82t5apHvT6AqN7bo8MUFKMdeSmeJU
EJlg5AKaLibTi6/GMNRkIOinlMSDZYoBuPP0vnVFOgbFNPqFTn2lXijZRWhojBSs
QXg9vTEwovoUi79KxJUXAu62oEgZU0dPeweH4j/+z+dnv2E4fyOxOrnFzycDXtSF
ktgimSZA7syR6J1WJut2uBtcZMtqH9zUzdpwIN0NT1uF6hgl/l+lRYNGVU7xkJx2
UfuBvMG+KyRPgaVV7eHPcI8F0Dxs+ktQaS/QGzGVa3WJ86yBV0Ly1UyEICSV8jPL
1dVbn/3bzfq4fp2R8TnIwPzIJt1JAM2047YM7t1Pz6w5oKEgKTvGkfvItQyslZMz
RnAyfEJjxtSDpMESM06eXrrjXVhh9BX4O3JRq7Ckeh1tV+FjJqi7eYa3fm/hQYXj
k2DKMj01MwX5dK3u5xXqCKp+ZPvWSzdQ87mdSpRdcJaOliTJam5E/ymXtAp1xK0y
xwMbNph7mVvIbGyPHvwyARISgAkh5Y22xbRqRRg7xY/L8UZ8hgTipRrI8HFm8Cna
ArE87OP/mXdRlDh4BZVDsaA7Mrju8OsZGv0rbSmz6puaSg/AXE99hk10R+xPs12T
TWjV9valcAMH8eablEdf+vIj+aLmdSaumLls9QEh9cTs7CJcMjfDrGWd3SpCZ2EN
C4U2MdYMndMzfg9bWuxmRTqPwrpvu1lpyhgPZZJ7WpI4D9v4xM+ZDlX50lJYPWjN
uw9HQolJSUUHaGY/xyRiRekEvjI26VNymIdQsRc1fH4BYDP4GgsI03e+beXlEt0l
NAnJlWgt/RqZLWmAyoVBStodlMkr6Aepz0vFrqZM95rj/ba7uzSV1PNuYYap5i6D
IytaQCQMilttgKvpBpiEiHkKO2LC2qkZeXfcsBQSrsn0kAQ+wRIHDoGYejVQ0iCj
Wy7VEazFt0CZR4QbVOFgqfkJWZfTnFtRgmJn0W4wgPkSK33XmoQVroGXhkqp35Sc
D9ysmF1gHYrb6u5DqzOc26TRYz+JZd3S5dv6VDHf08bJxa00jUYs5NBv9YI1xsmV
AarnxG6Bo+I5aEi1xgtzWydrDhxsbreLXLQkTOMmbsW2UbjJy1/zw2EmCqUKGWjv
Al7KzMqGS+IQJ8uPkiixGqs0SKhdoQn/bOJRbA36LCUrcJ6Az/q8YZM+hcBVWikh
mIkfe9CP2erGa8BhlWMYkypu6jlD8fA5ehqmu5/JLNqF2OKbu8Wpjj2z7dVJq9Ob
QG6ZPczLz5hKUjas8OnelNa9wCip0JX+BXQC3YVVbS04QUDgi/4UWMj9TR+yZl9d
Xb58pZcxMTFwWhbRBxd5hG2CElouc1R0qDWUltnONlzqu+hyuNJJXrc6x2qiuV5u
9jyOPxFzteZbFW3MF3Z3P9U3+ZGQLKSD7jxOR7a0P4NsOCpq4vkZV8/3vVzs/vRu
JTFUOa+pAb2Ui9yFzB2dNKd4odIql3pt23btdZpJ11Y0CMKcARB7EJw77J5a6ApB
K5v20tbi0QG0scAF5qaYYkuv210q7CYchRV2Lgt6fRU4KBX/4GBdsrlkU97uRgFx
BqkUq7OABe+QFcc1bxw5M2PeSs4br7lJAnxnlKAOWha3+MsbR/hI4dr+OQKxbBPA
P9PvyfY8+Ddirru5QEdFQKELdJJx4T6v0YUwKzbwbpAMEVrxNT5CljmTS8PGj8GC
FHwDuH9x9C5Z2BPfKw4ss911cfzOhtd2XfYBpSMP/IiwqFT0L9i8boDhvzT1uY7j
v7v4h6Ft25D4YrDz+ftfFeVUcnHQDRBjjXNxcBMFo+AflrFuURoaLLuK0hvPjxLY
qTLhTqRVpEU1RoG68S95mXZM/ioStZ37xXspZpcFMnQ/P8r3+uGiE8EkoOc4pQEO
yHJn7EKa3IFr2rpN1Etq3pq8gOViRvSF5ZeuOdu+IwuVrwYp4Df38yvhNStayoK/
j+RRlsk2cJJTQ3axYYx+pmGprRK+i04W/acbsCxJ7bPLFaNoPzUYXHFQ8qHxnuoQ
KD9n28E7cG7QbUMhSXcEdW6HgnbHG82kJg6NSJe5ubHaRdUlsN+IwIvXs9I/QYD1
vXC6JUxBVe149phn6Xyr0H7ZuCRj2PFfgRTjm5meZq8/Vo+sMFnv6EKUWfs8HrgH
i27br1zkQ4HEcGSfZatpPyVgaChx7v8dmeYVKuw1O3OzIHGgYAgFSjCWMegVtChA
o7T0NI3reAdPstUgqjWPCe+GjAKtFcTnasRbLXvKDCI1VTdCSAa2oNdVpsyqlN9E
5wL3kTlVR1xRQ5WWvDKeH5X3rTCzCgF7hAawWtuIIIBEH9uqlOXMaDOoURJAIDXX
1XTkYWWqIP7RKmCHWIbYHIYMXGsR74d2aksm5njM11ZKt0k1I/7f/LPHUSSJ5++X
6VbgzdDXBLr5F07jtEB52hpnYkQzWr7ySKSoj+9FzpAgQXAZeYDAXHGLaQhBHIwa
+5ldz+L8M/g8DbIY89YRzrpRu5BHwSwJ+OEOMCPgciv38gd7UeMAs/jNbq1/JDUc
PcwNItxOWO1f1+faRawRLkRHsteo9U9mkRfKAtaQYFIggpI2FnccQtyQ1DwcCOq0
IVrGIB5BAjYazlbfOVUoM1qDRIrvj6/WcaQJkvKM7NLIRP654lET+u+klNW9rrYx
p55jj+Nr0d4e5VrBp+gMw+J5PLciWvd329G291++O0kuT2SMq2uidv0loA+IJ3wo
T6Dos9M4S8KJmOPQFZ6wVl/sA9ziVDPDQHqd7dPhSJwpVC9SWkILyQgQt41K2Xpg
nM6OB4kfiqPxoAInbsd2ZdEECDvDUhLWNwny2ro1CeDT9ppVCl8krSkgneiRWPWf
ApD/+5WD9l9As98+KvoCgInpN+/8kGtnAw1ddu8PW4wTybIhKwfKEIIBv1Ay6XeL
X96b6lZeZBhHuow1HD2uSUeqCBlv57aOx2Io1ALHGRHwRPvKbCokI5JHWWoEue+N
GtDJWppNHA56NK3nonbx0tuuzocOVRQEhSx63Cz4htdy1U5e3PZC4Ep680t1Hre3
ZC6DxkvVAiY7q5QmHjMsyMC1bGZbsSB+8rzMETUlLVFpAc8EF7l+RS/zpipCC5yE
xG30wUL6imFG9pQuz955dgxPh6fkwlifFvSjp93q7dAyF+5MlzKRljxlnxGYqIjp
hZ9C8LmPnpYhttm3oqptyQ4dY6FR11mrDfoIRkgH34Z0mGjQmAGdB78OXCdror6H
CHOkfRnYn5sk2gWE6rIKYuGUMADK4uuCdBILtywLlGTb0+YjVjiwo/t++tYLJKx6
E34CbnEjCUhOVTyz6vvrp36toCP2OrMbjYIX2KwdJJuyGe0W5TFmfGFuPzy7x5iZ
WXHKYhvbF0arMyILszg5j70+2rMZM4wmh3KKw29JZKwq1jfp3I9abSx8m6X4roZk
8OPADMnFvAwPlxBZFTD9tBPS5KreHWBZZKhISCVn2dJoRZlEcMRmcxFioSQrTnMj
sxIwzgX33eoDHxZM3wKWSCqemp9cTntPkYeRaoPTfWoCBG62GS9DRq9I6QgHVMMM
9oHt2Ug+Ypx0KRGZH5RFi/59tsyLlIVr+ZiQeabNBPU+0UovH9my8h0oQWDi6hSN
LDYKemMpqDXIry25SrXJ5f2Knt/3lmAdVAne3YxjyQgrjconNu4B1xbXRqhiei0y
jSXS7sBty5X2LVKlGIenQv/hcH5bIN09ezRO4AtYN0We32oWNwouaj0shvLaUMFT
b0mosqowrk9zJ+sVLLnvadyZKqTzA8HoX/D2ZK7os42zMkcXJGErGKwGfCnD5tQO
UOb/XWkWZBByC6Nqj2Ejz7K6n+GQupuhoYi2KA5WoMacbp8luG0ZhNrQey/Ctrwy
IF1EQ8pGRU1JGsY7pVdyanqo//Bzr7TcWE1fiD484/l29B2ugcES2e+jA4R5DDhf
D+h6F6QOxFZ3A/chc+8JqXKjR48UWJhluWt58/BsVIbqPv6U12Q+A9S3wGNsri67
NvMvgE+MQZq87wgeK6bTMKmBNPXq43h1jMCT9DcI76BSpAMCUek1ykLOhEbK+UEb
7RROaANHYyHTGo29AQAvZ4OESHdpnbSFNqu3dC3tyRCyHI9okyU8ThDREjTwqvzB
8zf5RQHdZSfAlC4sSlxryoC/VX3HtDkB5JdoNo3u6OlGMWIUgEKy7wNwb/txBV7q
LonFtXj65Sc2/ryrSBJIE80XzjNPIWhIfzeBwSWgzO6c+znoL+Edz6w/5JSxFEI9
0EgFFLjMWAM6x9LsxdzVjUW+U5YxTAs5P9NSqDPMsIdnFOY/L47Mhu8sMzAqrbB7
0HZkHzqncN9aa24bcaIWDLgaT05uX2pQrHIox7HH0WaB3qvWiHZqgM02z3gqy4KG
23FmG+4SF0ul09vs+l42p2Bg3HQrVs2nOpuhBgCjxSLAcseI5/9hQWjtsWILDgpv
3WK7ugq84F6Apd5GH0xppN4Nrd9jBmOiBm8SNQOB2Gmew1DzaCBM8SJJUsUMXXI4
+2huWGM7KJSZdEJGp3jPRs44C+xPStNpBM7lx3AfNwZciVxPbdh6kWLssiyf2yN5
VhprZ/aLV2ZLRU8Zuw1eVN7V9MTT9ZQ/ufmMyxyOmFIA2GO82BFTrrGxlphydh+B
Sw/Edi3THmjlLZbuSpg95biLKvLY8/A0uDnBxmPBPZZSJOc6laYj8ZKvGZd3vBN7
CJNPfyq4zh2pCRNRHCL7ceoAtn+9KZYwO87jNBLQ5BuJbFVC8TAfoYnXBD4T/A0Y
bjB0u/zYXsrRaf0yS94pxPJNtlznBmuRzMf/IA+OFTmVaNWnRNLLZFlkdKWhj8vY
WAx1fS5VJCBqdpyCgDefd43YJUlF/skinA3jP4WrpPlQ/U4g0kmCMs7CSVwNvpDC
22cLWe+tFt+fPsRrx11vL/Ggf2lwvgancZfagG8Na9KAIZPa+FJST0WnqMsd+PHt
MCrsG8FuOduQu5q7N8mDlXb+VzfhHW3lxV3WW2tFIbU0gZtlPmr5g6nL8I2cgLlG
6N6Z3ZAFAOH7cPAS/FFHfC+2XAEVsqEC3ho+Jvhtl6szQzXR+uUgdU5dE38CZ60L
nh1vXkP/hzNRQ++ie7tx+xrbu6DEnQJ/CH+6TTeVWmmz08qSTMeMBUEV8GljFJGe
ZA/JZjs1Nhwf9jafLHweKl5EUuTNDxl5Xh0ahC9nC26vDhPmkX4l1JA181xvxza9
kZqLhq1Pj/ANHehH9lWrJEaySpfwxTjiOCvVVUsjq+DkBKjJ/Pi4X+qL6wfDDBJI
QqZ7uVrwtZDoxcd2dwLNifeQ/TpvFySVvBuiUTrD/UY4j7dZtky3t3IGWSHlgmqD
EknXJPIxvI2z7vNLqxwHedg1SPkytBgKKUETgEgxYO+5pgmutpqIRQnSGkZAYDDv
vODlTzUA0NXD8IWc2ViI4mIcQmB9FEOBrj+7/U9q7Iw64PLtp2CTNsmRX+fcazhR
NVpvAr0GTVEU5niSypZ9QGzFGlkIB+ttM8LSoKteXOqgcEeGaGgIKFyIXiI6PGMR
UpCPDIzQWXJcAcu/Tv0tzYoAVILVV5h3xT7dDiA/mkeJMxsamHiZES/wIYLcZihy
7rbVtPbjiLtmnekwEqEvNFp8CDr6aWzNOVzQ83cHmv6Oh6STIoCI1CcaauL7keqw
33CB/UPhpTBOChINfKT1HoF8wxxwKEmN5lpWjrwwinezHYk2TtGiS1q+k7VHBhp4
YviFICWU2edJdqs1SfR5HhwP/Z7bX47okfBtsKDPEGpDN+TpgfdcKyg8JhrYqmuy
FwTdtxRmG84Ak7PpZBgQrqxb13Z95MCK2AlOLFs5WaboTufncKTiv1E+kwQpANRM
nnER+Sch5Vaguzk+M9pTqmpHWYcf1AwJMZkruhNRvxnCBkiJi1Vj4RQqKE6f/FyA
EI+6GlTXjY3UORJYlHV/ynMpeeZJZ7LyuDLLdwsIfZQm+0aWsKnXKO2ArR5UqFLH
dg9ECM2g164wyqcY6LnqGEIeSBauOPw2UynSGQflbYz6KWDgukIqoUxKeMyLQkj5
9Uwv5fIrTrUnknUUKMv4oS9sqUpNrScNP5CZjl40Wdk1ROk5BGuhPWifmWlKCGOX
xG9UaAbFaoIztcvEt+j3W4MV8lKsax8TatHHCmcsHGCYJMDK8lkNBwHYh63dmN+G
na5j2x+hQaD/11B68ijPx8s3K+DJZuCzqMIx4Q9+x86s5YA+DW19oITL6sRVYftj
LGBPKrA/0xAOE2zTiuojp/6iczgiVl3KWO3l8bKyNM3qs+GPbUcvtnl1anigGRkN
evbXNyENWaxY71lqzGUCT348awTX0OOOEZmlGap6BbYynyqhLJ/mcXnaFEcBsXkU
mS7LQ0ZVO/iCwYbr5PQwd8OONVMyU8MbuDMTt2fVSwJCpHQDz3rK5iIqwXYaB1pt
75EZleAatsZ9PrWOS7dI5ymVuXW9H9a1VLJecXmIbgCWk2AdLCTxs2DpgAir/eyP
KtMpUo0lrI1mhYSWF1O6vZzhi1472NKK5xR46pfRYuGMRoQVmSsWTdcL/idWhfr6
QnbZshnwGRUS7xuC5IxX/0M9z2dGmwQqQPkZeK4AMWsVMqI9Rat1S8jqcYB6pUhL
zMbl18Io9JFviura4R3ZGx8geVXegoDbxPVj7jpf99xiUYx6JwUKLlojW0pmEZab
yTmoarRTW53mI0IvGIAJ/JR+hHtmPjQrulhGTb0UnfUrFBY9lhBhlnrCvho0yW2j
z4qdkcb6Y8dXA9TlKa0H6MMvVJ525Sjiptut6jm+UNRC3l7IvzuZDBA/Qf6seLDc
irpVcmIgWgJ8n9uamAoJlrhx/DGF2JO9sS0Bu3+C/r0aYEqhPCoEBMWOvgjkhvI5
3zEl+uQ5gEZ+awO/ShtdQDLyJkc9dS+5dfSbtryfLVjQNay850mar/vy884xj9up
d+/DeOgpNHW1yU485WZgM95RfXlSisFMsoDVy0xbVhac/e/dputqxWs5wITDRBE9
Cw5Chr+LFp0e+RirqAknO1POH2MEjsylaIdAijUeffTzhsqW8ugy7zQD5PCWDPq+
Kj4TYPZVGE4mc6FBec243XRaS7r82iZfuYZqkohdpXlAnWeLb6OMruHpMAwl2FNk
J+OFScgLhuXTsMT56tAkQPkYypkcPAvqM/7UPKxKntMhgFCTAzQuSu+5GV9sX4l5
Bf1sqjFJk/eAhlokoibatsupoTs3vW+IOvkorfqbeZJtLfXJwQ3FzLY+Io/wz0KJ
sZi2hooLNlvePs6fweooLi73HnOCgvgPRSdCM/ZHsbWzjz+ujXiujXU0GzBwkFih
MHLKoMjWtgVfr/OmQNsTbf7dZFG6rR6EZM6a/7/29JQm3EKoDheT+chop4lKNkMo
h24NHTkF2d/nYYyZNbHliRYlYh5I6PqduUKMMg+bGwV1+GlQz01yiU6BiXJg0yJv
qKWe4zgP9T5uYhJcPTLXzknTExf7MSamaUxqVrlgMWNf+MNVmyO1h1onCO1sA9Mi
in900d05OjHjZkXYXIkfFUU43jr8sepQ4OXgjO7Ix8671zMRFDO51kdZuCqVyxkC
uEl0BgHIbacshqwaSzxpvepVDh7Wo5NU0YFgcj63ZshMWkM3zLvPjOZ12B1S2e/4
KQPBrETr3VcCuyygp3EUldDyt4yNlyGbTgAr40r3mvJrCvrKbGZau99I8/yPkKBz
1BQXrsrVo+CWzsKVPiaRB16au7a+nqU15NrCCsMAmaS+2iZWeTTCGk6ohYxs4MrH
7jELCmgeLDxSnedVDwPiokvGPJMdtSoxFhiek/v2XQ9PHbQaZ8M7OF+A21Xxq2pi
nOWDOWUt6HjLcNZPeAJO9dAvZ/lU1ZEYcntszwDO6F1HyjZkTpeoDuOsojs3yRF0
sKRqfuiAy8PNkyKLnMqkrg4h2Svza4Wqt4u6z/FtLOOhUt04lAg4k7Fb8WcmARSt
Yvxvq2aZIUf0AmMB5t7SeAd58EsxFVRGlgnPAwvJup0LBaaY1bubIGQzxv7BGfHh
LMjZQzvwya232vJSDbtm95KEjB9Kxd/nrp2GOB58P1gRdtrZlaehWTSKBuuuI9M/
HXbxelB9do8BdpT0C6BGdlsgh7/njoV8rW/f+ss24fOcC40kQ2JmpNZTiGWuPDq3
1WJIhxqqfptpwdjTmcRa9QBUIXEaTFiLaUBpL4CNP874Pe4LlXMbxJJDAUBc6psd
GbrUuBSVEeafLss1uLRSD0tq5H52j327ITBKw5mIEx0hV3sY7qNMV1V5+UrKP2YP
wFJlcof7H5X6FgEiMVjKVJSdgPJC0+XLfX7eXJKErW2OS1bKcuFu/vKXlYP48Cos
PoJ9PJtI8ADabF+g3c/XTlY0PwiVQG9i1CKIU2rWqT0aUm8qfyHW9+SmUxdCg5db
crfrEd3xPzWN8pCvfbu+/xWSv1BHYAdM/sLkndWmYC4CJtHnMCLEzNSS0LT84bhH
Ni4ZzvcXvO5NLq+IFfyXfM92ydALMv7XtVk8pvCzG9B8ovicTdGcr+ktSNLJDDVJ
WOtcBtVTALUHOLs+dODLKu4x9c1RZX8Cx6rN0yTkbFHTSR9cEO6uYYLVNxxZTgAO
2kuSv4uoOPYMeQ64uJkPmC4m7ZiuOpHB/rseB+ITwGEd6UQ7P17OkSqjPaX+hGVA
ikkj5QkBcgu0UqNXCQf+QpHpk6uI0+X6HBVALdy8Pwetu72h/QegtwUtZ+ZiX1X+
yiQj3G1J5r00ntMXWkT08RTWI9MmQZXb/wGI+sdzefLaVFUMjNz2enS2OHbUOGyZ
/TqKpOhNCniMCmNYeBL82b8npz3ZRji9OFzEyqZM/Q5wbPs30DLz4MhuDGNMPIq5
OncblB3o7aKbE17TU/n+WC1/kHoj4/TMpLH0sKg2RzqVls5lRT2IdxiwduOEhMNK
3ZEZjPw5VHu5KHSg18J4lMLlqMZJ3zvdA5ZPzWQjSjYP+iYX0ADTAV1oF43I12UJ
Bgny18VDOlOSgivXA9wzmJRxoeHr4iK22ZoY8V2yl70ki2aGk5lDOta2pgbjVstz
Pw8kxQaBdSNQ70hIfWqiKSjWxYDhILhksa94EkJgrGhDsbzn8OTMBp8pX7yNMnyf
uVNMWP75eUC21NAMslBjuz/JfZrd0H726TZazw4LRhAl9qVfZgI5reXcUSJdgW2P
cK4XwbsvWQ6myF1UVRXWWwwaQ1VWloih+BEoX6HnTBD12GekQJByj2oi+SgH6XvY
2UK3e/MJKxkuvTyg7RyERaIrH4Syyr11h02X3laMb/OJ0v3PixA1S0VJtN35PtlZ
RpDDdY3D0mWv2WKv3CE5uMrWnInxaqDq9yQG0DNOrt8SQ1tAzyv0qgs6KpEpERHp
Vm4XdPgWXT4HlYwzqnLOpGJR27zExR+VZtkTvuzr/APZDK/MrnjhhZe80TEDXuLo
RprZb+mPXr9t0eHPXNjQITfmSeTmVoqrnzn68knEiMuKHGodS9u0ctd67BDBy0IT
c8Y1ZgUfBIlHuMaQR9Rcg11MlgFS5ID2dNA9ax4gAwYnGApaXi/8RTcdSKTj/Ckg
cGbLbtaWvu18//cGsjhHkWLVahFOqReYN2nu/MVRZfRuKhUCIJ7B1yHrmjGeGN+7
prWVMH9FHjoJ+8bW1zjJJWND6QxiePSZyoX/CLHOfaCgKifyw3QbhaeCJieXGhm2
L5TyVInooWeeKrKx8mHO2G2fitVrKRuf8ilQNnGf1t770veUMighpv+aF1vp/XX6
0iuQcGtH660Uy780H3+RhM2zW7aMUnsO7HbFSVSPsp1bN3+OSwR1j/FB2kQN4CxL
tcYbPp0wbrP8wMJNYrOTfn+V6+4R3aYfyTHMDdrvpdpf7ocAuvnWOcnZTX7xYuDL
zTQT8yAZ/VEtKyHWLL6LO4eH0uBMNxH2A4xs9srMVKkrZWNt8E3gtqoEP34qXVbl
Q41rj/0jPJzSZYGBWwGStB/GlbWlBwNKF2EkaLP4wsz0C3068r6hEYeCtzCiudby
1s9Y679FbqaknLAEKQnv34yR+Ygjxn/b5s6QZNW9cw5KtdZLfa22gIe8TtFsUaJG
ww9QioiVYXWaLI6Xkli5C7TcVaKzekz7RX4qKs3NmqiIAlUVdNN3qtPKiVygteTg
tNlf5vMCIbWaYM1yj9SR3eb++hoW12cYj/dPl7xyOu8MbxI0skht7iqhJg9L9UKn
0bF6Ii+Waa7DXEbRRelBtMgWjgNFxWeHRVMNxLF0vXCWLXG1n8lRAzIYG4kjm+SP
ZFOg5nhA8eZfiY37692DkTO2YVFP/VlLFHVAgs0/71GQcx/l/1M7vfg9/CgAE4tI
O0q+JtMLFVNUgvmO0bzsV/VQRrVrgI7VdFoVIc8ASHVhW4ooKNJJ67pHu+0/n9CA
LHsfy8WEf4qUE981eYLVu+6rQr1Jv7JT+ll/czqYEqspxP25hkz/6KRiqiSHAZEj
LBf1K8wxFlzpWQnr2CEwV4fZa8CXB/ygnQXKGpyStT8DrQQJ6ygrLWGnYIZvMGkL
Y5bOwr+cz/C3l7DZ5sEqgV8Zk8jJzy2L7jadwS/3pf/crXtatYi6xFkmKNzrJIFa
Zein3OI8Wncf4tGf3Tksy0Z/8vZQpKS74DEeuKOtUbF6NJpIetBKxREhXO0fku22
94Az+Mgm51aRsFNyqwmyPvkSZ7NFoINILCz3IzQeYZ610X53w0GGm0TH9Lo1U/mk
oijUB8r0RFaM1g1Neji8qVWClJhZ8sOGoqVHaGyLiSjPt243M3AWhmIR8RP6cYu2
n+v0vjVLwze1WiT3gnIL4V6Gk9V/oR32eJ/gBAdwQR7MTMWAzkuweXq005WjuLiV
FykfzNlQFYkx2zpNpEIHGt+fgHj8GcC1SX5YO9E8AHUTA8PtFv3//vmc2uLOQ6IX
KNsbDbT1GSwTUJWc5En7pOi8XCMhspIMQGmoi4mqwVfpFX97MrfvdV7ykyqLDUrd
JVhDSeyYSHlsYYqDb1FjDEU39KVTp74BbX4D8yYrXeyAQcokWijyEeij+TxWGX6F
YBGPK+ob/QvDsyjY6fro8KcJ43C4kcuaPR1YB1XW4vZMm9AHxz0gedTqS1vWlq+t
RBs1ZyvcdoZ2dOgphF1+gCQ76yQO7BhMDE9yzHQ8msbAILBDdxhpxQyfIDvTrVeY
pdHzeuHuLIzlUVxiMPDBLnqc5CyQMsfHhuZMziRHOOem1dtq5rRbFIgdsqUTV9jG
s5LUH5qkgDbbQM2ysXJKlJs36yiszb8MB5CFV6NIjLISZBMviQ4ZGsyTc+VNETyI
BdKrwmhdAZn68dfFkC3q2+bNuHQMWRqT/ua49FuwrmrXorygYEWXBfVXH7lFCyQ1
vrVpYqiz/NB5RcHhIw/BcESOHS/97khy7cjafNV1LOpuYxXmh8JXHGHYOUbSYQyP
ULhs4TQ287H+l0eFE6hUzKe1lGxu46m8YgNkI9u2IPXB8cA9Z28oYZ5vtiY6culT
gJpTjxRqnbimQ6P7YengzM7UyYkYJ3KAukuLFC3wlTY/s0NbVpiy3NCoNJhoiqXb
sr5OGoVmzlMCf/Zl7LOaARP0OaJKNVjA0IulWBUFU87mgCyYoa7CBPPlZ3Hickek
SCdzz4WKztaCu1rz8D6s3BDKrd1HdDw79NXToZ2h8UmJl/c2/NW8+CEdplPnN7lG
luLytbJyxRJ2veYdpgO3irz/BvTtGLNBgHFY+Y7XlxBQ3y3ShUWuWE2URzQscfrQ
PBKk16/CJHsG0Qoc1MUmlKB48l2a7zQveiK3maoIw5ErZZUP+yt/5y+zNVuNkRfv
xWXriZklh1NJbr/TftJGP9iPceag4vVN6r3UcR8H7f8U9/gVLmCi5wkUCNrR5awx
ROcuNjO0m2Pnv4840Io29Z0pbl9vy1T0uO4B9OWBUNdzRBik/YRoos+CbIEdxzIt
sCFh3EjykCi2qCNMB0aJ5aBY98gpESlzmWu4xrw1hRI9lac9LDB8qioyfT+pyLLH
fh2kb+imYeSTXBvP9EDXEVxMMw656AnPpsZUHsgd6bDfagvX8p32llhOQFFMx3Zp
cbgWdK/LbjRkQ/CDnV1Zjp5ATmbMo7DasN7HaebflAd3G3Ghg9uiMJWtjZ2Yfypz
hVKyKqclt4LdczBeRXXTR5Xa5EBNSPjvq2eRmI64zahZeJzzXrzASNrv2ApOK40Q
o8Fu7lj2sHZSNwTulo8Ibghgsr/w07ig1UEl/L39u/yZVAdlhHGPTsODARBo1aNI
ignmFMpy0vp5LYleDlDdrQDF5PdR1pFYy235kHqEGaQlOGrp5SoOR8HqQeRJIisO
JD4u4bYHnJGDB2IY9GYJP6Oww1wDNpRqSZace3+ZVgnTNnm1yu7eL/H9dlmCbwb7
r9AgKiDlzm7VXXyjRx9MFX/YinG9PmN/UEwlNYeCg87MY3ythjorQ3U762Tj8Yxh
6Ih8Gd6V1mr81+0Sqqgbogu90cl6a5lZwfDyhUKsZosxEKzJkNCkvgGVS7woyPbc
aPu4M9pj+o5es8Y1ztNyy+C1jFFI2HtojHvy7ZSJKVKdhn3Ni7RL5GHVPJvJQtgc
JpcoesULU9BnDdKfmHcOKcno9iy7Mi69zr3snNU4UM1WuN2iK5zMgM5bGe4hOKcL
Cg/vrD2mitlr86AyriDki/O+2enXrtQPGpY8OM9Dhtju6aqS5DwXfcHeyOwQAHdm
/cC0n1zXWTPW5tEYJsxrUTXkGAoRoM+SFdOFcD1rDgkqbH4aLx/mwZTJBv7mIE3b
HpCvJ0hi3DhIOKTy+LlS8vVpxYKVsVTzY+N2LBQB0vyy4Hub2mcYaNeFwimQ999K
pw1VAoHjezvAGV20cr+uEJkmG5lUQJq4npW3gzIkWg9DtssDv8jpzxmQVsD6kTC7
CYN44QTwPwopTQdGEb6TD9OmDSM2+7F9FYhfh0nCUV3oPg90iNb96SETjP2uOLBq
QkNL9pSD46asjoWqE+pzMLxR3YFA7UnNQSalg1C8ejpFaK5S+jE28Nih7YyGJUl1
GkIA4bLOGOUuZWzoEb/LrxYnQ3DkYE7rs8vHPxhniBjnKfRqTLCkNfS4oMlEmAxR
wegZMOPbYC0jjtvE/bsdU2HQ7vhgJ8E/3Ozvz/FKv56HNFNCjJ8ta8XgWyoua6h4
DFLVQsyTd3zijndaaIyDKlvNhjrnbRbhUxgl0dyC3ubNJKa5csJ/0/JXBnb+pLCT
FAGzzAcSv3tzj5TE7EMhqbP3uovxI+JJI1GkZi40LOulQZy5Ul8PDStU4gvIKofi
myDMki2Okz2DmJkGdih/lFtE0kTy/P+uqQgITCrJaNFIzcHcUA1AtP3ByhixBjAp
H8OV6F7xeT0wjhxiQvCh68XgXq+omJLA8AF2GjjJ/0wkH3wsCk5DSVXADV2x2OnX
XlBMctmqC9Taep2fbD27oi69BAPdPihwzfmb6k94qOPG5R5jXTzKkVzOUOs0KFcQ
rcSSz1XVAHaZA7/xnZ0BfyXALOKKHyveZhI9yMfsyNRFPNHonlrslgWOB8p9Oc71
G+Fi33L6TOqEk5joSpkJWTaajcJfjfmy1kGMRHo5xA5n1B5QvxpHzsvfqF1CtXTb
na1UhhsaOkI/1u5lRx4c1pFThVkpfU8iyq7tSe5kFMNTERgAcDrOj7KGwDGIPIow
5dcLk8v8PBeCsQePf7Ct+0J5Gc2BCd9fzLlBcHsSGs9ZvqKddAh0mhks4Kidf8mc
Fw18vCOeD0fMZqTE69IaxK9+qty/9y6NUdZ+3Y7qUyxFVT3yoosbgvm2oviReMfC
ajN9RGup1LO7H/5+hK4TpRbfhytuxCdevLVM00A+v0C6nZksDsCaVYDoaphQSqV2
OtlM62F3UJ0YVXqMp6JpR5ow9lynUrOcWXj5p7YDdSqnoHajR0THNsbwJ6BQulgC
7vByftQQwxJW5xSRgCQWflIUyGyTsdUjTNbh7jGrVqYZlMU6DqUGLtmEL8f4mwhb
HV0hJsr3709Kgz/tle0W2O2+8nQ/4Mb5coRS7EHbLNnK2vFA75DUAugYuWIaNyNq
0aBExhXwegMLZC4aPE7J+Yj4z8kBYVImjHAmi7h/eLCwFCLHEuDdWWx4gPl0AOK4
U1TOIluX4ju3fzw3DXnXgF+U/Kyur5O3K7QUr0m3Qvey+njYbOIBbNPbjfp6Cs6b
m8uJirAVRXU0dbnOgglBI6C77cJYC5H1g2WGzU0Of9neFvaDcOE/o1Wj/Ins6zeZ
Pf629xW0D+kQm2NDsYhOcToePcS7cLg7bNYSzHoDt6lP753ytOsoReooSYeCwSKl
mLSDTCV94kKZrDTFwCG9v86naD0OP5nnYmbRFPY7qlq2ZBu/oyP6WObfyl7VFlFK
pEs7QsmUOSaNf8jEm+GbwIhCLBHU0FyqgiC3IiiH9KryqWMZo3eZN4FIIxc9OBJ/
cHjKTIQ17vYGhuFZJJgGR2WpX4sdnwvGcFzGspGW4SmDf4CkcXVtVFKKTEWCJE+B
z2XhnmYISRj7RaT8pEZzX9xSf0wkre7hDWmBT15wve+BTJOhZJMre37uD0ky83pD
0oF8WkjKk+OWyARX7FvmXubrxBTO8xer2xRDdMv+p7UNCqDU/1hqShrUVW/8/CJS
AtCrxVtV7Z3s2FfdATACh37yJ58cEKmOMFNyIzaIj8qGCL9SCvHc2FPbI0hoCEcz
7Pbgv8McwMYhEZBAuHQfrqpp5G9De4SETGELFE5DkcrCq1OGRM2hRxjIgH4rZCsH
kyJmfH/hA8apedEqrLfa7doYc8lR0WbhuFUeT2NDgfuAWOJZ1k8XP6QsdHdgmmxu
TWBzDcOKWdytZvAi1BY4ydgBpe21yYXbwzY0h6w060/ZKv899s5ZI0SxtjiNQS1S
sHuQ7QdRBVUo4pfypBbKE1pDBtlc6d5qQWBq34+pfJlB4vJyEDN+XkJzQackLLal
tuDMwfuf87qTTE2rQ7V0q+rDYYNkxK2CKjmXaJt6Q4c8Ud0f34QOSiDMOL75LpKG
mD520I3rWllLkzqKcnRqUPyxhbwZPxIV5NybUTaGec+izhIujMJ3jf+BlxLdElOV
jD4H8e4YrajbJ6Fyn3g/37wTtmeMutHV/NL9huZGVxLX/LHljXknIxtytc5eOWLT
0zcTE3N101Lb2Cj/U2fBCDEbqut1IYlXFskwvAAxeOBN3OwezG5kPc32sW5qIlvR
O+LsyqTrspNxUGBebWI3QW/3ZwITO3e6SZ869ixQXFBOWpRSXUUfpyx4CYxX4+gf
fUok414iMhtcefdiiV4qihNXgXlJeyLE/Y0YgbejP9bjP6pYW06uop3rD3jfAO70
2U64xB4U1ha+y6PwquhX3slAyZuPO1OgfDF0hrbgilNBbnvXSz3jR1l8+9DbdBVe
az2B3dbKEKYErk1CF5the0oU1KFYMojatt+xJxgyVRFMYsXGhlq+d2AsOxqHRZn3
WK6UG7ZdVdKu5D/p+MhwlILMWv431zQFYBCQFEOR7gxojfpdRImG4z4X2Hv5Ya36
ByF0Zkf6aace14Ib0i4+3EQif6+oQbAQafrfLx22os5N+SzEdSHZxLe8kNkt6Sle
ThOMHkgeOpN+v7phP4ZB5Rj7yL2cUiLYajMsF7oFGqOjdjjryrmLagWzxCwM2VP6
V6QV89mKUCCI9NB2DSBvzbidmKlVm2Kqt/Qmj9AbMxrTEhCmmRu+sOFAY9jrNOXN
eCRrG598+KGLNAInYlu8TgAt4kG/JDp6M1x49Lz7ejhReaov1pC+l0Y+DVm5Ub8+
LyVi9KsFU7dRdFxfrU+x1sZ0XN+f45YbeIcGsa0uqgN+oIap3qqyDpaDVb7qQ2Qb
hsYJT5ZKgo5OPV5J4ruC9B235eo8zJ8NIPpfn7NrN5X8d+qVc/WO33AB1/grP7fc
YSwL46p0YsuS4arUaEkmvU83oDaV66/VtYVfLnUJgw2XZHLm/3TT95uDkP4asFrZ
K6jSMiAfy8kyEuRumVucxA39+OpPDQuR44HsIE4H135X6qPRqI3Ogvc75xOy1rpf
21b5ww7FPY0CrlhvbB9JYSMVXmVnxmW+VQKYvramG4wKg0RKxNP5ry0bjV5AUmDB
HwQSFRGTeX9BRPXe2p+owgT5sgdhP1nXqN1OCEUBuo2BE+fHG9vqNdhGMJjIYat2
hfK+7yG1bRWwL7tMCQAHGeb/ixGy9vA1vJ0vWNiWPTH1YnyJcAtpSA+NOLVhWAWd
cWnudTV+fGv3y8Hyb/TNCsqwTg5ZeO5UsdJl5ToUqrE/RViNW+A6nCWSS/spITqo
gy2FmizXNxbhnDmDE6KV2kbNG1nBXf591bH2fcZk8w1rcNsfYTdOG+JW0iY+wZ89
aXnulscGJG1LTi4FvLFk4gWlCYrfKBVJCoX6/PekqAH/UQaXzQUx54h4GOIzAlx/
ijo99TOUO3QOhSkxTEdcOIjKjDiBKxoZnOTOWLy5vc1MYF0+SnR/x2JTICr5238Y
0QJfvLiDypp0sVjCuHcg0VFr6Y2mKdCGDTpbR0M5aHTwzOwi1U+JRG6zUgbpOCsP
PY+F1CjOHWansW5Wjw1ItQ7N2UfEhSCmuKfHwFXfJ/XhZcIQUHtRLnVlQ+mZyjkO
9QMibIwIwiDbmtYakmDgMd3uWM+Sz8AdNlVn7GXxZiR4DHsH1BCooEe0uzgAiPCC
vw+zNEMyljRpxQul44bN63yKAU2Hc/FiYA869e7zN/cFJYVrGB+7Knlt+C/KgCLA
MVn/kOVlH8xuQEpOMOHWmTbSB+NGq98TD95/e6bjIZhD+h9Cdf5LPKFRdSSHdK2Y
LvfW/irAOP3FX58mEte0fDm/8x8kFVJkeh4SQMVQKGdW0Zrj+Qr5mIe705uzGRaf
0oB0AY//EPu8NhdkBc10q1CgTti1g+s212x8k6G8iKPPP0b9TfxM7BZhZ+ErCBlW
c7egTpJvU+doNIVxrvaHMDPUwXASjFAhZedZ2OwHadQV6Z8yU0/WfymqsZMMat8E
0tWVp/KeSsJquUu8TchT6yg0xlAsw8XdqOmhLvexkM5G71K+EYU2IMq9JF5gqtuu
eLT5hsHuZloEYYTiDRHH8zBVBOYiKAavY/Ff9sfd07SNrJMzEjY0RELM1BEH/YkI
RUq/ssOt33JZk1SJB68cpYTA3cOYfh+/bLaZE+xf2ztd5yUTo5echGjGNaA0zCrd
CSBF9VCXmuO0b3+reo7mk/hgYLJTXj27iXWzvauLmvgIxXGKI7zhBRdhEZdS2gml
zVh6v9+/EOrSftGsD9HnzsBqcYsgEsohNwPzKaagtsDdTcWzW1z5AtKPiaGMOSGB
RnrxBvQMUODBb9AOuX1crxwJ7dE8oxDwuIZO25yEouPV90skNYcE5F3m83EZz6Ny
uy+CJx7tx+hs/w4SBaqfElBmDWEylDzml5Ns1WQWhz3k3g36bmet4EXoUQmb1XPY
d/llUbKd2t4GPfzL7Vyrjb5CPz7eZzUUXD80xFKEdbps8BF8BhjlMBD5Xqx7d/3+
B+jUnzxXGZ3EWxYhZyhgrgVRqZsyM3JLUH3iTobSlbe2PWHmydqFVmr2XSDDUNkY
PYx49t8wgYt7eLMkdOMVwRsmsXVxTnmeliY/zfIRmDk6VgyUYwsk8R8NZAK1RnOR
l8W3x+oPufQjodvZeC2o/WrZiv5TxWAkLz2yZ9h2z9895Et6MCBPb2fO6u31HaR/
Qwaxxv0SDgig8bxmv+t6XMhG53PAOX8Ibt6ZGSfVnb0uAcXGxb29z7miOxnBgo07
p8s7SOud4RQEFptnTkvhJD/IzTCAn84NCWwX4B9HyJ1nsW9fWWdTEVXSkjTBzfyh
cH74U5VwrAhjkeqDspkUtv9wTywRuxdOoqHWA+RdV2UDaaB9Qpta5jTNpk54SMMO
duIN/gop7jqqdGmOTrYZZqUopRsOVfjfJngrMVVG8fvEf5oN3V7hOlUXyRjb5I8V
yh66bGpwuxbUdiQTzWTlpIPOncoLLZw6vprmy7cqz1X8cCKG63cPdz3iFk6jabMu
0BgIcavPQV5QCCEzg2TlyoNnKyv5VWZ/I/JG5Nfw1nZyLBHyF3EWR2wczGfoypVx
HwPcuG9OVu6B4s5Qk1W8bdTB76cH/+PwIN6OVZZb9041G+J4g2odDdPHqydL1EKv
qwIPcxCbshY7OdQsO/+eYpZY6HNi1gnasa1gz97zIynZGW5fvVsaBhvSlonoPkdI
FheOc6gVCYBcngpym5OsKqBnWih0ErliauXdfbbe5chaKRDDOMX5MuFMH615+XoY
t+AbhDCAvBcYmevMe4zMyJG1RaeQgHX2N2tjbcEWItacmG8cJP7LjTRgDjhyXa9Y
fruSNyXW2ejYm7+7liRNh53h54Gdrz3FOSURkENb3y1PHR7h35Y8IrakK1jI3cLN
i+6QUfzykgMIF4giDJglrclxNnIs6KrjtS9h4KL9wU7+15SIZhW+88y9GOL4zNYF
DL6c4DJ3E7ZvrGqlOjwffoa1GsKrNoxRZbAQB1kNrKpYx8+ZSMHbIB0FMylVJCoq
lYXNNBP7+hlooMWItLQ+D+XLYSyr4L5OOD2BcIAVWObGkpz88TyqmELdboyMXScd
T8D7BnLglXIE/yU9LjAWAz71JBcwraSclXQjsf15Kpnzv23OHQxL2usRGbxOKPhd
qu4ArPcx1KOigLuVAZBzEiKwHnRm3zUgiu3g5QUFil+M+qlCxq2q9+8wGdjPzU8N
OXUzRdctznx3CsG/PNs/BBd9oqf+tXtgH90+Rf8jQt9iH2lMp61sE2E6R9MQ9/Sl
ilXfQg/cZ+YvLVQR3ZobAoVSaKp4InLA2zoztCy09QtIqbiXhts85QMmwsjr/+cB
3BhaD391jzzMk837MouQaryyynQp10RpqifhfI55PLasrZ8PBVt8spjrKoChwUfv
H9HeUuVMbT9hxCZD1Ms3OTizFdkf+yGbZgW+9Rq8SYCUruhcWkkuzGOTvRjQjddU
GMGzdFxrGs0QCx9pbvmeMh5TVChny8aNkqb9BDCtQrXoEGqqPvju+WLnTvHNzHI0
WIvAASeyrBBzJ8DtXQ7q3hDQ+9DoHmD1sOdQz4vCpklH9FxLhF+EVGFPJwGusd4o
pV9hCp2+h9ROOXwmAkQWfVlTmsncRXmL+WMmDkkq0uqVX6xiqoaiK9PTbKDicGIb
gUe5XpNMsKsNhV0GOnFWfVszV/hCgxfOSAFIofJJB8769h6UOTUG1CEncVWElHWe
GzK19f9k3qkJtJ7KIXepB/vYa6Frv+8Zu3S+rPEx+j8jYPPyXxc3UFalNRkVjSOt
yOUcNCNv1Q4s1nyaJnYdJ1J/qrUUsdzOtJSO5f797sqsU7ztj1OiPfBcWGtgArMa
odnTjb7ZbvmnYbU6+4r/Msb6ueOStlzbY6ITt4tMQkozfP/3f+FY9CuxZffeFyfj
XZwX0tGNTZfSRivz1ePCT475ve4lPB15Up8sFmA+eqVgqyCseH517zRQwjJAyFBM
wUNxUVz0VFBIx9n14g9hROpgutoQYEkd9RGer4xkT4L4p9eEaG/VJLeY076sxd6b
wuDfmKME1/QH5NnufkDd2uqAQMyRicr56uTADGnlJWD0X3ofvd2VCoQHd0HC/J3J
I1oKIjr1JDv5Ot9lXSAwv1HEu9UwA+VrZLlJO8AD3hz9AB75wdwbkxVvybw3tTyD
0yF1aTptB2Lk4qvKPwY8zDblrdwfMI2i8VvZK+bT7cd9+BI8WpJYV4DzIuMZKmo9
1s+ZOsner5Y3ruT05S9DdF9qZJiXeq+ddUTLiWRgoRseL9dp5QfNZ0sCLK6oWmrK
CMgYzI98S0XhL/2NM+ViTrI6aDRO7ihs4/KjMp84fXn4FZthq1I18lOFijzVSF6E
7u2ntYYgTluc7S+qbcEJxPaXFwbFZU2amxXAVE7WMBsKtiKxlAiVwHTiSjWnU1Dl
Mh5O3U7b7RzvcEPW9Tx/LAH8VlEuKpcJdZPmyxjk2yibJzb74hKHY2oPOJaXCYwN
Pbig8KmuVsk4TqRf3yszrat5RfW2K8hBIpRl3Hi6KATd7z/ui0VYh16nPyHwD3w0
HOb5LaWmir5AWCCozfV6P367mpMWJSHGa4K/iA6jm5pHZzjE7mv8sqdejYNJkfK+
bVY2tjUur2HP7xIdM6cbdxh1FsuYvgs2JNLuYRJJdohdEK9SVJ8UlkIAOtFajQbB
f8A4sNuTE/9J+MZ43Fd3jKUjoZ0g6M5VPlGNVR7dO+4sPyioalUM96h3kcg2Mg75
VhqGPu2PHFRas4KTP2tehPY1yCUXXQJVleOvjbd4KQNhmk/Dh9/oPaxEaTy6yXI1
01+E4vTYL0sc0gyrb9rJk6En7NsTxoXYBj7+BtSSrXM3NDlQZS5Glk8scUADvcfU
i1XYohk0hjXAyjC+4t9MmeWBgfbYCE4hzLv8GF2je2t9phh1bYFqA5Oy2YEpEneq
9FWHWwpx/VcAcr1D09JWftX0MLZ8v+Q1hRQiryk69K/5ES+Q2hP7aPvSZN23S3ON
QBF2c86kAhiIr+CnzHNtWYvw0AnQdAoH94KQwODP1LfY2TEY2J0CMUUuJYotsayI
xTQkepjHveIQAI/7s0tlgg6mbbxJ+YRv2ldqm0MBw2IUEr7w75OXpPFUG34IHpvN
BL7H4pHG+ZMxcfT/VE73jRAsVduAl1snPlRz736eKdYDIjeDLgn84fJy3F7bTE1O
5DSjJKhCrkpMaYd5rniofSpsZ2zcgtiF12e087FRykuyIFV40lLsXpwkgHHGvFPJ
frXIbEazhFAoB8EcTN2u5LGOJLr2SEf+t267rVafowali0YSYqzjVV3cSTXcwEyo
MfzRAUdO/tBqD1H62oSyLWmAQ13+bwsMGATChp0nHc2n3Wjsx75drxaPvojQ6Qjl
TODglvbwQJvYnlIL90KkRCKNBTKzSlA+pHWmFz52O+NiI1DtL1Y7y0Ku4rI7AJzi
duSSUqHfjfeZ5kMmIIUfDGbYLaTh1DWXgZSjJBJI4CrloMxWiX+XCJS6E3aw0Zez
atGdWK+Qsx/y+SwsbZzlG6Wru6jh3s04iWiOQ3PAlTVFBsyO2vX1BFxzBDP7b3Bz
lLXESe9ZP+z5J+zU0PKd9x36n9BFlYmzVdfc/+yoDMpvufvVhcFAQrjgVZsmDe3F
INa634MgMwix+3a9K1CGKqn9DbO0yZlxegqAWwVWTZ231QXQdettBSWyp4+urcxK
GEPN6jtadG3R/7jCwbo3w1502GyRdqV0jwfK31Bx9fbYd8YIqGV03usfvWcmDJ4X
tHERvNAYzfjFpYXjSfXuOwyR996gh+TROhV6I1YhgG0NHzkJ0TTwm996DZ3tRKQF
VTRod6g6KaansJCmCuQb6tSwTqMb39BFKXYX07LRjrQ/LPMZM2mOB7Vu5eSas0AH
z1iOjd7XSAk52N/Wr7dUb0vy6iPmF5lUKXMOKSPHHck1tQQk6AKzqGtvYHtG5nmE
Guoo9xqOjdSTmi8HzGjUMM6HgH8q2ZWrMnhbaTWnZgQ87+BP8vIPoFSW0sbOOMpX
5AdElRIGQ9ooQS6E+ITLJJYf71wTnO+UokyzsT0pJSW+Xev87B01ZeJlmm3RzHmS
Ks8RO3qz1Rv3d1cbpttmm7dMAnt64q2MW3xqpjdgIqPvL0acNS2J4C006uJymIt2
AuoQjRWHqZylyprYob5OCDZXUsWrh/1Gdn/wNPCUHHpQK4k6aKA5O59KVcjtfZRy
K+As2cuxEtKgMCBmytl8tmw7cdJFD1M/D8AAf8dsDdw5e55E1k/Wf7RoCjozjXJy
bPnkFvqTwRNU4jFvhnBJTq0tVDvARB1W4gsJdcSAWkgCmNKvsXfIRlC84ytTJHc/
wz3VjNmVf+H+5vX+QyArdA2RmY0N32eLG0iI54HK220rqKcOvrcbkXXDbUnC6WGo
hq6OW90blLpKqClydJOfUUE3F9ez7UURUQNcye9i14b3bYvU+670ml3DQzET7INj
uuyl9U6qPwqNXWvMFfhlsYBZ7vo0i/vAAh7TraH2DNmw6uCL9azpFEDsUfmV41iB
SfwO/KfuAqFi67OqoLunQU7svAbkImNP/HoVq7Dlbg+iM5nbcgglTOf/oaWg28Ar
YzxOoEoZ7dzAmwcDnEHQDryTaaZr4DzfI+/QmPBtDUb8giSW0KsQm5F2H9DkNc/P
W4v4esFx2XmVNqX4Yk9JLC8IIOI94DNFzkT0Oj46BcCidMVbcT+RnLlY4Fk8Pv0p
bPxpQj1vPu99MpCQsE6DDx3CVhfvuej+Z82oXAZ/x2yh9f/Mgw+ru/SFApMrzmnQ
PlO18x2Zlxm4ozKskAAXu/0879+C78NDvDPN77BIuKCNjX9jiG1i68Na6JhB6L11
0ldDuIIRcd2e1YY5WpEcbWNhiR19VTptUXl19ira0BJlrc17mS2p8nj2lnAt/iDP
kJw1zxs3HWkhDzQWSP8WbZYVSvWPLhH4zTuTU5TrKsSvt0aeRZk9cIq4gCtqV4J3
GB091otY+QJnIlSXvVGypT+72/p0FtArQ45YRyThd+Q4UB1lV71zsvgtvVC6tq8a
0MxGjyq96j8/GdejhyDlb3VOU2yu2UnC408v8Nm99IXotOx9VfiIo9kUlJ3RZgYo
C5DtqlRLxI65fzoZCEscEBHRCqNaw/u4mnJ9xLekpTRKbmIZsxUMqGheNcb59mHy
eCflhYrMTxVfIXaIYqWHv7y9wQGX+sT6a6/B6SDmDADhuYIbPCgnwY7Tf7bZlQHI
3LthCrI2HlGMZRMn1xNdaxGcPgV6GfH6zpvJjnK0W9CffIwhFonxQa8Qty5Gu7eg
ZZhUOjsc9Emv5a9PmvdaFvCUyTQA4132IRIWx1tWoDtYhZ79r3hKTIH43yQytdiJ
gG80DavWtc8yfWGj3If4S1SCX6A75rbIGf2JhhxwgeQQLOomuvcufLOfresr5KZ+
UEZyBRhW93S9deoXNhfIPSv+A/7sympllFhwE9u5Loj/WsYVaPeecUorgC5y38Im
Q7L/DhXaslVisbn16xVCRQddqoKQBI+ZnXlh27fMbIlrWC5iy9mocqMQeehFQRpP
S4/jkt0cZUiAWtqdeYoRy8442yvvUbfCKqitlwGZVP0h2ken1MNDKPN2qIqkNtYn
qk85Zr7miKEqIfguPNgvDqT0OWZ7fKa4hJ26A7GJJHaM+JwRudd94GLgGZE/M9D7
6GfeVDX7UfYNWaw6QW1Pg2KtyJiPWC6OSRSD+y7zvBWU9YMQq5LXlKBSNdCF+J85
KCZFeKe00o5nRmuhlo808fUySvB8YjvX4glVv3VstlK1E+EYNG5mtrSRYkgC/Ykj
Ji/K5m8HXo/xMHBL/0Zq6sQDgAlMaE/1PWgz3VD0cds0zGz7AJY1dItxmcJT8yBf
HTgRinlPmUfkUT30rvcbhJL9CW3C4a3CDtd0i9L6fGFNN3cbzjZddYkcqD98nxdv
czQ9EnvAZE91jHZu4+x0fWZIOK8ggjMOdGYcvYxhJ7acJQZCDzO5DJdoVProS+bi
sKYx2zPB3Kt+7GuxzxUOKmwfH+aagv5BJ9zABcvlY1TzSUdOiRNyhojCT17ygcN0
6gdzpfq+b/oQr7Wa8z8nd0AI1yP7nJ8CgdpcTOlshWcyquCwKcxeVvenUsxfTauh
qZLBzGJT/pCqvsaWSxMVID8uX6cpNv0EVCc0JVEB68lQIdWAfh7mBXKTHd6FbpEq
95S6Vu10MA2uqaDtsOqXImlfc2UOqgp3Y5JUoTYiHfK/sNckrOI0teKvneGjTDRu
I4x+tdtprpYVZ4aIQkC231k2zYOfLyRz3brPHp1lkkCoo5ewh9+8Gze3BgMYwSxF
3NZHQn5qNbzlLYRXPRpARF7eDZzEU0WLX6PSHHnUXUQg2TzjtyXngFignNc8SJOk
GDl7RkF7wPcuKcYGxHacCW0pAAJ/zEY+tG+wYtM2UF8DdNJZXmaKCOxaBxQ0gFhX
NEi10tyCiBT7lqkjIpBcve7YQOrTyVW16GcHrMgzl2DMnEwe/Q3OUmP3gP4Kt7Hh
D2iBXMekuFA4fZaLu5b+pDD12eX28P9oxRnTT+QRE6mjnwU+dq4/4V/1ROVTFgtY
2dtZAmrWLQM1S8L2M+PjBSY91D1ZiaDlv3VT64fs1ZLZOR4boZGJ7CrIso+Uz/Ru
l5dbV2k87efLOFY/WmtRwwMbPzi/r216G3bJVmqthWemdYgXYAhWNMLcVza0xkXO
I56i/LGPkQ58wOrV2/qbAeePk9u4nHbNwjoR0WydxTX8HPEmZCqZv512c1ZrZWDx
ACA2I6bnE8fjQzhq6pLUNasFXyMvbYY8bbg00t9xOrRJApfQH66MAr2ntRRKjl5o
yd6CkrzDa6RHof1kkSB6lHZLVmL4gYONGEozPSvb42MJmbioaNDf8k59+5P8c8Kx
HKLJ2WoMtGPEXoNnXw3+AbL0nt0rwAMg9ONgMcTT1oGXcINajSe569jWQeuQJ9iR
M1iYzfvEBSQxA9eOCcYt9sqvArx19I/EI7cCb26eyoULsYcQyoJDvceHM7Y1kJBw
ZVuYxwPXJebbNdvOYbI7Af+IqI6VBPcskbyvbGv5gbbbJ1PBYytIooyOxK4O+Bbe
LiP00oGQBYmfkH0eVIstQ8dZsQpEb2XaLSO4jWGqKosmQAZN3/cRhlTqai4NHuUS
EiYrpBijdwDwLY2CgaX/dhuAT8VQWtx3P8q96GnPEF19xHyebHzViMGK4vdoe4nI
m6B0wUNX8SEWF9WFQrZ+mwkIcElZ+qnUafoWalFDBzsrQWxRPi0Gwo/nT032Nb1/
tvy5S+FIs/lnD3+W3Wa2hB/ZG8tR/n9FhsnZNClgs4TmrK9X9kVypF1hXOH0pGP/
ZmbeBaydB+hG3ObQ2qqHHufnV9y6QQt8d09C5NrEuwu9dZWGZvwoKpG+zHFrcgtY
iMMTq2PqStRbU+Y+vAXDVusMtJ+d51ZN78OMIHphy102NX4FBQn2AM6eD05I2mUN
EcLrl4p6fOiTPiK0nB2pkJ8QctdGo1qWVodGhaLOAPTvQC0EFdTCiBxr4mqLWG35
7uOFWdhNjc7CLUuTjrxb72l/ZG8aSgskUg9zqGfm0LyQk1KSl3vQ8PmPX3ftgtNg
BcBJPY5Ml1AshOjc6uOzZIExibbH32udnM/xA9GEHyJ8guN8rVkNCzK0lerucKZ6
bfqXJI0PAu1QO/f32v+mhvFZz7BgI4VP5G/Jf5kU2dMr4Q+7HhvBfzFfc0+zng8c
5nb4Oe7pj4SyO+Xf41fq0I1j2LDdVoWWsTtWhiyx/3xRzpMVTru0gCcXazp+bXPR
2Q+UvyajQ11z46jMqlgDfaycl6ZdF91XVAetFcRF2r+dimbgigoeEVNDx5HRapKZ
JFU2zBn1QfKC5dc3QbH3d4OJYWPJOlkIXsp3/LtXd1QaZEX0gg+tWEiHbJHFT+ND
vOQk62eaIhK97J3t3MVZEUJYszUVPxOA+dSZHJ1gyUORTIBlBoPnle3wgp3bawcG
6G3U5lOC4k+hC7PDibekLbelKYsX4CGqp44E5yUaBu8Us+uKeToqNCAaoQAzytca
NB2LOmSh71wd9iRpi4/XtqWRAchLBgtRaeTtU6Z1mJ9xN2ybisbGczVFIWHsif6u
MezjqJLHCF2ETCxHjG7glNzqXzOnt6ORTvN0aLFboc71ZVM97eE0ES44txuD/Mqo
WvaMb5Iw063x8ZEM0LyoKULeIgFtrejAiBwVKAmOHwJ6SNisyXBIu8lImLdZ1o3/
wuMd/IKM8jkUBlfXXd3PaFoxlJCr3Z4AA94fTNqJSNkDHTOHEYPVEn6PS1oDJyas
jeAXmo/3a4KKlDSgdq06YqYKuQbw5cyiiLXyXmeCHdHf1vv+u7g1ORvSesdG+DBe
ETV+l6twDdJ6kCBh8vGtNo6r/OTGqaNSzrY3IcXvIbJBxA6tG+MM2soiCrYPZ5oS
n4JcLYTxlvdWVsYq9xplplXbH5Q2S1eQWj9Hg12e44eA1Db+9DrAKplhF6mVJrYM
clw9vnLUixBvfB0Pnwirb+LC4ylBKMbnJcvaMO0Cox278MLjd8KJp93IsXdKtU4C
DSVKVu4fFEgq0UHwsHQvIPeec7h1l3KiYtxRURzK01I7eo+LJs+ctplv03PlFfNQ
VGGxU2qdbWaIdnWx0gH2Fyx6pNPpxdR8l4X8G+hea0X1xeVah0cwF/IEpT1y9tml
7oqxQpzjwKwJ84hB+C7NLTr2uPmI0o6kTFdoy7Vpdbr2gSh+UJXwFnBKfKHT2nTS
kVlolZg2XxE272+OMQHTOtJ9Y8sH2/dOIjafl9veSqYUu2HSh1Hp74EuoHeRV078
JQjfvQayc+UDM+im5dPUHFYKFYrizy7qJdarKI8hQHWWRnduqdF9CMzNq1VW/uE1
B3U2GiHxUcVi8ZN5aUJgKwSNY96ehVReXldIqHrzxSd3jiuq286CPWYccnhWxhZC
glA0Nq/wplwh20ywqUFCuas980nwaXt2B0TOyWUM3SEgWY9el2YvzMRLShXOyOkP
gpgp5WgrAhWnvTp7ixWxFR/htExxpMJGLno3LG0C6vck2WhPg/gy7sE0p2037B/r
4OYsgJBziTocdLXNfHgRMyGQ5wkjVS4jFvjmuHrnefWU9lyTb5kCfVjj53V3t3yo
WCmJE9tohKnqpPIC0uzIFr9uVqdCrXENC1/jagScf8LcCGNOMXI+4d1V+AFbqBuH
iNRiv102jJkfcn8SzX/aHK8FFW+ZrrEHc47T2cfmwFZ0R0Li+PsVKaIkRE3guBw3
YpwJtgIwDKnHtZCP4zKEwroK/puJF5orIrft8Oufvs1lx0pexsXJWxw0yOIFAglJ
eFG0C4NdomWphftu61PtR2/8cTn/EGM2VjKHtJZz1G+8e7UgMW/75kvIViMsXu7E
Uk8GwbpH7q++g2pr319SQK2+qqEl59ZXJ4K2kIjzfwD7mMwbe+NwyTgCJ2IiodeC
/voqm9zKRo+pBDp/q/ksHgel5wg2UrYDH5INCc11+YNtxwvbIDmdQYMqKFA1k+m5
IqECQDvrfaiJogLtDYQ3xhb5Pi1BL5t+4sCmH+co32NOwBjCHwhayjeOA3r14l58
mPTqC5tphVm6/btS9MvSetGV/pxCxH3B8JBJ/zxj67ILr5x5HOhMd+k45KyfxXDb
kMm5NmMVsU4LnGAwMTMB8yKUiOnmYfuXPomoB8KW3eD6dNalNIm1zMv7qe1Kb9ut
LJOiMaD48wMKTyH6cbxjHv/ibu68KhVmkSyABqWeHu26VSvRiHN7E2j6YsnUdyeU
wHsaUdmBlu9eSZDpTDiGehiuQLDruvbEVIfDnpcJGYwY1UWm8kwCDjXwwew7VLDj
BsBmESljw00Dv6+w64We/kdzJqZN8SSXJoMGZ+3MIc8havvU92ho6s/DE1uisb8U
ljvg4Kq+iY1dvmz5xsMSaEAyJ21OhPRfzl+aib4+Lj/zW1huagDLmej6qL3fKhT1
MZszx4BEmw177FalSFXSsCNYBZeC3nWeghpJgNQACN+/0TVzTCZ9UquTO1mHpy0W
mg0eKFU5lSWZfRtgNbhRnDypqJImeBPhXsFJb0e/jRXCpIUTaZvrFrabL1JnVbmU
Ml+A6CroyuSzzfClIoKUwuMEwRtdlZcJZxaEhRo0siuI3pEcfAOmopYDaaWX+t5A
m0/OD4kd9S4zK8VMEk/IoxfvDaGrkc5SYw19pPPb/XXIFcki6a+6X9IK0txR6Dx2
GO+klzeCxgxp0epkRLRQ/2u6tovK71pv03kirsSj2yIsnxBTozveocn72AXXCC2O
IhYxQLdVREwrja0N/7ye2EAl0yHX9SMSDqjqHrAj02baKXorVwebiRxAqenFsecb
accu0uSszbfYU9YxKKxvPY5mG/gnOKmr1IHBIhaNNrSfQXK/sF5CG47dSEj8f0dJ
VEUMXgXEl4SuzIAclurJLLl5t2a/Lj8Na14Djy9PPegDt1ldXc79c24c/2VWowrF
sBo4yycNzCNpDFPJ3YmdfhBG+nDtoVz8C0b3qmrE3Fhiv7dUJ8fIS9kLH4NSLQ3R
Zoa7QuizW92EfZmJ1OqZ55xwRi+XycU5FvbzIy2bTVLa8cLXXRGcSpYBuHf/ZBfv
NnO/yiAgj6Uc6FNrPeGlOTLGI0k6K1PMzGEAGdtrpGgFFHoB2aT/SPl0Iz5Zzb0U
TPxzkOPZwDZUbWemACxyjCEVj5bdQTJp//fGTLIQxdf50VMBTA8Ew3Lb7EElzE92
jdYvwaf97teQp76e9Oqn/e0Dbty4qtDshjSd3aix3jkdl2rtmt+dWX/9FsjThsdD
4qQ2K8EGnZT0/5pcmVRzdKOYi0OO8kkfWdXvTop72GndGgqxwNzhIieGjx3fHD6y
SckxxypDEo3Im2cvDqnf66wFqW4V98KNItTfKyKwNzKSQV2/Nr9cp14HB6zUFLtu
P/aaqi0xJGFXzOZNNgf4GNTZAluG88iGRGOBolNZgGIf7SOZtpZdvITBQxVpzlLn
EdaLzELtSX3a8P5xibh94iN/jO24anZcmdGSPt8jE+fQUqsI0CiQ4tf3IHc+ecTk
gMpg0Z8wncsFbXwynjiHRMizYqugi19yebzQBUKzO3O9vxthdhOVnb+V1G/plMaS
gpSJSVEIR97/iS4S5GGRR72Pumvox/0RDFxCyFL7IZvD6QKx3D80++07mB7vhkqU
WeaqePlRm4OiRXoD9OFMPtFAAtQNBKFPa5oyfxHoa35i7Fzqh7ZLPnvPel45pLOk
k33cQs0RQEJCqkjfPpbAKq2kCbJwuYH1Pg+oRrZbknr9YCWBnGkK7NpCoNlIU8pG
xrpoaEIarc5e39M5cymzqidN1ipT407xzc0jLRgYvpwR9/GudNcO8yWDkGgRex5f
oVI5GtMQjTgD4rWFbdF3o2zg3K+5nOVWYwH8SuSasLBOlygrDf3fAjLDa4U98ani
DLEARkmEzlhvOamg50HNZdtEkrAiO/rJ7aO3CzPo9JiBtrQ6HKYD9gZcKwiGB7P0
gs3/tPHf1qEDLezIlmm0stOGqOfRDJjbsgeEyXZKiDXNes6sX8aibIxoSkR3aZeI
LxUGjA8xe2km52jBE2U+jyTISASNrZKWdt4/F8SFUHHvi/QdFERpavhBVZ5f1jLf
4jf14Qq93y8NmkkUmdv1r1dRVyUgCQPLUqRVPeV4RLoEFkmLF8EL2RlbqAd8zpP3
VAso4l+ek4AunEdpxscznzwkhq7ky+8JC1DlnUniXAnqrVmYqOALjsEjLFYvMpzm
SjyE//kJFtOgZoPn33FSzn0pSiq2Bf5F824ZSuDRnEMi57uH7NkScyJrpp5eYnBT
54fYqqBfSufmo+wKEWPB8RVrrvQIha0iO31sg95PN5/V2nyJWuP+XtL4LjUpLo/6
6nSrNyII7qJk3UqnmFTvxelAE1W3iOdS7Cd7r9J8IjcOJw+eDKU3bj9n4A7+HpvV
mNuAehIZ/nIA/eCIlu/QS2MXsGpnFvSkiWMgWGEHGny7Ru+eMamQaGq8EDp0mm8N
u3rF6cmv1bpQ/lRqyLMs7tnkmI+AhletRvzhrtt2iofD2PwxqGfoI7vavhAAPpuq
WTMRpmg98MkTjYWtJlOH01jiNgQJarY8bcFZqB6sBk3XLzQTrH6BeOonuUFUNWpD
oDdUGEe4YN9hJe5PAGAkFj7W6gAXHeEJ6Yr2dPBVhq5EGFhfQqDTNBMxBsOVjiSU
/aMtwk4nc0FFyWm4R/DRYVykjyB7fZqCa9oj7jvyNMiTA0pDn4x1F6nED4ce1P7h
83HNdmTjmIVgfVClxBpboEJafiCehbQmejDMiDFHjYHE3zuaKVFZt2VhHNbtpWEU
lCHCpYrwpsYQoSqNJjfCo4zfW0RBUkiqelqbW2h1IKHJnNo4yPgW83eSSlfV+8yj
90kZ7akBjYcOGwjboTUPzd2Q4+owQ3fMOkslYMlA64qgxu/Gazk5vC22b3EANJSq
a0Ix6CoXmuY49znASEB2ukzPCJ3ew3o5SulZBJZxVedPEyy6aACUxIHAqEih/d9q
cuquRFIIpRLMGhIymEQNhkpdC6NgwCYLLSEIETRRzCGrqD4U/OV54VHLFlSBGk0t
C88AZj0t6aHPSb47JClf7SZCg+pQAjSrowIMYHusO/tnk6RNUQODsgMabHd4BtnC
VFKUeCQKLxWLf9PSnkToIAWRgC1R69zTN3fDXXf9PxZdnmJiEFoyEbg8WqQAuPec
d2gBBsARQxy4r7LFqS3J9QARS/TZ2gVjvqcMyQNOvF3U3oq1n8A/Wrc5fNvSRGNx
R3NlmCDi/AWyA+FaaaeAmjogblxP7cl+ifn7nYjLRGN7Fwo/ukWoGWZ+rzrNMfBS
1ABbkYdEeaY6PPufAGf/EyYVXrJ5nz2A2xRcVybYPBVMkZFzaPP+2K0JeaLHfdb2
UKMvuaC4MZaME+HqI47L4Z64Mvd6TsvxGssxyvKcRHa/+cedgsrQq0b7M2UQdEMw
VxPHDe6voN22qASM2Mku6j7TKof31jt9/X4YIAtQaBAjP31nvaB+SLAVdR8irhKS
zkFj/6cXaA13RD7BfBphUCvOBjQa4j1vBn2PF0hQ1JPgIvfzhhMt5VuY8dejTMso
mu13DoQVzxZ5BZg/SsspuEcJjbOcw3wTS5j6hLaKBPAPp0gbf5cq8GweS/z5RJKQ
nWhNokjgbi7bMYhB2K6ImE/idhL22BWNmsACjU4zgckfV8y7NVxwg4oy26AjNTjZ
LXHHqh5Hyuq7aavxJcbwfM7+61c8ayZLRpx2nTw7R/m736Sqk+NPMAj2bI91Wlh/
SKwkeiiC8Q5dG1rZTz5kW49wPJsW/DDWPXT8lThtO0gIcXR7eogSYVJckeFNNHX3
hblM8Tomeif1Z2Jnu+kD+tiCa3/MP40Ob3+BVjyVQSbR3SNpkwrimY7OVe8bDP4U
v2u5Q2eEDqIZLKpFHCoOi5+X3sjTCKStl241mS17ZRpJUtxm8LF9bfwTSU2vzDNT
4ZopN4U534OjLpbw2ezCenByoDM+o8KNYzsZq5A431obMiXUh13wgB8CcuSGhRO3
gPkiPEKsefqdsAPu9QOx7cqbRjH1CNcbQMFRh6w7bMIcSsphWPL2+RJEYsugnuxM
6wgq5IQL5ptUotjua4q5oeWUIqf9I2ukNCWDZs7G+D7pamol9Ph5ZlNykkJSehgc
jTUx7BHUsUNLSDkVxacC/QEORYUgm71oi/K15ahLyxAHITDelGPex1diVLphVqA7
NVRxHNkdqDuEmrp6JM7fK9DBrpZNdDdWawiF5JAF7MTxiHsgUil6j2yfh4JpUQXz
Qz8eXfLrCsFpXsO/eYWqW8B2yl7gWZETw/JiRduyQ71+OfPpUBXRzzBVidlKKfpJ
hx8EdImvb42SfNmVaSk/QTTy76mwW/Ed6k079dEPK/vsnajToKB/lC0XFCUPrbgz
otu02fcHbytmWzTxNX3XqE8yfTsViqAWfYX2fjRi61L4XG+2OYC+k9LfANhT9xsp
ZmzbbW5W1aHPJOG7YpUxAj/0EjetPzh2iXijzOgUuY5Oqcuqy06yEYuZJIyVy1up
OWVdy3OIBeO8gnO/iDdPcWe7t0iBUxEOis0+S7z06B8vn9Ul6vpdafSaiRIOPBnF
nzKL1H05Q7PeoE2LpO2WFfZJw6W+S4wt0In+lK9Uh5JfZNsSTuqu+aKybxaCX38x
ZJ/4tx0K2TrEgbbl4Q/3/O0viViiC2t5veKoCINDOBM72Zu8T273Mp1NaI1xk/AP
NUdvVKfGdo+rWigvapzc+HSb2MAJ9pZ0ekUg83Hbu/vzYk6lxuML6QpXDn4CCACI
N5BzrtZoiSjjWHX7hX0pvy3uCqYPj3HbnaNl5L9h4ZVm423mnEMpRQdr9ixRU9oy
evlWxsJ1llsFwaofBnZg3xDqmUZFOcyA4nj0l5nx2Bn2jqoSVhQFu67/A4/gTP5J
QyKkjW4fSR680nqoqV4I+6kLS/2PXAILMYiOpra7aduoD75GyA1G83WSCDIVY0dY
7tt7X0jiJJy9vjg4Wf9hKvLGiOdGx36RZOYVUjCv4nGXb5ohoDGml+vxlBwQc/wV
kXGou45pois2a3xj5O9eRCeb61FQU5PuLdrQlnuxULAZobxf6XcC9Yle+vm+aHTR
wvLYtN22KFs0umOw+X4d2jzzhSqKZAOZ3CYQNIgBB+EqcwjlRgb1ukWw+2RQd0H8
R/zPf8z4wGqYpD5im9EMkNsXBVLweeug4Bz39/TPt0YhNEyyZkkMDz2TmcSsIPCq
iJYCglZ6LDwKm7AnyupSKAlY6m6r8Xz6258MougM+LE2czYYCMRGAKRTIwq/o4m4
4PWJnocejb+HhfBSLZ+Su8qzqQQ0mrKqW+v3JwhZsTjdDCTnG3TZ3Ku4bcDho7UY
CXiOlmA3pmD1iy/e+L6aR6azBYUl+OSgXBfqVaw2vYSZutw3QdEbaD5vx6+i2SAR
4Dc9O6vcM7a/tMdJQmLw9EW8JYyNwFcyaPW2B266mMd4yNNon4iFOKmpPmVifZNI
D6e6i6DdaxYeRz5ek/8zT5sUohILFkbYFuMzqbwPdVUgOjty3U7KWdc9eVLWh1bp
mkxQTcs2tPvjUell1kOnm5ztTyJ/lsP1YGlINfLvRz8Kd22qGiH6anvUIVh1YK2S
AWPM5FR15hMeiL4rcLfhOAhEU15LJoXtbuaymSKQiIC2gT3vQ17o6rnoWvcBQu0I
QMeuP671FfHGEwFJ0Phr3oirXTRyTHa09rOJDl4/a1NDEkkO2vZ5TE2tK6lXGDZB
5elzqNF7/TfQT5MpJ+SQ6r+zEHS+t2nealqi5K8iamj0XFXJVFIBewKYQG0qpJmm
hRkOy8sha/QiFUhxFRr7nzsErI2dDQS39MJHCtdk/2mR2wRnd8ZcsooKurHFU7Xm
hXy97e9qYyJvAOuH6LJ/M3ONfoU8Uu6Of0qMqGC3IaUUa14DlL95Dmbh03CDDDl9
WOzqv7AxBgTx7M0mt0l8h6zufO76S+PadG+ihp+mLtPKKGxEXryS/ugOXs0oTa34
Pqdv5Cjwq47dWZkWb9QKZYQVWeDqeJ1p1yGAEGN1vFp7LH74eCiPuC8vWN3MGRqb
JaGiqvVts83ybh1nWGIuXyjohg7qfc0qisWOTO8awSCaqmZf2CjlKU0a7nBpWP7e
2DlByS/dgOYypbdmrdAj842Nn7icKtDVLieO3NoyMCBz1+dRtooAHF6+t5nEZA15
kDqWUOl/3XDF1Xzfv1OnEDG8rh0GcuYRUeLzUit5CBXXrTrG9NX6K1XpxYMIYb/1
th9evxNuRinXB6rS63TfvTZUl87ENSJc+XKyTIvrmnUIy9cAZjbpngpAYlbYpbdm
IxhgKXjuZZoCcLMfhNMStJwwIRjW6uS2AnIx2mUN+1DZgh3ue81Ku190lD32PC+a
mPLprcMtlJkejSkj2z7ssfDS4tvwsEjAMH06o4vejoqF4uti4uae2vkjjkVMiuj2
Os5HyrvXCKHnnxSVzGr5zeDjcdEBaYcRjwS21BXX3wcBRDSMDMTUwM8+wBHL/Cj2
NLtlg1ieHrpyKeN9/AyPtBhY0iYdrlVyPK2ivqsitgKIDrIz0wZdhAtRLzDsoAsW
BCX78TF26qZZDepcBYEzV5uxxkLkpTqeYLxF3DSAcZLy0mx80IIfMDEvD4Cs4GNG
f7aOjyUt0DFipEkuEA/opOWcgKz00xX/SiKtLjefEKMCQJJF9AcIcNQQzkRWn5rT
H1ED3jZEE5gTAEvA0aaTayRuXYDFODcn5/lCBDA6P8EKBHWSzaZZPCMj3LRvNCXu
k7r48z+RPteLzPjrXUfh0WWDdsXd9BSZccaN0JYDmShtI7RFn2JieYFPetFugtXc
h630/f6mAwit8UYxZ26ZWVW5qzfl+JaTUdRkhiAQpp2jXnkaTxqxhbrLB7cjjN99
wSOFzXceKOGDPPankx4iXUjfyJ7o/j0ZgLbKm2Tm5egqU8vdujDiXTL83A9Q8t51
0vxjsSkVadR5/N0txdGYhOUdWmn8yzROv7lWEWBj63+i90t55ztNJXxStXvZ1SKk
Bzflqj7cf0jArBC+7Xk6MQfXqQxpOMz86risGQ41h8bGYacB0dQvFvV02u7qnqvC
mDnwT4IdcaWgN0qsz+O0Azdez3uFVJivkQd43WwKoIN8AlCQwh5fUu7rQtzsP8vG
MgYKHCI+iMo7AyuS+PH07KCI60Ax3SrPuP1ZHr3gnshjBZNDIm+O196Owua2wR1W
Tx+WnLs3bbqjgzyXnrV2hKJ0U0lhXG2ypDN/sdbDJt/J13q/gNWMZVvoWWgLuZp0
yfFsZfrL8U/mqaKaFTgdhvzMa11IwR6aaNh3TKEdlZcfCER0M7dpDTJPGUNq5V3d
UeBTQnMt/aLfhcO1OX29eIyraRV7uPB6axLE2X65TDIL+PRtKEDG8KWCEf6NGPju
OfgaGbfMdE7lNq1es4CvMJY9U3F/4hHcWvYFDONvzwSslAoLiVFUj1bkRmfFLN/z
lanYknBWiWcfizAWvc6kXcIhaNSEEggkk5hZqJ/q/1ZI7Jg5wiXgrVEycjqlU6Od
/okOUsnEyBSYEj3dnPD83I5CCMyNcKwD+39Dp+sqHmrhWvRWjtRy5q/Apv7JPter
9hLt0NnpnZJh5M67w9kYl28UdD++8yiBQepo8rU9roJ5uXmLLpVBAP886UqmeEiW
PJer3brJdY/lIyqG5nMhM7ZOmjmr8lbffIncm7a/bFsJozAobcSu7MxdjjnsZmpI
X8zFvWQizf1a7ahmCGNTBci/1nuAhYxf9qm0+D+Gsn8ZMhTF7P2Gitc7Sb+O5fjv
lyhV+v/t6rSSxFaWTn0sim7uvXw8Sk+0X04LAct1aQjXi2fGf1+hRpiZ1/srgiYb
BKFNmp2IJzOKGm9Kg4HMUnPT7BwrtDZQpdRoQA9e2wCnqnpAfdtQOYzam4V2o3Ud
vzMItQdvcAsi9KfZkwk7kuQ5f7HezWY/CUTrlaX8q5MRFETZ0/9jGEaIi0H6Kkvn
ji/s6Whr+zw2nc0l84t/c6Zyjj+zTxOqkoXGItNHHP/cgwz+uCHpd4tXR559enAT
lqNT7jpY+3HHxMRIw5eCoGN0d6Ogv+I5VF8MVdP4FrZoTPr1KJBMVobDADFDm7bU
FuN8Az80gCZc68IdZG/CZcR09j6J8358m1037vSvyUDN8eKqy1J1rjacDOC5Gk7H
wULulmvkNvB9k92tV9OGU/03SLeil3PerqPLxNZAswk6QZheHWBAEBqaTZsUqhQd
iNBpHgYAwf1vogjyGGXdNKntp2ZCoaaD9BGdvNKvXTORv32sbpi4c4Air6B8jIt2
HGjkJkTx/HdtqPrFOQ36z3Ex/jpjCOuYgebSnjGASIGMMFVPMXwvbepw2LuGPZPz
sOScW8YWiAftvTn9aoEuEPyT5t/h9SvdS2i5qmqpwa+wmWI4rdwtWDk9TBUDhW22
QraqFtwRbNGQamnZ8+FmIEOn8oa5PCN0zHzKMSsKw0NXSWHimb68ig2cTPDypuV3
Q5J2AxPa+CnEhbZ1WbF6icHS2Bo5/a5NXoEqsOsneRR/yd++i7f+xTpYnXSdfepo
04lUv0TAIAExqPWDK8oB7ofyLUUuqpKeDO7t1SvNzRJxNYfOgh+o4m0CQqP4xADr
h8v9rPLzhf9CXMHy4lXDe/64t0zBeofhb4Q/5gMOT5Mqisd9PmtI3o7PfVe0gfKC
th4AcH0hlgwlxcwcO9v0kxPIwZVe56XHQIw1S6D0JFxfWEW2ywbGqPjkheGyort0
pgNFPcB1dBVMII1z4pBY5Xo5Ldjfuomi0nPOGEzB6LEHH7RIe/rqIOXXMN5iA2ds
8sRvMuATCQ9RXaorTVPS6lqo1rw0r0Gomijf0Xj3zAvNqT5hgKnVanKqY0deP0Zo
ZGbPmQfSFnGHvxXaVg0EQcXPsJj02wjTc1UD+lEGQuEmMfdWQji3fEsuanux2duI
Zdb/+QnGz9K20+/8Dm33HVtKFaK0+YHskkWkL4hxOOlY4pc7WDVLtUHhgiSeehCL
HbmFqykZY8r9gTkeaMKjjdSRdzgMS/Hb5/9F4uWHonCfcMBCsHXupjSYwSf96Yhf
3qCFPpWw21sMSb3P21NigXOSvVbgWqNVPndQVYmUs+7OM7m+g7se8eCCq3tsAgkd
gOPKsSQCEjWGEkNRbBKhfwclrdORzvn+WUQmeKUSTK5UV0g4oISGrid7KA48Dcja
y8HIW2aGa1PLAJnPRdCNsW3qzRnroRU2HOtGcouHLuyNfI2kw61DQWgR9suPTyMz
gzDZy93CN2DQW0dE4BrqhpXzCEUYt60Pnnw5sGSop+APnRDH1ZQEXYVn6cRsrKJq
EZ8hg0AfUgYqF4FsYPHOpYCQsh8gLnaXo9qA25TprUr41yitUZqx43RSATYhlbK+
a4rvnJQeVuaPAnAeYqUA/xPvZvDT0wFN1v2tV18j1jczHR3+vTQnUJvx/bLKtipW
jbwLHQIXlCxuTUtInzSRXIVa1InAy2NToMy87BV70evs9xnbo6vMyw7hdo3R3E/q
zFTNbQYmoqoYfCObZ8J2NQ5N3MnIm4/Bi78CMHg+SW4JlmXuYvDbHmIyt00AzW3L
FW19RmN6fm+JuOj6hRRy1WKQZHMLIYrVTsTy7yeUy0s/ym2PU/ubwwjhtN7IcKMD
JhuoeXe4AaFE2SWTqNFGkIEjtCh5LcpaW20mkMPsyrNPlz2ibquF3FwinUCokVH+
2fQ1F7kwDhhaHIWMZFPdVD4rvmcP2uAcJvwfXa4VZAXfS5X0WOrYyUcjdNki1Hz2
/rom9m+iRnBL/A+eZ1yVAKvH5BrPkHc/DygAFfSj1jxuvy4uv461vAY/itTM2xdt
yICDORLXQ6SIyflvkdgAnqsQMhPzHRN+YbWX4icJN2vpFZW5VJ+uioiW+rRYJ0fx
yxpivmam3D9fvmrwqwuU/ZfpCjOcYJwbIiZYx4EXe3kxg025haSa8BCgtQdhyK2r
jnMiIyJbSs/GD17S4HRPsK6VUvW8FcVgoe0774XlcOwSsPrPQHTbMVAsAg5+HsBW
i8CurHXBaxiHqCNUMZfVp+khlPSQpJAnkn2i/2tiCQfYq4jXA+nDnuMVht1DyxRS
kmZkHEym0l9HxLjK5stWQ8Rhgy0nFUim9U22CldsCtFGhN9bWK9nTQQERj8DkMBN
RH2SDO/wENuhcgeYIIjCLuu8ujvLa9BLpxW6uBFXoY8LDwjIGBY1937/9E8Bvkxr
n1UByLYNn2V2v69OMYyEvDfdaGyoy+C3R94a7doLQrjz9EyBbEgOsPvr+MCCXxAC
Tx++OzRDqaVEg2JLbDA/KCZg/IAaMWKdB0+JS9X8IZi+PlbRjLOKd2yCDrA3MCYd
CU1n1C5sNSiYFlMF+i38C5lcN/uPzN81GaMApres73i8mN4q2c4fYBy71W3+T+KF
kVVuVKbigP8Tupo0wu2t73QwJOJNIMkD4/cB4KtEDWaDVp2ios3xdjl6/yFc+94U
ibZJZEdf/yYCyY2nYyYfZtOEgBlOvMkkC7H1u7ajI6OVZkxaxNLKCi4ynk6Rc7jI
TmPASinfiEDnny1fx4eg4AiZpVCOwoci5WziY1qh47HACd2+lObRjre4+Wh3gW/V
cdW38VE3Sb+qUlwyji08w8/PiXxv9CNeNIU2jiPVlQCbqVpusuJggDCgEqZi7iTJ
ylQ06xxokUwu5G0cxoB4stS6PjIW/oQ6C01Bn36bNNKhuqXdnicOrpIiDAlZ/sS9
2spWbsvysSpunDLTGqmBIU69rfVWVz79TKy2i0qK/D4ne7hKgg0Fr5gJIL6jqy+H
WBWS0HpFzrzjIPxexMxEOQHHRbPoJgIGo7Aea6v8fcjcKvi+HnIZCPZGCECvUhbS
ipiunRK7jrHC8vAXcM57z3rFoTXpXSdn4ItnjEAji22ODuvusvrdlwqnGVII0h0p
KjfmQ/MIHVZhN4U0oI9woL4MNfFIOWbgCN424ziJa00E8rva5p7YRtjro5w2kJGa
eZPk8UP48CAoCHXpWunpasN7g3vP4CEPQpCNLq1+vVn1YXSmm2Wjn+D4OYkfmMm5
AQxP/wMZcR30BssWunpYu8ojPoxsoKXCxn+oAPHzWoIZpPtLvGH5TNlYBO5mHf1Y
ZertJQLcGRbROKnD6yDGGFs6jFjx2jU/SeSOrJ2ptjhqZrkgmkKzlwP7jp5tRR1Y
4h9EnRV0sJMBbFLlweMQawhOCgJFDo5bjf4yNETX8R5Et4+026c/TNYP8YRGJ2VD
SiW6KNix+mfdt+8c1vJ8kK6HG3E5+kMuF0O+4FjXxNxRjmMdFqysCZiCpucfqDWn
c5grfRUwsP/ghoaO6c077bglwFo3oLQrtUBKa0HupMVIqKUbNHQzw8LB3CytIqbr
o/PcHTc00ifQaS2I4dmPtdZXrh+Gg4I3G6oo5ttm8WmFeb9QmPejMms7MqfWXyX8
ZL8UjR2DXs5TBoLWpyVNZM8eMuzkLiJ7Laeg1u8J/3lf32/wcH279jBK0AJ3jJxX
7CtYpWjcmzikWyjDb0+tIWjv1JvXUCfUnB38ONbROoQkBCwm4Z+FxzGLc+q8zmBe
FU5hY7DZyQDR5o+KLIfhcBhXyLwXeRKipcc/QPRDsQ0+XpL1k79HagerWApvcbu/
zg+yhbjm/2d1j/cEXwFCRHUlmNXOahIQmwExbn3rd7Jmzc504QlEL+kSCnePE4L2
tF+Qmhbsn0pmT3rlLp89W6Bba2bHy9p+yusVGKvmJ34Y0wusvsYjroSmUtFTtobD
Ttw1qgFaESFZfkNocwvMyQxZ8svdqaPq14yg5JYx3GzR2Ba6JQAzNmu6+aS4KIhX
0pQzJ6G/qn51Dgu/90JkdyFS84DSu5ulTWWPL4llIwFXdcHqTwxmuFLLWK4V3CZD
hdQqe9nDXJcFm3Lhz3vfVENR2R1zIZOtGY+4Ai8LjiwaZJuGHR8G5sP+En2VCenm
TOr4KvLfTFPqlO7B+HJhFERyz0aCODAjA86ttcsDEPoq+dt2dnF5qrErqo2YPwqy
APE+7GzWVFLGcV55h+lKOcfEqkfUluoMS1FQQBFv9pRO5U5HYDlfpmgss3OeESQc
X6CvM/MGrqv6wI25Xx/e3+TSvAs57WM5UauTQMV97YPuaAMtYbt0Ff2xXJO4rnz/
/5iLLBxCYlvJVmHrJsFuBGvEkdKL9uohgrCER+5+P1TTcuT+vkq8NU2RPLB0uNA9
F/Dx9umMyTSw9qYtuHWNelbJEusq7EWcjuBC6rcm3xCV5X6J0IP2PlGSni7vZvca
PmzLmi8CohIJrTiun4NyrhSN/ydH6ZJ6STtDDUbYZkLKwYuaHhaml1n7sf+ZltWU
SzOMuchguwZASANUO5ISdt8s2rconUb04Jl73KlFObO19FPUbmA2aZMxhPWe7MbB
KeTWT5aohxGPzrMRsiMCfGZPWbBWQvJvrxzV6B//2pxhCVlPNXRKwe4ol7F84VkC
+LDmulbJpliSDm59jGbORmCpYCqy5DEpVfvjgln38MFA1+Qi2vG//o77jCvGFPM7
OOHbiX2TfEFPFzBTdyFsLgMz12whsqbV8fiMaiaym3ei23G8jb+NRhaHY/+B3x2B
fq2E2WEzTdVUgxOev6J4A6qkXpxbmGeWXuwYJKuhx3dlOjm1yn5H+b9zBKFOwc+6
132cog3MAThWCDLHf6KuhGaY5J694Pkzrpi/gylDjrPAIyVVmm03FKDmXOaMyb3D
y4C0XDuR3BOY6tOLbC/Mq5wtNx7Qdpe9+UFcBYfEf23UoCrqZ5XVv3M/pAqqh7an
ETJtVn4Wl3R7v07iaU8G6bqakGyl55jbWHGLKlAiEyxFX2hQxjUvXE8UXHBZTyvf
bBm1pmAyf6zJ3nDwc7irIYeQji+ukzY87pilQS221svYkVYCpblqrYh5BZixu4SJ
6Y5kQXBOaVIAqyOG0Hh4e49S/LoWM/Bc2+6MNXBitD0wOTHzxkD81I9qR/b42Vl1
kOGneVYnLxAnlqTQZ1a01hpApQxh9GuWbkVf4TvO+Qv+o+0AuY0QTqW6XSoWhr6r
A/ftkqqWmil4RJP+daYwRXJSR2xdBbH7jRzsn2K62E9YOZGFzj3ZdDwqOIzOpLcj
yF2VRt/LYioPdzDNgI2gIdJHuJBYX20IrswFlS1bpVxRvKyUzcr1t6VdKsASkL7L
rTJSMGmYdqfLIoG6ad6/idHsWZUPs//J4Db9Y/lXrKCrHLi1omBVpR00c8vW2C+X
ASKDTeB6pDk/ylDx0Vf2aQikpC8u4ZMx/WuWQX0JmwqUTjPxokVHISyKN2ni40fY
NexDFTXoA4IlXJl8WKV5HkPWNYSwUPUUo3BDRPY5N+/KN+MIB56H5CwaAmnMeFSb
BkNBcnerIn46BAkOsW6Tj5JROK3w+3+vTnVWKpXMsCl8WMKGdQmzIrx/7x3P8Rsw
OjHo3OcLKxNHZA0B5ZMToTvXChRx6eFMtm0nJWGFZ9FZBMaROZgvYcA/yEqUnmVc
hpy01uBnYnhWN9Jq5LSu794b+fRs0PQXI1Izox2MKv6TIf7+ChrGu56YqmT0ENZs
kgDnGc2HDgEAK3WD2Y7BTuqWnQ/dxoeWcNnGl6opwYmlY8RK6v50A0j0Ms/ye2iG
d7RboakSZjN1+LYKA8c6WqmOHycG4felX943Z8/akINRCiQfLd1WLrlpCL9sFCYR
Wr4Mop1kbKNg4NswNzOypOziRK2/cgw06AlnAozYtt8zZ42TPPD6Fd4Zi9dSK5VT
mfbBWHS6DeUpM5OpcfSYVrf5WSy4exUS0SDjfVoU/DxgcPnkypKObu+8vSUVMpRy
761+d2DA8GS4p9m+ZDU+cv5bEE5VdE6PvqenIFOaE1nciAQXwQLwL8KY3zlXTSwy
FTvSukEKkSy95TEZnSD6PpvRCod50iSCAsKUkwspzO4Wm7jbmqYn/1v/wJiaDw8X
oxKVpmeClNxyt8aTnSMrJ/drpKDizVsktyE3mAtbSrSPAKztwut58OEZ3Q7KaNS0
NFm0duEDu8hYJrBdazpo01lzamWJ+Mzs6kjJ0jdn6YsbQ51Wg/bIi8iWqdQU0WUH
k/OOZ5O3yUi288J04xRESeQRsJQaFDJmmsD//iXJVB+yUkbIc6POKJuRBQP+m+Jk
Rc/h3ogbnQIc5CyNP1zNlLX2PceunaUxoJYjB+f7So7RS0T0P5+ZmfXUY91tqsb3
CcW7AFijrbdvBgP4YmUvn2YiLjfa+6HYKLF6rgiIZ2EYv6hLcUCRI06+vb8MfjRf
8pWvaJDZd36koZCglBlItlPb+E4UtB/SsEsrujA/M+AOUXV+MT9bBpSHWiHA0O00
n+XTW/+lfXSD/gymJ9E68krwrGoQ/h1hcuwyfd8BiVuYNYaW7/1eWNbterDkfm2p
09r9RHEmyQFX5DP7VKLNf/HM0FIG/NLgr9jXLH6Y1PDaWLWdbYhSwbdHW4OBWNe0
kFwgbZgHBUA0STlNZv9fjgm1S1qpq9KjgR1oM3/neyEvoRtWe6m7suLobJmjCHso
k0oXNC29Aww9IkTZwWr700Lg8mrc/f0/+kyA9Sxi/vE55qoSCfa+2bzZ4kXanFpv
8SjCxPinVhe0AUj121PIYj117VzaJU1IO2HpZgwWS8kmno+U37BhNKvPMPu1VKb6
suyNuiToNNgSz0PfVpOwkx08cU771AcY3RENLeFNQuo7NuSzkcnx3VaTqxLJZGr/
8FVXBF6wLviFRCQhvVjpyqT9rMLRG4hR3FBDD+bxC7UH0A88DZ98K38S0+NqQZvB
vpWIGXC+aDDf2atfgnp9uJ+d8jPWqOmRugSVjf8ZBalrTm5E83qkUxFAHdq4m9+s
WWotQnwhsIwUirvRdFaoNMDl/EilSKmwRANfbdAO5GS2xSvaAN5zruR/VpEM0dwC
63rPrPkfpw/85fbXQH7O/IsHmKe+p9/nAuJEfuhTvi6TC6z3Qw5NdOJjY47TSQwp
W5mv7OkUcIn2Noun4HyYJ+UWa+R/Nu1o5LQDnw/Drz+LMsrgIxc2SxlxpRjwEDS4
/JqU1b0JD3UteVKFAe9We9bnXs4qo3/bilTD9x7sZT+Mt1En2Nl6gTsMadZep3Lo
wXlkl392fpeBAv7dCLiABdU4G2fAxKNhycd3IOrZPuPUTjaT0qEhZppQBsXMM7pv
JPH5X7ssueaqo0yU6zDWyKCKkJjNE/pi5nwpx1icyp+6x1tuVYn7wYSI4s0vMVoq
X4uIddDWHH77+8T+gjUz2OMV3Mss58hTz121aZXmA7KDbDtqfRTpJhLd4WV/KG4z
BjjdDJ4ZgovvS7QkqeSa1XGMMFVPfTrmyFdWiQ2JiisHns1HFbht1X9optBclGb4
Fv7GV8cb98zYi3H3IAB6Z9rSgLeJyFfSUFJpv2Bnnt09mV5WNmJyZEhEL8yL9asS
Ot0woBQmp9ADsS8V1J5d+uk7EBPadnPXqBaKtir/a6dppyumfDdF/OvTvmObTJ0m
uEu6IxkEtn1HqzIvrqk3oELhLnB6iMJTGqUAvEvREuwaw71DZhXRURJ4JBtSJuTB
nZDE7qUw5GFCbsqJwImg5pur6ll/QDFOrKd8tt5EcKQkP7JbCV3jtRqjju7CLMm+
Z7zZyPdKpT5You3UpfkcJzao7vTAetldwU8x4sVhTgGbccrafUsrnQ2+PiO1K5sZ
Q3o6hSNiyQ5ELiLLEsVAgQqZuJyRhqSyqszcq/Hi11fDbk0Bed0F+WbTLU82gTbs
42/3RWBdPGqIBUIBftrLY4q8fhI9/dx0goOgPFw5ZCcZCzLK44SMGe7QLt0EMOlk
1DajGXHAjAEVXJxh75cp70pWW35rmpd2ubchbLjxGIsXq/E0IyhulDI6JXX4ZBVn
FWvNZJ3BhmyOrlCJYRAGt9BkHpHdHFv5ANgenC6/4Bj5pXrLtAVuQeZz1AQ1HpbG
lqKiBT6qbDqTuccxDgIa2GU1qGCGWsc74i9uimOGF8jYsbn274hyBBHitIa217yV
AJ7yw8nFTqIZNmLk4CYIRaxkAVVUz+LXovmeMTPliOC9CdEYJdUOGg/VF94IKv37
sWbxmDInNfXdzP/kAUKIdmLRMgN/GtUdpSvw5/kWHvQ1N10X6O3qew8wv8rKrvcV
BURjcijpH2L1PJqgEo9hIzPJHT63Rs1FOZA1zKDb3DkyEA7G3f/TZ8z8fc5lhWbu
ldusqlKqXkQ4E+cMphZlgjybw7mTgB1sKgbiW4qh94omX5ezyP9PpFa6EBB+VsBQ
/aR2F8nobUABfwJgv40zLyKQ5Gd2ZwKSIcmVPJ5Kyn4AhtcZ3UQeLQrBDmIHueie
4kN541955EzyL5aMrQlmjB/NtBXEqGD3m9GY0OD0PZ3s0yE3qeURggIT4asQeRv7
b3wn2FzYvjFAEqPuHKyvo1A6p7upasBzJVFnq2eaDLt7+lfxRGD5ams4id4ru4U0
xbuHc/Y2BkycH3SlNrY3fibL8aAeEsdSdWqPC7mp2Hpes7uohYyZQmu2/SVvBu7f
TFC5KIf6cfpRj5wUQQv3mmJEypFik15KHqHf5kcrPcM14mQMtNn4HkzTyGov4tMD
1VXbHU4eJJcEn0FVexePKIQ0LQzH2q18sI4iShHpz9oXGDjenSPFl3/cqf+yEbt1
djN6DEQSbY5q1NH5t0yDD1hWa729DI0/DXfjENKi3WDEszPdaY/P7Oxy6x+SRVed
zBAsguORjdGhPUtVBHrewC3Hx4DcLQlmrX1bNy0Yyi947aO3+UA/p/W9I72K94wk
97yqRUdw/3wr4RsAGBNIdVT5u3+oaYoHaZZQQSW3HmKVat8iYWmu7dwxOcYqaG4W
8xD4R/OQprp+rUO9+e5qFyB58b0622Gp38ruCAZendYTQwwSppNuR+cm85qcfv4t
STKbGkVEoBefCkQYXsH5oBsKMIueoZi0Hne0gqZ3itil4pnpORFXUsUPBupGVLKN
4pXJUnpEi4LnaXXDIRLQ+19ABTRpSQ5T401odjdk8P4MA2yzuP4ju2P9c/A9hVDZ
U01WfzGtM2P3sY1/lVIHjp6IfmQkA0HwkDe96JdLVYi1IN/ZiNR4G1AuFwxnP0LS
ksn22zG/LBm9K0KS6aifHsTtJA2GDME6r22z2IQnuEcjyYCqaAEtoYE2h/7qoX4E
oXMHQCkgN4Tnz5On/Ktm30bt5EDdktgtZ/t87rG5AetlZqCVJzRbftukjTLEQ3XB
rrDNVmmOlGtKfziTam+e7LNFV8Z6T9tuAAn0Vt7/WxPfyXEX4GyVsEZiZbol2Dvh
5uwu8Mfyn/BlkhkPgvlzFwIrRXDlWi1QmgFUUnKyH3Ud3XwXS+04+3b+K8RYO2qy
OYXq7qWI0BAi5S3zp9dJRcL6+JLxmaS5Qu+WZshydUrn12zT6fRC6NyfqzVrobNU
5e+duHR2PJIyXyF1OhM4yik5580yW6S332qUy0Cn6yioU/R5/1LMQ4IN0LMM4j48
UjssjTubXv9DcpZPBm7AEloPmN3R6/hnwM+WD75zzuh/NIfvzlsDanodOly9GQP/
GXdpUz/KQ7bFx4KGYrzCsVJQB7Z7FhT1N3kb2JN2H8nG5ilE8jkN5LDKOdwehfwB
1w4iX1PGlhmGg1W298eQiXdL606vxQZzafvfN4V8aypY5rbLxtu8+QnXC/4zWSWT
zvh7IL3jfdsZsB+SV5y7Dt+xZH7hV1bYVxUHODrc+4dxRDb91kUoWVZP4FoerDFP
2nz6+980VHgW5ykQcHjZ1lF0hJFsDN66po2iidQlCumY6J6UBbAVMrZZdEp9AsI2
uN5VPMH4jfpJFmobE+WZaeGIGFXgHr9MC1mJn0Be3V5PyLMk8BW68j3gb4BE/Rnb
EZuc+sWAOzbZ4Unk9DQx/tcpfmE6lGZtCqlVLN4azqkYvYuyZHyPCzzIQsKN0gUN
4xziKGD6JIwjYyu1YmG9CMN8x86+XVfxp4Ea2lc0Lc8ma0h+ArHu1o2O4JBHyScv
RV9Kt/+IMjn/i47f70qxxvFostxm6QKwmZgU6VctObI22qW2Vzk2LcKqiF2So1tM
T3uHChOirjCj2s7YuzK3c0BaQLpenatvFzqKpW7HRFzkzbwm8J7MSW6daMF3y3g5
k6Y3EpqFXNsiFLmHVwarsfsqHbT5JSmini/eHqdGB4dniQgkHjZcVQLUDGprOYZ3
DCJrzoLlCUL5iLpDb2PJWxWCMH60iWvsdaHnucyoye80I+9XtBFdbTyqu8ybYwAB
cCg8+Oib6iNTpTS5IO6m01R9Ob7EU+MURJrUQlAy3byDWorAImmRMRlPhpuxd3G8
hA1wj+aKi9VSWED5fy51GNPbCcJcKvJqeam0cRUs1hLKMUbec484Rv5eCBQOh0E/
glLhmWtdYg/HyA3TlygV+/6tKe/9WaBm81QCfTUeR/ndNVyEESj6IDI1LOHGtmYz
8nuYGRhFrZMj+ErAeZ9/jceL6ReUFEc4SYBA4k18piOwj24d+O0lUJVYzsjrub6e
fLgFIaArzDUtOuiCKTmppsPPwYveC4UjmrWXAfR1bCvmIEvFm6zXL0uBxnsjQG+F
K3ajA53nseAe7cIV/hETI9Z9GQJsPWCr8SYkk3nrke6Zu5yqhOZ9danv8anHBp5q
5xSPlfPlQEnaha5J+RbNSzyrLVP1C+q2ktOwBLQh6Hz26AXC9pXcFzkPmdO6Qe+O
T/Plo40ejGJNQyVbaE17PpeD0C9uVRYlcBdkjD76AgEvd7EPAEeYIBjsnu70isTw
rSnEHVi6a4QK1khyjPEvc9xhHo4dra6Vl/C6cqTqJKGx2oKFHx54MkYvwaIpWSRi
pyQ/gix+B7hmhL9qZx88vLP/gRNUbgeTycqMhbwzqnUQ9bVDoO3DCxUn44S3uXCB
80gd3ZfsscLi2vmUhlTVSrak9Try6WoqEMvl3ARy9sn+ARajxGQGg2KQyuAbPVxc
FmTtE0cOljLDt1tBpnZZh65bZB7jdRjAzFOMQiYrt6penmxo6d01Wy1bAa5hUeUc
AXvdCkP9xcPo+JWx5nxm4eCI4WuWwU3yv2ojk3GvuQnZZ1PBFCjdob1L0PKg6B5O
KfYvaWFP6+61s2lPhNE2U+J5KhqtdRy7QvBoE6mAAkjZoCG1EBYeUsLjhWRlpA6A
7tYaKSkqVvvWnx7XkkkyY3bf3cjqQvk2Zbz6CbkE04w+hsyaP74TBj8AZEDR4/g6
Gy/36QHJZipMrE2ptkMLEc3m3flzvWf9hQ1uuGg+nmiehl0AywlRe+AStTswlYx7
5HuhLA0RSlJEf9WN0F8ST1zQthWscJZOAK028BHDXr0BpXgEad7F/Gm2ew+ZZsgk
SGJ7twoqwHajtQAJerV11n8vJLfhBuvOvv+2irKN9OUpwTtIgjx3+DoaeTjj3eAV
8LFqPepGz4ALY9Nl5hz8+aR7R50BD7Fd2AXQOZX/D/KW6ktTNiwlqqkG2VWC8djp
gq8br7luGgtEvPpblG5Ja+ndIYx0a/NRxwdQncoA8s+ZhCzrAGUhFHzxTjRGS7uM
6siA7k133figr7F7/zwegHMg+fqK+kLRCMcF3pZasoRxJ0wXRiL/K2afFquXBM3q
VaFMJHscORwpqCEaf7fZBfN1JYFhVpCD7P7Xm0jQW4mQQgPQrhgXD7601YUFJDmx
PwqvtV2zS8heGNoV7dfdbPgIODjOpELyetskCNnffVayHz3Pj6FrDzgbpJT1VWBe
QiPuV+FfpV2HswudUxjFGuX20Rnol+fo6owlwG3b8wZhG6++YBwXVO16AK1lFAbh
7712zbuj/RnvclBM+u9CH+fhGB1MQCwjnK80ZJ6J/0Qn9QMD2jlFoOF4H9ze2msM
rpmvk38YIWBN9sH5d8Sq/YN33iVsQzQad249rIhCRHlr674gxc98cScInK/PIluf
0lYTe7TW6Ss+R0pXwYyD4CO+05H3trVffq9+okXtMpv61mepgatD6t2srfWsITSL
DAg9u2mZrfAE0vkXKXlrAN1h0Et/Oohn6ScYSd9SH23AFEZ40tohiJsEB5dwoqCt
Bx0leNDcoph8gLzPww6rDGtd+whrk5jB6qtMzNmHhAHCFUjm6kGMmeZWQTtEXTft
8wsQdiK8yCR7iirdkBR6glXI0yYRIZ5hEJZ/douXEz+5aIz7ATBfarPAjZlVG2yC
cFD0aoZ2JobEFxlsZKCecIz5QraA7bCnCnemcfgsxSDnxmRrn4M8ew7BUgxqEcEW
lxP+MPPM1wEsUmpMqg+BONQTw5XhJaJWfq8Aq02KYAobsDq8wB9i8NB6aLrrZ7Gi
PGEDl+0OABG/85Me/Wfkv3qJL2PV7zvSgl9NNy+9VMUbJ5akVbuRqG3gVP7AtLR9
vjULJw2VP5LGbZvBh0P04gmMXGd+4JJQrnGD5VMnDR7tCBrejOZt8IvUnDezqblg
9mwFJJKtIQudiIi6iClrj0DwIPzfAmQmb2sTB5QOeiHci03dFlzVhq/VMyyTAi/9
/Y+J7Cs4uREmnWCivqKwaLdcAxXziBoOJ3N3j2beArnPpx5kbo5DMuh441F8q1uW
iAyVpuH1GnHstGt7NKs0XfiynM+B970WjWGQztS7yhnymzFhe5dFm4EhXgtIr0Ah
wUH+owImYdNwcLyqPZw5vSc0mEDEbK/PnAhtNY4PmSpQ4M615ovwVNvZ8aWHuRt2
5xz+rXN4Yv+8kJMjp5Qtly+yhWzEDsr8PzyE3D/xQh83GhWeqZ67hAZ/RsGqDECZ
lxX3hwW3eux0ybmOWVvySttgrs1hmkW61yq30gDhv8zbuBZ5AMSfDLBnUrBv1EXW
lIZjRkdilPzaKbp7oGDw8IRiaGhw+YWgviWbBj+++ghb7NCsdf4vVIFzkyU36j8X
ovt/MZgReSQCWpx7OCDjx/14ijG5IrIX9rC3wGRE5BalohoZnpvg3YUtyakRG7qk
Vx0iS+LXNIGer6aCgmUauH9SrXsTs5v5QnqJQ2S68h0/PRSnAgo602dxRrbcAs/J
UrlDIDRdhONonP1r9R4Qm5HZxp50KCxbO/IdcXI9tB7hpJ+3Y2ngRB45OPYaGu/G
uy1nToN1UAfgVeCmTBJDDPf24kjuIR6yd0lcnawy09eqxs0171sobwlOzu93Kphc
Gv+vZWwZN6QrNnu6oZiaM9uIr8MwEgQWsq3EhZZ9sOzqAXA7hDFKvcmjvvz515qz
VyCnQMHeOwxUj3Y/f0Bb9DGZQ0N7ZLsCzn+yWCG142sOZcJK1ShO1rrM3sJGZta7
SUAzp0hyHWnGRpsDPyGr1Gd5mQ5FsYyGNoT5GJBbGBpimuv304toFO/yhngF81VY
Dto7gb/MkQ1lvoDLo/QBRfRaqMHoHeNh2aR+x2F3GLpWwAu0mNLFIhlOqgGzBfu6
61Zuwg4FkQqX8LrIk7YtZR7K26Eq78laIZE3g+JcM/ky5cPX6D1nBDlPFKDP4iE+
erw266WhwcYZMyxovgR1wRilSBGQMOnAivGODj3Kd4laTjC+Jn2nW5IiSk8rY47V
pfDagguaeS9p70Q+7VoMRmbtnjtMvjLLmGtQI5jMGN+BrtKzICORIyPW8XdKxOFp
GTXZfihX5WY7If+qiqIiBpd14iAefdVHQ9voWILTxYY3yMxhUndOoJxgpLPTSdrp
Drm1KWuhVh+AcWGmb6wHh4JTF0bW4vwFsMxmneY1ov/ZmcMieFplkewDmhROe1/M
eJkKhLdFnWLvVWTVlavD3bhOYeqH7TyyJ4HE0hUWReMAkIliP0MunxMiVl81Ehub
VTNva+30/PkIJNRxsK1bsn9f+GZOaLozLCJj7RYXuUCPhj7lyuYsY3wH3ElP64Ge
QhABNNNjeW+DNleesBGnMfL8K0J5eltXb5AseEC+07Y95m/fO13ZlDg1ieaiaiDc
tYMBJD9p498jCYs842gG57O59uBgKdJfqcX7GMYyIQMQs3tg3OJlMWlzo3emH5BC
zuLOBJctL/IevVCMshPYmeylyG9E7RQb2m8/U//G6YkBWlYuKqzGsIxEtB/NTbrO
qBIflv0VRq7IJVIjuG576cW/S+DBVXpjmMbNG0urOE5ENrrNHV/y8R798dGraUuw
ZdNBDZPhyBSzNqtRk5+kBIzQ5O3pxsM++7dc/dQ5dkEh1BwEt/Qij+PaILrkRFns
L16RKpTXS9b76EUAC4s2ukASpXMwPCX0gbRr6hQwtbsL7fKgW1YqhD5XyV+Gtan8
0gkJzcRPjqIqc1i91dVbbGGWAoWMcokmIfpbQ0BPYvZacGUXUUBESAt/Bzor9h2l
ykkaGYk4hYjGvRgIXpDhqPHEdqI+TZvtYAa3SA/zyb7PwraVcq8fRHBnnKgY2HAx
9xZRrfFB+2Wy3inxivUvxCWLz9vj8GvK8zagAkYtqIF1xWI4T/utOQFB6HygUbcu
yVPKhQAi7jRoD9dJWcxjGTfkLRZzHEmu7PTQSDzFAwoaeJcPkEfoG/xJRz0huVWj
UYkadm9mgq3gga6nHnQy1N4mZqUje6qGnu/ZMqI46xoTIzYlmh25ab/EreoTKtTW
70hxHDmH/nZiQ1HuXVf4nGQZa2sO4dfSHWU/3j8k276OrEjS6H7WNUcj+3UhAU5s
3Xn25P+q6O1vADnfX7xHY3j43h55bWLGnn82MUlUSv+XeNzU6k726MfKnjWp0XrE
X0/58KNeiqbI+deIwtzpMx8/Suq0qqGdjFw/ScRh5vA5cauYlWTlaZ60Bhf6EaNW
A7fSjUM+jgT1xqbq6a4ywNynT0rkUIg7JxogevaEoFe/QMPxI5iSPpmXFHYWJm0E
8DJuo+m8aZfv1l85IDCtybDI3cNLHhejZN4DIMTznEuRfDCL6YShg2FKHzDnt7UA
0O8F9uT7ixssUKD/886C13XucXRfJVjTj+ozjP4EQwy9/7wZrFP17+0NmpQuLPuB
L9YHEEjXOJAyfR41TpBm5DzdGDDLuXciiVc6cBIhFvzy8yODX/KQdNzRRatF3Lv8
iyScMFqos58sVl0RCr74rFkos0/nd4vChXVBPbl7d3ijt09iW0b8qBRCUwxYMLkU
E7zvl2jepwS0LtBlBN3g+h/xywGLg73YyTG87akc0Gs5rLw2CKfZn8lT6r5Z1DCu
fX3EycZBddA8CDPMVzPl2eesrm2MgSpacHK2B7eem4qivxZ5VfJL5fAwahH4Za/C
XfcQ4HUC+gACXiUVrFeaK8do8LLLSbnWPtpVATjLC5bdUVH198Fe5Q8rA7wZ5cPm
J0afMr35dpq5uCpI9ayoggIT+bB/6EA1lJYAOU1m6P8TsI2G12w+bxo0reE6q8YS
oj5FzjZZdOfpZNyvLCy4TsAd4dhQMOMzIeWBxrtGatRCMfh+/F6ntoGP2EsNx/w6
vavL71HYCJ0BPZmmjLW44yDE6GoHjBDRhGbJ+j5DT8TPmQ7fdt7/iu4GSqfuX68B
i5r4Jiu8UMXIN83ZAhsdd9A+HmqiPlpRIS3F1XlqFZ8yF/T/+EjfOll5OJAkmLVM
cMBhU4xxEH8CgP9jmCXWUapzA9qgf1fVjvnUVswlcClzlV4/qqrNedTXtbqNL6nO
s/i/0WLpPLhFUaqY+uDNxmlIBhCQ/K4lqFbwvYoVJO9BgKzCH0M+oCWDg/YBr92z
TC5GaJ7upHZHgOIp/nCjIVPvJOBIUpLRxFuNcEXUozp59JAEQInLqwOKVxCGLZxI
YES7+WFlgcdUJUhiYuEzeEoNig58v3YPBVPf+bkE/OZy3Ia8h34w5qHFQkro7a1c
QbT1KR1ZBZHtyIuPPkkWWSsW1ZnOyrggKiPOiCTBgKSaOsUDAljjYTfRzccq3X+Q
8+wqWxA2Nr/k3rHM73RGkwCsjZfQ9HsGYTDIDSlXP4yfYnpF4Ld6XyioSldpgBAZ
RWuUoyZyzNwvBweQ9ymfx9eBEOBdCnzKxDZF41VZoqZyaN1kt83KfI6Xj2vqjtRW
qt6YCcswPVYTYH1JPvOzXhR1/u/pJEqi/RBboacOA30/375rGPVEHF6b9t11pnR/
mBMsT82wy2kn4sX81Eypkmdc1VdMjeFanLfTKQtGZ45L4nh8RKV6YegibQdg8RxU
KNZJq0sUL6HL0eigfKt6jLI+J8Hci5GUgWJ7fi2G8DMQDb9or7tWYx5dXm9ACj4j
Wm+9kBGitE4pvRi+ueqFTkssxg4UmpVaofMYvNLzWxB+Th7Ww+fWDqB/CLwWKifg
VLrgyqaQHuJmzTdHLE4o943P8sCevZal2VcYPzQ4ji8DugYemp4KrVAxMFMbTLKT
m9zHc6YqlMNnLLyyLIz3jnMMzMxEunGvGSivO4V5GCfRxAMVMELobYJKB7+fxyxL
2t4kjUlWgXrQOw+NKmVGt1bxi6AAeHkF9XePCe3JE6umOU3Axibo1miiOTvFjuUi
nE0LZlUNngspOWrDy9s6FGi10b79+7fv5fL4ReXGHXZWYciP0Jnd3mYgYAg36ggh
1v8+1PXn1jwHom+TaeRFsnabI++Ksb7V71uYdv7zwEsWZ5USIeCXTryPPHAHxzA0
4RmhzrcfHNp5HI1eXKpVsKdV0ScpzBKCMffPJi3yVtYkxXxWnTWiEmPMJGrQPr/a
bQ05qh0tu2TBp1jwpaEE7fHtjjekqbtX5Y00jZxigNH7vLOVFu4p2y4UG4vwP2o+
OqMEBUXd4tgR3u758tGkweGDp9KzO4vtArWIjxk07TiBKIy4jRv88j3PAG8cnxcF
svxFJGEwdI7ccYHijUs3xf39dUalT/rO9UdE1vfxs5EWihdONNYU36K5vg4RYGBU
aHtSeQMMaWshaUcXla2vjMBiGSyol7EzxciSo+kF2CL+3zpxH+EAFrPLx2QLuFfS
K9oOoR1es2iZXFBFv3fNr0KChqtvH0DkkfsjURVQiWZAnMnDafqSDVyIkp6tC3NS
Aigi9J/mradamXydUnxT5rQ+Pb1pICOqCpalweFsre/qOfaWx7Zs7Vld7IlBYCph
oD3G6uOn0WpM11fEIJ4rVfgQurtG/0p9KISGv6j37AK9DvLkaqvqL8cKyVagqAhQ
gy8qmc86PTRzGmSy6fOnzp9AOyR3NmtXFb1ngro2yZWbxPQIXPYQjIAAMids9gcA
gzZbSiUUuVaw84NaRS4t0qg7xJeP1cSmLfYVJiXbtUtL9+V/AxyWOf5kSSfLixOF
l/10VZXjCiyDpdWEGIBCm6QnaQZ+FNiO+A8ZbrTw+MJ8tJ6hIG+DakV2kfod2xyc
JxzD093ntZgCcqh2xKaDav20SIvMqnTdZcjLiRGtgAcSTsjui0X2O1vOygcxh+5b
4QJiOdY+pTB7qQwTr34RwHbi9uizMLd/V1a2tM6Aog79/Hi3l0JuMLuPe94PnDZW
KQYLeuMV5W8cb/TkAiZT6rqn74mOU29kewiAazIrWFT3sGbWhVRQVJYIu8aXD3KG
8VsAfvP1S10v3wRqTXJSdPPZ1JU3RLov+X/yF24pFZ9NZ2xQWoILoCrryTNavwPg
ETudqpR54z0JkdHGn7bcxRhP3kgNxwuo7IXRQKyp2cZiR5Vt6KtQNcrLalYy1ekW
EUnbyHyDjzcBV0IqJZ5jFtAfV/HVQPHu+eiDuzLwJEWbtOyY7CCaiUTHdTnRUrz1
qHPvIx0Z7/3kjxPWpxRDsZlkS3Vquza3314qbG7VBSqlhpiLpR55Ka9YCcs7XteB
i7FOiaPk1scQprpU9Cw+xjIIG1mFr6ti5gMreEonRgYzGyQIjNsReW5bgp/Kem6M
7izurnBQ0hx4T5iEc1kQErIqlnlkcyrC1z+yYrXFsWF3VhxJvj7vvL9NyPy4P93i
zGseHXcuApQZirCQLVGbSy8Y6M2M/IYTYFwgKGF4kNS2othEoM6Lz7Gw1ffV2GS8
Ch6wM1cslqBLAUIxtgIS7FEZ9Qx0lrFl8pNV3Fkzw30l52kbi3chZwbeBWoGwQE9
EEkWbLjtfd6basijpFwUcWSJS9a1hBDNHnWed0QmewKSONbir4vOMaZzJizCDs9w
M+FmDf5+R4yXsGRe+Ary45f6scW7VH5LnuosUi8l4va5OD8KfZyMzZpfagD2adVA
6jYOamSlQ3F7k4MYzBXSLdBhR5BFCmNuAaqp6c0wVeLmKGkNR9/BCxik99N8slfg
bfKkU56oO5APBjQ8MF6dVxwjwNxnz0nm9WSkNodJQ+cGV0XBr5sV0mZlikmYqb1G
zQCjLwqmY4UFzM8ddAG9KkK4rGTzD7wPSf5PylHRFm+XywnmymahJBxh207BiyF4
g+iZKrlxppnKEe41BoXfVd1ogjDx9fsXekp14ArM8GhG+37uhD/tcZbo36wUkJZR
9RWOqMR9x/Go1VH0k916pgERJj5IUb0C5b6b+E2/w37XA28eDf9mMBxTdg2An8aj
Ue6emtsqiehMaYZ2Cu1v07A29tlaFq8FGwM7zfyjrwu72XHZXW6/o6JBKUEK7sb2
hNvtGO4ZdHgQbHPWaXqnbBQK53KfyPn9CBZszOU/IyBgUx3aYvBb5yXX0edcqMu2
vYsOQ0p7udz19ce2O1biF5dOL1MGx7dY//Eolc2cXAA7t8oDbJTcvP0BGRbjhrbB
tcel2ikTurrGwiRk+rIFxuRl191n1O7uO17gYbNCP8p5f3k1P3tLkHymgriQidLe
GVknQSVwAH/664IBrx8X3MZHKI4Q5Q8/ZFuO4KAGq+YrOpQaW7jEgUF/W6h9N3W7
sejJ+Mm67KaHCw5HxGPq4x08yN0lNKiadOTCEa81iK4B8Z/NdaxP8wK5UbIDtNpv
H5v3hLvHQStlcRW3nbi7wk63Z6bKGQZW8TW1Nklxkg5IsAaVFPgrBAlklP9P7+HO
t3s1c9Vi+pVgYNrI9hfyywgWmBPDTGba/OfPm/DX+B7egd++rGLT971W9Ep8I0rJ
XhHwbJAJ7bN8b8Jd655ILDNfIUloNxlm8F3ja0h+zh2S7ev3R/lgTjhdF2Y3NWev
6MiD2GEnB20ELtF23/72JBYGLlSjftEjPVA+cQUq6StI+Ay2jn8bruB7CSO7q2Cu
XQNNHtrZEyFkSWxMGUSYbM9+6gMi5pkIvwTky+bkDbwlGXf1WqdW1Zc+jYi5v1zo
QozRWPQk/OhvMAE2n0EjkxX4NHQuMB/zGduSYVBxP9CEv/V8GMIfsqCSilFKtFwT
BqZ+PGxt36BboqvzwTOxPe5TiuR3SiJ7xqmD78gBFACNfts3IExFsP7TJ09vEBZ3
Go41yg0+xi7UQrkwfTmE5uMu2BNb0sjBszYO75jUm8bLWwh0DnljQTM/97rmtT+0
3pSsIkZcnUaj2DCcsRIOk64WjyEVcQS+ZDd3MPn5EFB8Ij6/XEd2FMZNhCiaODCW
US7xe/Hv+crsdGWW0XMfNdpzPifJmVfNOjgKL9XCB0zRvzbYOWtcNaq/TPgDHKYJ
1UKM2LNdl1lIcWhJX0czyJzmca7uNxlpMZAE8rYg1H+HtpIPKTrzdH0VJuNLLqU2
ua+oXxVcIq5wMN98qI+eUMCp6vUXlUXYOk0PustIOKO+9stdNLo5Hr1lxz1Byl8Z
Et3V/OHH3dGXhLt8cXbrr8vJRApJBOa3tIkJDySiNEB7Kjl5Ie6ZSJDL/TkXMTQP
/l7kYPV7DGiuzc/mZ3CZlhChnbuVAvAOvgCmDO44D3WIoE/z6FDqqw0jjgo4vWcc
Ul0NwxA0C9sKymsZW00M9SQ1nYcMVMn1h/wsGx/GMXcF581RhqzV/WdqkuaOzkn3
O4pCbirngZP8SQUOLnd4gEFqx/fOfxnmYasfpkNnPh8dg5y9xk/poc02DFyvoE4X
4wqOlbUvVCfHMoJC5cCu97fzynVXVSD+bmbqeNGxnGSQW2kuN6gSd30Q1Y3LrcoG
xwFkjrm8/W1mKJ/LWsmrtKF4HZLkPFW++CBOQcmpE9U8H2l9HIRjk5En5B5AZbPg
+6tJ15imS2wkY1gDHNE1BXLwoc9uH1EcCErEwq0sR0H1QIM4zv+zE7Vh+L728RlC
6cJJNR8W3ce0pjZd2tQ6ejw/ydH2GhDNSpGXMIBgCNCh32f2y32oWJ2iqQFB7+c4
y35+2NaRfBSL7C3g9Xr/L2sLqT/8M6j+V9mnoGxKHjD8gfohVaYInoro89ISVfFf
8WF4JVL0AI9mZljH21LNkq8bzUZFR3lbu0FlH0gGCeynh3RbsHCG0LjANkTuaJ7N
PDMsNfBDyjTgP8dYtPPDcGg2G1T1Ychn2SYyQnaxsebWtOkM911DUI1d7TyOGIO1
eUWFIzslZ5ZsazqITWyvl+SX5v0/DK/umizClMievYMhC+J+NPJ28t86jbZcjNJL
/M1eCPkMmF/vLUuiPTISGYtW3BXCmxnLKjVKswpZeu0Zdl2A+RucA1rt0JEMEvN8
6aOnmoe1SlnJpyqej5tQu7oGox0hwDmo8QQAMbXCxQQ/lW6/KPTAdPOr26WBCdfj
5jLA6R1hzdszV1y5XzBx5zVLKO2IbpKWx8P/medxYO7wNShwVEWCbcTgkJzuMx7R
C3dkpAIhN0xTh52OFEEhejQfJs+T+IDZiuQjagA025ZCtgdqXOrTs4Mmzm50pnbT
3AA+jvfTSY/Y+kms6KOPs6Jhp0HVFaOeQ2EY16GKmccqhXQTiRtuxcp0XgMep7JY
0IK91xLc0yE3vyJxRR/bjd/0nC4K6ntMu0DjA+3D6epR6hl3Ghd0dM6r6oKSIri6
aCL7eZ9Ld8QYZy2XFxTmqej+qFl3oH0Qiz23Uwi6Vm2YBs572w6+T+VL7C+FLqba
33GciAIc2aKsfYKfj1+1riCZAm3OUMD6BRNPaVWGxNNOFMhv5y9nyFTW1gjdya5q
lPNWYzHnZKizv70ywqBbdFSo5AM/3j6MBdaCs08YQ6qrtYCTFGdhnRtdxLOb06w4
3wUZR3Xq93P0GIl1amqJs4gE/DUuE7lzETkGH0P9sy+Ggc4qfEb3GVSCpRVdMD3P
JS6ucbTG7E6NmHUWO9psW+Qgf5NBs7u3YKOW8cBLo8FXAE1arK3sYB94IqcvtMn7
ccWjtEfZ4CId6Hd9lu2F9J3wxE6C/1/6ovfyphiM/XS0NIQjyiG+oglDQ+TlHSdt
My0Izw+AlY0MfSfaX1d0r3sjpEk/v6W9Q40UyYYt5wBqOT5XsBl3P3Q+ylLf8AjS
JW8z6RDmNYZsGVs1+ieqjUll1J8wnunCFbWZ+JOfHNDMNHx6Lh14O8krNWQ1OZJF
prKcWZK6SKkkkQl9NrZc2rNZc8MPcBGYtYoY7R4V8CduC1dUX9/GOba576wYX/+A
oOHfJqlXJjkfwKc1CuKWBVVLIHVgoKmbItQhHKg5ZX/IxEXTa+mXKjZ8QrYNs+5h
Hl0YNC6USW/ivij9p16z7wc2JydBxKSgcxrN3HPQ5ggy3i3UIFJlBI0HX+EAZQUR
XaXLna+J6U2Lrpd88oUDnUMQ8U1wfizDOrCf/JlaHFrlZv0tSHJJ+c5NM4N/FHW8
oYfMOHWIqE9sW6ospt278vhJdgMY1CbZDGR5Y4ExV50iyI1ce2FET0CQdqLH5LvK
20gFhXJhrUe654wlwMKYBNbeSDSmva/xcJu6bfYulEzrrQnC+ZCmRK4nuKyfkiKX
dWPlqSlfyfyAWmagAluZ8UgZXSNxMB/bdPxZxUfZ1bCj8WuxcPF1alUhwZ2i+WlF
14IE2AFjgGUTUPKQSsZJUeedIuf1LrL7+nWUiy4KGDQBY2g9IA7Hm+4XfhnePcku
M0qDPMSx0LLkLLGg3QBmijaBlvsYzdr/LOtUAwOFU5Ur54liWLgCv9Twzso5mbxg
Une7PTdpPzZb7RrlrxJ/FE01N4TTaToid8Fk+E8WZbDp/famIgZ20w3bSof6tz4P
KbYb5Sm2FEoNZpbM/fSlz5+/HbrqSOX2lupqlnfiQOZpfQgNEYf1/UyzAXvarqSK
USgcA4bBwN+cC3LoCV1vsCqQ0tDIIUPyVhJ8O0ZTbQkiwFikSZ6FHAxwVvRrRAWD
v1SX+9twP2/4/532Qx8qOniThDbyWRNgjhMq0xkf8XAUCXpZgeKrPy6NMcwvU4R1
PahmEzTJv+XNvDkZSH1Mu9E4G7vsL67H3hAIJ1bk2tRowu2CSOYorkWUacHQj72m
/QWmduN2VlI5w0Zrnp+uwxLWGHay/5ADi1T+GJGgPUYEGkx2obXH1TXgheynrjFq
t2z3C2uG5cz/Oe9Mx0LLblu2E5TgwVEg9ATmRWoRfAo2aHpSjAsVDdch4ofvk0u3
rqu2db5C9cZ/PhhA6NBewYvZXSyuCzUkjuqleLButDu/Bh/xF2cuJ4pW242z0vNU
0H8bvP/2Ucf8Ik+c26yIP9DlMTln85MCr4DJOflydcWRGiHfrHhpTCq4EbtGlTmG
2LLdOOoS7wMivpyPaf8wHzdaoY5eg+SLeWF2F3+k3GDYQUTWpFRCWvKNTXuldrhg
UZzVbb/eDrl4xLkvaoKUdTOCuHXbSRX7A6pITpS3gbJr8FUWr5IOHbbxeRzFeArW
5tQVI+5kIGOSWmWmXufLHkzsyGBwNLF2pCkAbNG0IxI5aXmUyy8+N3SkONmZlyVG
F32DfVq9+khB95xK/yNrJfLNivqFibQ/lTF/svPH8RUqBm5fHCPzbKE5WhaDOJyD
LNeriswgsX1i11LRLEr5vCaDTFWWbkr94enw22S2zvlmMu5Kbmtvjj2KF5J1eosb
WOCh2SWR9/pQ6bDvHiNQUu82xjVaoG68FFsd9k3Mcgrbn1HbkdN5A5JZRSYfcI8r
8/XEQQEBC+7GCxrhzwrW3BRXUwKrT6QJRCNL5syxdTi3poRJtfwDFrS4HA5OLOQC
d77oLda0wc0X77avdFBFNzZcYCWcXnwPQqLm0jOFaE1RBhHZD8DwXcpwaEWSPuY3
FwVx5c41CNUKtA8dajBD0UpifYAX5Ogrew98jemUT4yWwPSLkTFTN3kkCoijk9yO
Btxt4+P8Prg1ayOchdTXmd4mEy39tnANZuEU15cbR/BZANMWumG7x8xOgEjYSgUU
FApN3K6HWPCUKhmOIG+4uxaLaKt5lyAAyK3d0Q9HOlIf7oo/kldB46HC497Ir1Jo
FpqBuqHoKMqLPzG/b7W3fMi7/KsnmDS46he2wilNpKN6zHlyxF3ASatEfHzDKpc1
oO3+XNVny9/HhSGR2h7EMdo8HRvM7jqsQ5IuaH3xh5K2GHrvLnPpdfXPw1oynUuO
05pyrg6muDWAubCHFQ6imWh9sjly21GCcqHatc9HzM7Vy4d6CzcKYfgXGLtAYOWh
zAaXdmW0AWJY0svTQ7dXgbB389P37jxficVyNtG/NbxMVHDMs86idLMfVK3IGwnv
kCTkwAaA+PpBk3siHpuodP5grWd5Oyj50EObUoJVtbxvg+qYPE4zUAGBoeY68QYB
8Lmuv1fiqMczKoE6BTYvjKTiHcMsGTy/8Ryb8yKopzvAc8ral2XvJaHXTk0qrvb8
lafBczSLYgS1hp73pnKu2zmeDivZlYuPA+z/YZ0Y3Ou0/A52NqkYjLd+q5GuSmje
j7n6nRV7Lli2low9h8DB7qvud+1iI7rFNjq39Dz5atoaytsF7AAnAs2hXbVhnWxn
rAo2aayKLjdnB3NP9+Atx0CpO0SzyYGxPb71n/lwpETLjaekmsMa/fXK1hTDz+fk
FWLZQrOuWg+ecY+VEVMC6nsLQbTaa7M8fh7aLiGfXq+VSzKF3wFr36A3TLi0m/wR
o/4v+3wnEF6XL9yblWICKkyY0bOjsOu/29dqikU7j1NDWwkX93NIZ+9wOKjcs+/0
10rXWGY0PDIeN37lyIG603KeqpS/u8hh+uB+C+klWYgmVR8cIACEE1YTmm1tW22C
rGKviHAwa9tSHSIwnicgjaCpW+OQlY9QIdHssD39hEe1B+beA5Ahh8YY05udRMXd
8yhsflcwpgwit5wMOrSaiRwGh5PmzdcIC+SFXuTZD/WI2RLnWPXu4KBjAhWxq9z2
O0oqw3r2SPFMBTjw5eGHAM2C+8WWfO/sk3kP1sER0s5G+j64DfFxKRrzMgCrelg3
zD04xi639NdIuNpst/2cMIcJBgsLLjVvwmfRxKfebkCzDSkL6wDSnEWO3LldGSXG
l8PdkMSTn75fA1CCQWtTycMisXba3xdDcmNAOFo4s65fMbtKbsawcf2ovry8zo6c
EeyMg3cP2v8WfVE278/Dt7MZgeY9GMPYudtZZIkIkoVbUcG36RWogEp6W3S2tCY8
1rHCIblDJaO+Tgzi3Abrcy42IIaOAMJQ1nXbGxrKWdHqBUU2cz+8SgzeD2XPSpXf
DOSf9XcrZlKyMLgSGuRCp1Hu8zwaAYWJn5t5VWROELMPqC0ZEiHduCoiislfQ7xq
Seux/rXVC5fFNMZg6nCdj8WpTmi5gCe6qN2Ylv1H56NwNdDaq+DaJhYfNN2zcQ1V
Y/5yXSg6KbYo1hwdDTMO2RvPkCrlO+3aY9qFkNGFO93R83TvgkOl5o3elbLcjCTH
mnOb2n86kqMErP5M2S1mvCqetHVAcOFRooOk2QM5SwOxlbFKLWl8QXqgNd96ggGU
mgBA5VQlTXQNt1/DJY+37+M2nkNoLFE0Sn551/iqYgIeucllXcNOCtm1KHD68YIx
CM+JOZZlG1g1sCRBLyFCP+VyFQMPFT6XIIPBrBKC4mSnt7MVV+0P6HbP8qHXzd0Q
MQ3bDWyXvi1NNHJ0mIWhXJMX5e/pzQXy3hR9h4VlI+VpscXvi6MG0fXjj4DN9WE3
7dGm6Z+eYZWFNecYQbxRKUlwECymVR6Iuwwh+m6EkEBwSpL+6vy9KM5zlVnhdgTo
ua941brqEKB3If43YnG4M5QUnVPtl5MyvdoUMAESvohg000PgL387HYF0Lu6gjH/
BMDr3Pe/+HOOKdM7n43C+EyGyMo2vVrvpK5dpYefJaMBko3FCmNM4q9YVjjZ0gLC
98FpDi0miN/7u3FppQv7vxLPaRugefk0b+CraLu6EszOHK7QewPBFcpkgvlRgJf0
9OtbC6H7t8F20rRcTmPWqFYvbWnLsbkDadi7EQ0Yf9xsiFEeYyjpnJe3wugyCI+n
jjvWaHM3gsi69BtWeY7g2HKxvTtmyGseeFqdW/TFFVcMTKKugnhy7d9yV0Txy2p2
Tu4ufK/1orkNmBY5xrhKqoSFRy0f0fzpcVH55uQnNio32FeAvn9VhCrWeOnVJBNP
87IW0atFQzF9OMfedvaXtTLGe0bQ91wn8lrI6ujOICB3V3MGyqeQN09onPyrI9qw
9zPbMoZb73tF6jcoNcAYoYdKRmJAQA0OZlJF9gPpF+d7bdznjwOMQhoHYLQeCJBk
wg/oH724jtl3ccFWhSa4IIFwUGdCeioimu0oJc1DpK/M1iDY2JtaeE1ILSQCI1mj
XGLpXVLplq43cTyknlfazABjp2frOzpfR3PdVkURNY5UTtPj/mcr8OAu7QPW7NAs
yPvpX7CQo3GCJj9sSB2D2XQuFMfOKSw6l3r4h6S0f3UnRwtv1CSt3AoIpYF/eJ6O
v0W1hvSKWcsC5eL5GPGSNVOx697HJwqJ8z88lgO6+hoIHdyJFtBP4/aCZwfRjOHy
jtMVZHxByb01NCmGPkqvyowzl2eUZv+3uNdD7+2Ir7SHTFejrnUd1+mYZsUzQT00
Y2+lz2pipCNfKF264SEdQnHd3L5lldXIxb4vJ7p+LkgJ2KqaTxy9oa46ARE2x65/
sIGvgrQf416nttnyC72iURam6GfYXrjmpchhN9GQ2HokpEzfDnjonNfk4BcZ2UQr
Zl41ebdwLIyRsc2SH9yoCqCC+iuGWRBgs7OqxaLxC7oEqt4abWpN9TWjUyK89ctX
6LJzcf40665vF+lMu5hlUG87Lexuc7swmxGLJviBbYmdkWUfCJ0zZigabUyEVW7m
uXxJCZP8vTszLEGjWagNMKJ0iBcTLIEhTcYsTcyOttugvqzFtpLuuNuv+w9tvk+m
E+pSL1i5W11r3cdokv2yTk/dv5Pye4Jzc9ePylCZ+Sg1vvhRcUJwVR3t/d38a2IC
HTxa0calcZptchhgDtuOuSL6+9/H3K6kW5KWo789hNyptUM0VSIhy6ppzgkECTPE
tmTGBKM+QrJ5bv8jJ6l8uyluFtGhW1FDXSSFJ2VWMUJqlMv8g5G5zaqutJTLXwFa
4WsxdCo/v5xeGi32N6MklxzMXQ5kAJQX84p+sVFsn7M0UT6rmOETSbJBj/C3XJX0
JYkYWjSKzkV3pbpwBytEDqt9LJvUrLhAdl6oM0fiFauETRQg/CdjZAFD/m1bqGp2
z836tcgjVFTCA8vmFCDfB+tBNh+ki/klSh8xuOmN0g5x7wRPF5glD365E3VjMHwC
94DdaSE+mGsdI7Ekq3b86A+BdTJ2xAXhSsHMkPJ+VniYlf1sTW1oSlCFyubpOgxg
I8+40CviFXhSt2fg8RYMB5y/q3shEzXR2pdh/6BpDkusw0UCJDjrA3sD6E7pHNia
0/ly15WeswFRcNE+/Ls0AFrVTPdu5jDA/nYLFDfNQwfwcrk00GlvTntnSwyN9nE7
32ucoqP3E03s712sg8gVlHJPpqAhesIoUhnI/udSPhe+h6cgC6j08OQd8N7GjfLl
USqhVpcMhN6xgopNShj8FcaeL7nCL1v33jrrtLXYG1f3+hHC8pahccELQHjZLbgD
a7HwWPHEm6xnNp6jRXILXKnQr0EyL7uZ1uwJtha+CcF0mOcVZNr81DCDaev+Sp3b
Zl8uv1SM4i6J2dX0m4+nclehI5Ec5smC3AfTjyFK1KyYF3J+YyJijqK6ImWToPCC
y7qiBrftJX8d659KGOZSvhWzq0ZE1quqRGwTRwSMmyFveQXMhQkKikTW0Oh5D/hw
5S9hCtUz9EVkcGd6/+r8f82Zz2L+t/Z8O2Rh19jc+ccbAEbZ/Wc42GHPAdT5xTiH
CpmzzJiQ79Stvl6IZKl595VrzHwcKo/jf2XtTmKdv8JvefqBoLkgmcV9A3NchqKe
rsLDZML2CuEy8Aa1KC1keba1t09lD3JwyD5OG8FWQWot7eTWiLk4OHE0uOgJ83CL
epPbExTO6mfBwe31o7RM3S2HJcFPIPvpxLCjNVc9eY2pyJj0qaAAPDf7+9R9HywY
2/u1vxacshry811ZaRP2CVXQ738AfcMX2nT61tcFUOFx/Lj0L4Uc/hwJiky2IoWj
m1XQ7LAe5f85aKFvikhGnd5JD0KIKcTcYoUaWZ4jG8RCYBURV7VgzfjDw5fsuCHI
MVorEfW5R9BlBIE7PTDjQV+r8nVDTRSxBxQzj6F7oj4C5t9tF9Xg00zDmVM2J/Dd
kG5D4ye4WqxZuXnVfQrXdMs9jSkxKUpBYNeysTJHYX2AAZo3JNQ723zSci4EYKJ1
4A5OLZ75Qjk1OkGXzGHwaZE4nRVZeAVk3gaSUXSUzEuTdivqhslt19cugvATKSqv
ryO+DyffR7iehKDKt5tkg7FQ9IiFxUN1mUwtzfl1N0G5kyBJ8rBHhdkilEVit//k
faXAqu8Jz8tqs9CRveE1hKl08nodxE/uVMtb4wfdkuDwQIIazaiqt5Ee4RFphY/V
fYN+zZH/1ZOqdojwF3RubLwb2zKhyUs5fck2uQ1qaqf+fB+H1BLfYS31WVVEDepB
FHEmPVxQ4rWKqQwYcDwelVLXM61cQCJVALFw0eUifWK8UJpcPymn5oav6KuF1GfI
AKjxV7KucViq3FeBapSN+eOhkWJxFg2BYM8UD6EN4jztEVGsmePlHvvb8YeGUUfy
3DF03ustg08wIlabIGb+hscOTFoDd/EJedhRLjF0Vy8l+5+wsT3fsLJpTSwI/1bA
c8ofMLtNd39D0AjeU6AtBoiEh5TMDSKuZjAc9oKvouCCxNrNDTSShibv2obV0nbH
xgVWk6ztPNJ4u6DZrses5AhW9jvBg38a7OARNfA2GTHfyyNOdGXUbQbZ4Fxf7nlB
m1iZKH9PleXAKcGvlX5psvpATEwXLt2wpu9HEbeeczbJ+hLTDuw3STlz+mwzKeSP
3gKkqJZPWGELrqXSC+kZ5Kdl9/iGvHeze11CLY0ccTBxa0sY3UhjydOLDkSdMwhd
b2yJlh8Q/4bQIIrsNfQ00BYbeIj95EYuH4iU2DYh2YhA5TnUyLGS+PlKyf4U3fc+
NYeizV8MFZXuFjZOTiRdFjYxLSIQK+O/PG0wsMVNTT39b9fo7g80nyJKcgucFNcA
i7Q4xYVke4F1U+ORVvLummZPTwhllWdtP202O8OlHCQFkCPXkZ0uxu0Ci/HYyBLk
PMmN6Z9RkCPLFInFm2m4UXwIaiclwgkTu6kG7e830uMmkzhqU3yBdW4ariTjE5Ll
debLKk2tBlycN3mL07e9CnxGsaZIijYy+TQUwqHmNPY9FpTpLF3GYfOlDXIfha9i
GX6IPeagRtGOdbMAYwRS7xWX19c1dEgz7FSDltWy5lmqcy/3Gatoijt+wlt+uXmP
yez5ztdatChA5XWou3D3nrQotNyMbY4SA/hs8MLyP8C26K/I6qPz6p7a3U9v2pTT
mIFfaolyfjAWuBcZAW8Tb6mWgEwF7sfwY1GbEBMlNTlwoPVhDpmvn9IFh11nODeR
BBDE2u/CxhrmbQLiyCkVypWf82njjPa7kpjQWPkwnzsJu7g0dVrGyT3JU3PY3xj8
N2U8Ytq3arz8Lz2BPaQZ+3M8sFiLuzoJH/C1AFH9V6Yzlj+95/QY67GBX3Ss7fu0
Ap3kEiBCU6maJeGqZhuoK/C5adrz4KDKqW6FUQW6rL6A85TkMShvqaPEKK/P3tmV
NYtYhIGnI1ULmhbXX7xmc9E5MOFd5ckb6NR/5/uqZQVdTM+9I3i9RnyYWS2gj0hg
zAPyQ/t6rZJFg6pX8XjfwzrHiuCbL3SU+nG/a6dnZJZbtM8gKNCppXAg05fycCwD
Q2L//5mC7M0XYRUg1V9ycZy1oS+H5vcBTJiOf0bAk/QE3o2D9SqYfYBnM4UZVKF3
HAeX1jgDvEfa4aq0qVcjYwpkzZGsyJ6Ll6m1Csbdw6dFpT74UBtlC9r08i89xMUd
ls7/WFNJsmwgXll0QeV6+GYR0NOSmcFjAJdlkjvCdfsNeAD5aYdqT7bTjfgyy52V
ttNxyp4iKwkmkaG5OKcn0hQsiAiVe9bbuoOcsWIvAb86I+hvA9qHPIuK3SfxB1W1
K/yfQBEf8njvc2odxH2EsaQN0D4xu3yrMDqUCyJ7OiH9crj05ZHOOpwrRN3Y6hnr
7iyEhnDg+w/1WDfb7AVYk3d/wufRaQWJQiLfMf9Vlz0W28/6bUoGHrJuyZVsA8uy
mAAb3k2ZFTsqh9VOIG7QX9DIzUcFtiojSSsnLnkFL1ICjaJtWbeYlpIje922WuOo
YcysOpXPnWOBep6mCqbeiX2fPzbrmvWDxB8Vdyl66hxm05b4GdYR7pSJkOjiuxw0
kUjOKhbAqX1PJzRCuAgNrVcY2UsVPf0EJPVurQNcsgKj0tM9/WgmSQM1P71y/k/W
lPCVdu60eQ4X2aSOAePBmcHEh5wRVcBbuxrVuzHN1OtsspIb3OBSZwYiIWVS5uvX
TEyfHaOspXPnZCIsw96s4fD50iwd/5zqPq+7qMg9//GvuhFvEK4Vh+Ze1IFts9r7
fV5Qiaqbb/gnyVQiA8FclWCiddfz/fMDV2p4VGwqt80nU7k2sbmFc72enU7FKaVP
A/8GoEqwmz15p3zR9UBlR8nSgFuSnK1nrC/B2PbwKYizrPpqBbA2xLn2d3JttmLH
sJZmWpqwSK4gQNfpHa7etYMSeQstaD0uvWrqlcWvA7by6hBbSuPIY6M77GCLeFCC
VH0iUZlUt2e/RZF+41yrvMELoLR9PzyjvlSTZ+tvFB4FXb//ye8AxWPp5aoCJd6j
CNwrX5o3YRM+Sed6L5DUXp3A8U8p3QwLhhY490sLbJl30H5FLH7dbPU30WotiW9D
s5voe6BuyQ+Ryaj2IBH3CZASH1F7xDaq+vxOmVH5Jj6pWF9dYwcep32KrtxucsYW
kUPgY7SmDMwFjd2M85WeMET20SFRdacQfjGcOutJSpJX5+9hRB3XrvvO2S7IUbrJ
e1an8lojk5jl5WZjbwVoCl/bvr+TtI7o4RT+zGxM/ZQCKhM5+jv5lIRrGGTZaf21
8QAG0QIpQuKan0gskq5bOpYExFxC4kADB42IavW4/0G7h9YpNiyGnZsdKaoK8JbT
YqSKKLtxCu3kRaLQhnJwWoVVJQH6QLPGZgej+blh2QyFL6yoahi4PWIN/77Qzj6W
sHH21f+knvRvxy7XOEYIuF8FyBDvvmKfmvMLhYXCqCHd9jVfDrp8XOa/TaVBLgtg
gU3P7TVINqe5jZzAZWjBmVURdRQey9qzVMOfc3M4aHLmeqd8WsUCKyI/H0atrtxQ
t6xMuRUyx/h+XUTaBootriIu9R1muURwBd82SoJ7E0dhpsr0dPDssKmqTjRtoQiX
419Xez9UsyWD6Ya/ep0RlBmDbytXT3mOn6TDAfaVyxNlSBfKIcsAA49YhJWWFqq3
ldZUri69liw+TqkoSjmBPSEAye7oExHGJg8VXchrXF9BvDtlWzzr6jTQluZaNhKl
H7BRf++H/XCLl2gyP0zRpdhTjqTyuXkAi04UCU9qs0ZoHouQMUrHDvrKGDNVO0wk
RLG6iO3aFuUuchYTQxStYNft8/D2XuejQ9wQ4dyINDPUn0qkosaR7I15IjBPj2JQ
JXt5m5iDPjx1/qigVJRE2GEfOKYITv23qEZnt+yJj/5vDMZQ3s0y1ZJWyQBNyh3Q
KQY9hCXBo7PvGMDbjG/JFiy0ogbk2yvWzTPb+8adeEnxs96/+jUCahsQVug/SiIU
oCt9HovjPp6OsR5g7XFNQehp8MKQOQ9ZuzWZRu8E/HyOuGnBmAk//Xdm88krbhrH
b7xLBLZk3qv2uJlFm/63PDhPcEPcelHKhcDe+zTFZXDcI2I8KWFRhJYlT1bNnBlr
JjqFknQTaVPCnxkZbS65OrwpNK6c5UjtJZbftLFISzn0hSTDuRF+E3YKgY8WJdN9
oNlUOOS+SLa0+jfvAqQmH80WrP1rgSz7E8dBAmHANFCXxPCZoq3tqAs5CchCbhnV
8URrTpggChmWlX4sBtXaQXvlCNHU8/84BKbqdw5Ael/AI1QG/E/eFl8oDdVEmYbD
E+FfOWaeFjO8MEQRbO9Svbv76AYJlQS6x7Ejoem/SORlZCGOtxZd/HxVzg+I2o+1
UHaDR/zkzgP/uQpjPfI3vMuZiuJmyEP0gF6zcG6ODUnr7okrklTK6LY0S+bHISHm
tOnUPrReGaQY7EVC/vf5VPEeXzn2VJPEmrH6pH8iYBeIjcXOmljx+LmmsForQDXu
VsL4eCa/JydQ4J6yzvX6yZ8nXUrnIbA7nhn7SumG5jQp1kE27J+eCaAYqGrb+2SK
U5iHYf3KtgqR7Vnvu83BbZxuW4pUzW0yHGXVf5opmPVv0yoPP1vAQVkkY7dX+xFk
x3Sf123ybXuDEL9jmxk9mYmbdeWiy2Hdk0gJHPFt9Ds8yjxFQuqJ24d8CWp4hcRQ
EJ6Ath8Cy9csG//oUVtg4gjybixu3M+e47v9QHIw+F4DL/b7NyeCC8p3lGrsB3DG
vs1RNnm/YG05WYoLdDg8u09W2N9AFTHMNVWYU8Ktc0h+vhFgRnhDMd9uz8ShEoTI
oEi4O1HxFaUeEhwFaIixW+IJO+1PlGV8MMjwoEoHBt6MUrM8BH2cyO6L9FayEP3h
6oTxsmngTTGpzqcygcbu0upwurkgr8yjrWKKjD3duIBphgMfEKa1JU5Y5BMrOHmc
yIsmT6uFa9znTlcMvX1MZYah4mchngHBVDOj+hK6dHe4PQdHDCBK0ruD3DyPSBEV
51evtq+w1jmvrLGTPVg/Vi1Kt3mL4FuHJ+ctRKxF7Dzx2Xf3hndPrJXwsTv4JDMw
7dKTBFYxwmXuknQQNHj6FDOHhXUIYtVvypK+X+zu3HjNbqVj7WilqFMNQXNP095C
Q55kbKV8f1aPkz7zhsYyCtXVguCkdXYNA2VaJ9MBoSlcCpt1+lFFXzvXsHlQvRjc
1yjy1MlopEaLof9XaKxskc83tKHy6FSwgrwMRCW8H8MAelyjPvRkWbbIgV1E3ft+
q0c4Ec3HwPy2VmIlYecyfYo5Z3qpSIhEWjBBkxyhVaVTkUA7T7IkEsCLrETPTbxd
0y0xnZr8HVIByPzCiCTneKBYNv3tXPcoe/03wQ8+CfHxy0bzMR/FCaUsZ2ulCU3n
P2RlmspyN8YyaVc5c+VFcchT9U+dMr8ednB2yz8kWkX/ZbFc0i3XMSViwsTqv5sV
o2Wn4oRJGxnDjmW6BzhvqoYOkT14l0xUwgjh+L7TPtPCPSY6tBXQxg2XOLaD2FKk
MyECG8RiCToKlyLg3kNO/bfq2OQxho1xLooVfwwwiEMpUSpwpihR9C7bkDCDJ2a1
PP2OCSu0HKOrYDEoNkclS78m0n7Uzpk+3Q0HCDAk/3qDHwIg0KB5twIdQRX7a+S7
gaWQE7IVkKHLltq94nqZAYrTSDHAbTHIIuDkV54GsISRL2wddHHU6WwEWnZc//lC
KzSm2Rv/HOAnQmlgkJBK8ZsGc5RrENA3A3hAi6Cb/NdMw+RDEW5EnlG350ohAqzq
FPrH3rbukPcQuibAbEb11Z/43H4EcTb1ZfdTCBGesQUUZCOIQFr+OxVx1kitGBM0
1jG0F2zf1PwFNKZIUMLRCS6j9cBpk9AXwFDMkfjiyqI+HevyOQh0Fb/txOqmCm2V
PeohBwNz7c0Emxc46bJcnCbNtGPFqfAhTgil6eq6ntGaUC0swmtkHa7G+s8i70l6
u/VSz9L/r+0WnW0F/OkMkj8awIdGm7qBYEAPLh1jRJoT2NBG+PyjVC3bEqvAeqgH
mXIppJ69G+5PZ4LIKGEt9RId5EEfLrFMbZLTNm44KoBcg9v2amM1dRlqAU+YbtLw
5myHEQq4wqOdQwEnkiho+jiZAKi05ym97SYQQ5IVWOxOmIDu7UZEXhJPUAip7McP
SdOYsIheC3x35XBs+r1z8n0DCD0Tx50m7KDKb7PLpOqlM5Xcds5CpcynXiUJb9ff
BEojrGdIhdf1hq7fWqMygk3U9MHEoK3PnVtpl2QOFC3He0+yzM2AUmcLCiPMHhwz
cyZlxxDTY8nmK3m00GmFRqSItBwELpid6FK2wLq9b75g5LEqTGi4ea65IltYvehn
Bquy4khWgiK9o2DnFl5AGySSmMDZUfbu5kuQRnXkWoOTl6p4hbLx+Az9wYQXiGRE
T4b93LZH7Dm7Lwv9BQb3S2q7UML3gXreKTuTZT737O+QOtEoTFz2xW1hN6kkrWid
zAFItN4z/PTF2Ko1Kjzs9EOwcVw4tT1jD0ahpmXJCGOmn5K0vro0qNtFx/8ZuJCT
ynGnJy/pZTRG63Bc+qzYDgiHvWahmA2hZcTwMzl6GVc2+HGIc42rpTJdT7s9NMhU
V8aNs9/N0HWbo37fjULnGeKRvUy9FHgAAgq7j3fxv594Ji46Mk+VMoqqAkmZ1hoz
qlohL/rkb7JHtwUa5ITeqNsqUx3KJo9T0OjFF4oIMhpf00g3WZEEGr+Q0pCWXjnX
0zX6/GEswwFRnLViodeB0vy0WCaQCK2WX3E541bNuP7tW1LdVOku8qoIluh4kus9
qZlQduGS+hx/zBIvXfrit4UkKnPkN3riSmWmhb2u0Ts6LZ/wX+X7vCSv6i429gGP
vLmxy9+wtZYhLZNfpRVfuQy+QZeIyzoJABAH3iIBzPib2mwD6o6vaIDGi36guoHj
6ikCPaFHX1JibPSzGScgmKOIyfLzIBJEbov7BZkJ4qSG5iquFrs762BZI2p9a0z2
PCUlH6BVM/poHpeurwKs3JvK0+c+bQaoOUZpnoyIWgaCtMmQ5QR9m4rV1PkL10/V
iHBbrTspJ5RaBZaNzbIPiDFhWO2lNq3J8ete8/tJpnslUJqr4fo+YGxagCzamNH8
K58JNaE5nL6aXe5I3hHJLh1xRSLJBl78sodcdoycDvGoC5o8uiaPgrlLrUgiWxil
d46sjsRSi4N65iBibH2DhkSJmsI9Cm+fqOiEX8eN7ZTNZaZ73RR4tP0XgFMLJXYY
aRTtaLkOZTgAZ0+uLSIUThXc0gWP3AeFaac05gNRcZrkdTHdRaUpmHhKaw5a+8Nf
dzBR41GxmULib0bQHBIQsW/TNtcqgEkolaFrlejvUEf0qT5ouOw9Mur/ZE6pISe+
TG1T3nnmR2rSOKYDsdXn+CnAQ8lQUfRjqYFyx8i/Iv+mQUPbbtjucqBI30Q+K/iM
OfzUjdrwhobH8noKNro241hoVj5gUJd0eVIO6+NN1hK7p7WW7Tkty+X+22e3539K
denKmKRuTUt1IBGEdpsxm0GGMPJtxBxJCmwLwr0kIm1MW0ABFmg+f1W2zb8QpdsS
rKzyGLrGhTxqB7wexOO1y0DmFcWbHSndR2aflQVCiKDWoPXVHWvtWk2smnFWBlCz
vmVqGm5/PEnWwH0BlBdnLLxiJVZkgRZ7kGEFtMS+QeA9kEhOnPZ1WPZ2vgGG2Ge4
cn9l9bwEjLiYijG7jo9pRmUpnDYxKAWRQvx/8/yqJBAtC+M/OhIk01hjvwLtGzsk
jtipKDO5CbqmJkeD0dos9L0LvWiJYEHQZ3ljJ32sS6UnIqkrpjmySlA1vL2pXNug
dkl3OrWyV6p/6xbOb++kjFof6IuiMVck7IYIlJ7QsecvPUa5dpbLc2tyi9cc6RRM
NXchqNc+39nFvd5PzDmlQTnIsSJYC2tZN0Xi6JyiQw78juijXQwwfm1piPvD0nkm
N82//S2pdCoaw3iu7PEoNsF52zapghvxYLnlAJ/6iOZCXuD/cAUBTXI5LNrZtZb1
waFAEQWplRlWgKh1IDZ3wfbJ6oLeUIf4Z6AHJV+uT9FwO6KXsRx0KWX59hwGf45Y
au1gLWJaFerBzXzSNqLoCe1VnFQwQLfLNPa1efHjkDv61QGT0kqXHwVQ2ixq0mtg
Ad9n96+L2QXAFDhQD0WklI2tBCYJUjI33YyzmccNgDjkKfBeRbDCu4lHfEDEoi35
+p17w1SLWUgam/5YFSMFyf6lblfzDQSNZwnDURP4vxtq2NhdBXGE5J/s/M/Knzrj
1KchWJ77GGRq+NGysP65Jk05s3QfJIAmo3faW6/vI+b3FPfMFUvSLV4x9iwvRgj8
VXUWz13IHkDRYwTs9vlDeh9QSCeM4ivJ1we2fFtGuNk0/Grx6XT+ywyjp5/Lazts
awlQ/FBjUwhRFtvtblghIEZW8J5iXI1VV3GK/rjP3U5p0ztUa+1Q3B6Fip3sEdsR
sSDZhJncfvxX2uaBR64x7vxEa/N3vuH57B2txNIXi3bQPkb09mIZ7GiyxMM7fYiQ
qcN7KYR+zmhsa/25o0Kxveavsr/+v65oL9jpWeYKYKRtyLTdluTczyx2S2joZqoA
fcStsmh43XKd1zvrzKyvPkIjyptmZ5uR1bUXMZJbxuc2NrUJyBIdjg6sDZRNG8Sf
VH7pDnlqpkO8Au6HNutIlID7nodomB5KMlDEBFdps8gIzQ4MhTHtCenUGJGkg7CI
ql7SCgvhWRPF3BYDunFqVhzIMFAHcLkuq8lpnonWZT7mw6kgfUPwNHxsPJIBNClC
4ZU8lbnd3OLyVYhIn5xQyImJigfY351Tr5CjcCXBBrF1yubOu/eanMTN3v3UH86U
7sTL2Osk8rVHFO7mxO4knDzXuJt3lJfxD5zCkY0Khc5QVgxEl49VmYYkIE69spJg
wPmf0qniG07KdocBveg8753+PNtXAKErLfb/fc2WynPXh59ehij+vn/+9sMOmORF
cJoxoKgKeN0wdBERYcIJxVoMr5BKyQlE77QCOGQO4RRYLSB6GUDa69zeHKdKRmMW
5B/h/csFnCznMWwA6O+ckzWJ7BBIb0SHs8UysQLIvBLNUK3bLhszNPp4/DKHCf+8
8NQHlOn7vfN+f+dzOxnJh9fUdEZ0P0XsOsNiIYYVAS2fVxpwKTabeAUITMuUzg2n
+8cc3hYLQuPy6vnShtmtS/SvOovU+mjye9Lm+ZUF+BQ3erMogtWWZiA0Ax30oSxm
fULntElDp17C/KBsp1Sg+0pIY2MaVZ4z4O1hPGjtMcvdlKPitDWcDaixYxwWeBwh
hs9Pc61MFfelazgNrmzeOn8U0n9UlhycQvr9MBjsmCnha4Oc8sKHj4yJGzZLCP/b
kDdk5Udo/ZfkKwPPDgcVcUhkMbFarc3z2nisK8gRyVCsoQc9EfRcChdnsVpJyJNO
gBbvN5eh4qOnZDjOrDwdE2kHNZs9HWb3P2wSjBI5QLL7IR3GPVKWVAVPyFcx2lO0
gpqiAtpM+i4/Jl/fTX/dMdl5TydRLfCZGCuKDj5DwRRJQx8j3BvCcobx0mk/qCaT
Y9bVAb2OHGCkuRLj3Dg8ezfhW7MC4cAUkak3p6p+rZaQrZT3X/Xs5LVYIKj2k6nP
vXn4NickgWjhk2dy6qpjuFlESr2w1T4duURPIml0fgtqwaWLOt/mI9JPB1HPmXop
+hBGzq9B2q1CrjVZEmUa/uuMMHguvtNucdwnEwbcksA4BHI3t1DGBVwa8SaH8hKa
hqgorn6FdwEu5637cJEJyoWIv4PEL6BoaF8+2mmqKsCy0MGnKiqMU9AGV0bWAnzC
7oo67clFXZxGHwKwcdf17KcOFwzGQ5OEuwqZqDvLN79EuzqAx3zEuFwBgVUuDVkL
9RwQweeHKEiQa1Al6iN0YQD1jiTVuGBbCrey8mekqUlO5/EjyBL+1V6SKrgD0/mK
it/6eTMF0cfhDKkmOp4AiiPQe+kSaRjajSzCfv5eQhg7T/rM2JkKH2CxvP1cWmmQ
kMLCdj/QquRD+NvdYuWtO5QSfH5shcYNf9XReZIqClFyctP0HgNtWu/wHLN7P6od
BAe1bZLrXwY14gzQhZNc4Y9AThUojpez6ZRhnIVKyUXRRyxdf5aFJCCIpc+TgaHi
PwKGp3W35VYvhmNOFIhMMZzHCOGd8Fc3KoZ5mebj6Oh0uo63T7oKHf1Fz7QocwVK
b8Pl2eUe0KIe7EBlIlPcjGfIEaEd7zoW5MOGUlh3uIpy+zWYD9M7I3L102z7Q30n
5aTq/xWpGrpkSXIWOmi+Ya3IfMQ34FQ1hw1j7lsom4YyE/CjBQQ0cPnroix1MkV4
GtJXKiTI7EXLD3C01KziFkE4Q1evpSTdK55o78nMMqgAPZyDVasWaRt+Pz5c+pFS
C2p7uy44CR6qdWZeWFZ4Upqz51sj6B8b4wcgQThnavIqJAhRLmFqiJraSdcFMrXF
9qDFlL/IjS4AIyq0kxm1Pau6Ek6Q7UuOC13OXJR7e9bAjddcU7FsuH1qWgqcZA2m
1jV++zwPzBgZso/nTOunAVlQkTC8R7ilHrEROjLzfhu8zrbmwhcexoIkGDCT1SOD
2nO4xe9Vmg7LOuZL7O6r4v/ChzqmUzQA055256qtB46kiW/CwFENFOhXQ3yIvZ0f
58JhVjKoDUarJz+6U/t3iF6JqtOA2WhvGrkkoG3OTlZts0ABaxLkVncbGEmYlijk
yD4Z4TVZD1yKNNmu7/M3AGtVNwuqfmGAu+AOW8i7yyqYIP4jWEfhm7CB1GkTMulv
fpoQNY08DGETi/GWtouFlcZZFO0T7xJyxY3TY79lEgDBmflSR1HCB9OHHAH4jUj3
yJrNi6hQw/AIeWsLaUvg/138bthZcVF8Z2OSY25nM/I593ydwTa+zU2o+0PlOhEl
F+c9Vp5YJlO2H01CUpT4zPobmWNyCT6EtSEcGQGnDkcS1a9V8lmCcR4U2TlVQE66
DVb4gmdg/TKxBkp4VawJpZ1D/31jMVp686fI2dDBYlVa89GYv4cNDz0tmJQj9MoS
4+dRDMQBJ+MMwwD1ZFMKvxQ2c2Sxp3z4ngM/o6FyK/Mph9lYd4BtWv5oPsa7+oR+
6zK3bst24iZ64ds3vduCQ3AE5RlXFCFN9bTj1yt5G2s19TJwfNpXZr9yK2/Pchyy
p0g34oDZ62IqdPonBJ4WSpk5GXcHdgP1I0HNahCbg3RGmRUaTi7yjhIf7dEhxfXn
kd+K4bFlSafnMNpvIBTu1Zln7bYaM8g5e2uPWZTJsmd6ScY6KQDnWEMCPWv66xDC
HlqmJYw0duGm516CsOblvLz93c1C6v0VNfekSy6PdGCcCf+DpZkTn82tFMzlDdKe
G3FSG8FU4QCJjJQxElB3zgd56wrvO8Wf3eA6PMTEYg7lVFcBxJs/ejGjRXSWFKLP
qAT44MN1Nnx9D5QupIUFMDQ07rEATW1Hv6T1kGTrvNctHFwMonAljVGn3i6edf9I
setjUDKFI1HldeFOAfqAlhWF4x428fW+VXUjvm7hdeo6/uuSqjQgzF8YJolENlbF
9QKp8NA+OB5Fl62sNtWKIWQvbso6dA2ersf6In/tcVjlVLbIve2gm9Br1QpKnuhD
7c7nk3AwgwI/8wfcnYQBw4Ap8Cgoy+dx8YDXmyngt6AOJ0CJ1mROujZmPACnDaxF
mZoCa2NgENHYYJ4lj8Pa9xfXaHSZyyUbJ9jLJtNYaoBZx+DxPAph/u/Bsyamso0Q
HrvjYCQhcdBJWK8x/iZc7qR9b8U8nH3Kk6LI0Iww30Vp5411wQEGyscTS4sKxKpv
aDHhx6x1pSUgJbUyJWChR5MeDVbi4aISCPce2CqEQrCTy/toZ1qnNOl6DBbfn5l2
imbimMiWPe9yKAARbtg/6EPr+kik+kTy4jBr/l8NH6tTDSh/MkleLgnu6qucOb9j
P7TfqBjzdaTWfC1rgXPDsdCk5SYZVFW8WwDJLEgEZqfD9Drfi+sEmY94y28UxiKh
nK85ENFksvVbeC+vcrhX3yK846CRDTKf4QtUA2IrOYbxO1f0LXxa5ZdmW1p1fM8k
iuyk3AKLEfrx40elQUtF2e3b715xmOf8aM2TL0em7iEKCwP5ppUwooxEH1OEFnfB
5iwNf9ze7jTRkhDeegXKv1FGpg/OfWk1cnLg9x1QSUzL0KXiCKWY3PS9jAYavd8G
53Cu0HJ2tBiG7OEG7gzlnlRrfE/Jiv4zbTxwovtnt2xk0S0KjkZQ9CUpC+6udv4U
dfRtI/4DG5iCaFN87Q9OWkVCdvrkeRpQohmOWqbkyMHbVO6LXMay3U/tfgoBy+Ee
tA84EcFP0Zo3Xcs7BFZHXggeQKU7kxBD8ACVLMuW4JzG/GCuWhiR+0jd30PHiEnv
WS2IpIjc7C8MtsF5Pr7zeokhYt0vLOPav75Svp1AQyxhZNKnBjsbaorfXNa/zBza
aB2aNzvfYNBZ4F9QV+43+XeRJ4pMhy9vgbI7YZNhauYwUTQ4rfVKO/6b7qBNlGU+
PHeTvQYt6dBuUaTJWv/vq+ETV9umyTcJfFKUGW5h859v2gtWSFe+Zy8HXUN6w/NR
bkTnsN2RZ6oaF0V8pE+WaOoQgyF/MUaZgaeMSbHnDkeFT+iI26RjOx0ejNKSXD9Z
/DwenMCWAmlRjPakHBNfsUjW6B1Dm87hshszlXeB2KO4h+awVKw5fNYn7G1dmGw2
Ykjcqav/EhE5XWS0Zt/0XGYjr1+lE0RtS7BhiWP6aOR9Fm4TL82SfUFqK1TQYzEH
jSxXqLgkiY73WhNAbsg2UxTJPvQrZU0KC2QwNReQ6KgGjqoiUIvJgyMl1eHGKilo
vu0xRKbFU6yfq3+UE3PjlCSUMMAit9KK9iIfguJn4PJt9Yd+MGN0rETD3Ru5P8wM
CwPZa+jVed0LwJ7rXVu20xutnLKE1CXNkIuQ+hjibIXGXzn3ddTC52r6unGLg8CE
37okvPoMGKQ/mEmMbWfvjB7p54ud3qD3QbKtJ6Uq4MVs7wxElRi4iB3xcOdyAajL
bJgusHKa+D6MrmqQBYg1amigG1iK5Wu20p1TLb1b0K4wNrWJ+rv384/nFmqo3Tgd
p66Qw1VFxQd3GmpV86DWmIpzsTAYepBA6ght+xQ1guz1GV+vU/80w0J3FhMz9ERQ
WxLkXWiDbTrbdzS+6hqQlBimlVcnGZ2d6JPuWv+pVL5Jl1pgoAWLMIlIbcc3UkFH
ID8/Y8pBtwVq18FsIZ9AFufSFoa1ktmF1RnABgU1fk5GeBs1jFu0vOeDcGmjTqa1
H8l5Ux08ByT43LCRYN/VrQCVrrJxCjkMjEHGoLt1xkLWNNcwO+c2myuAxgc01V72
91H0cM8vV0Tp2JeIgFAGXKyhKxNpN2gAxH85RBYU2Aqj81cj42hG1wdEgUKcnTjU
C6id4SXqj3NLnTSTBeGqCwn8r6pNjDSGxEAmAZ1Rtsol98loS7yU01Cwt3I7IbT8
hXBNZmIl3Dx13hANe3hLavQ/r4VxMc5xFgMilc/seetb7Y09D5o9eRWSSjMPMUOR
ttBfE8WF4SbgCjr54jEJNGeXEao12umOD6lF+MXdt4rWPjAPuTBUGN34bEaVWD6J
cI068Ba1RG4cgCPr7EKNfAdKPL0rTeRkjHX79Yo0hjIhUYq36XntQ0rg9pwQzkZB
Z59uZj2x4UCJzoYZaUIkC3DAaMsJrbf3SkZkybu9/lnuEBollSa6MmgqJAFhiJVR
Bdd698mzoooGtLkDN4ZJepJqus4zJKVYNfkduT/H+hVZ3JR9ZNY2vtorCxlcne8O
jGzyuLtSzWuymfJZPs4+jyski8TG16tHgjZm3t5541Iv8jHQH+hrwGXRdymUtDfh
OrE9qe5p1hFqFsiRFmSEM7cMT9TAAZAyf/7VESXH9OvuhB87uuNDX0BRkymfA2XD
zA2OeIelFZoctsUz0tjzV3VeY3YrAPRTiaobXVyf36/csaJ73Gk2hy/TJFcqWmZZ
+A36MxfiQ1XtMWrxhQj8LFnGlOuGgHH/1sRfzL8EtmLSXgPozs6grUZ6kZAV2xf1
qJlKh8sEC/e5yAUHrgmd1FfqdV0ipve49A0Y4DGjDUJc9nrYpjSIHsoQG0EERUgZ
sqYm46xGmIvwnjTI4eYbVTlCMGci/2/mGQ4tjvY2fLkGmT0gKdlmm+T0YYOwTLsz
b1SUbBKDu4tFYYvIWdgXvydNQCqDEWTOLdjMVxYAvo89VmTfOgU94GKc0KOZjcKN
A9Ysd02ZUjPlEEiErBXG8n/CMWozET25Ae9Td3kA11IN3gmSHCgh6qQZ+8vG6cm8
GS4t4+ZGnxywAAMlinLrIsb9I+yQ0bvRL2tZKPNuyUMRTDi3G/l3Nfdty/uu+6lV
+F/coijdyeTvYh8FG+IR6aNH4N5ln55ljFs3T8dQX7trh+/MgFNdq8v5ig+v5D8p
3Sell2k7O39uNW8x9aWOk9yfZfuaSHwuN2XPllkxy63sV0STj09ztYljcqtTc+qn
qFEnGlWPDJtKWg0pvZC6JUltrXnoxU5K8WHV6uVDr+MzDjBJF2BrLGSbNXWBBdD5
+wgMGgUMP3WQF8JOxUINlakRxiDTYMBUaEzwE6geBWtq2awGXxuRZxhUEkJ21H9A
THiCshzvXYlYHDdnzSm5/XgAEJJR0ZMvA0iRtPQglJQ4y9Ht3ZkDfOmRhEiACGfM
wvvHkFBteUoD9wJw80qTe4xGDc1OPYJeiHfaztjuglD8FF17Mn79BRWl8btJZjDk
TSSH5zaKdnxWizePJp17t6QGz47amsEturK7BCNAD5nfMNuweWSbK2Tv++Ns0U4v
JbLjHByvL+D4ALm+c1F85/mTo9E50bLpGFPdWW3TLZ1iohCR6lZqCjZ9ITI2Sy5H
QTUeDlHrPhnh7d4axAN12Bx2FnFlGgyKHt9IZWinCjvBDtOIeiB1rtxFc04IXUnL
OjkORQd0sbgIxYtEyqpdWdCrAjaC4Hw8Rj1NVfYD2oEAPDXTNKIaZAOHlyMeC/Dm
qxeQJS/z1jTJ5msfEFuTCTPp2VVam1RgxmbJtxUI6go5bLoZt8a/9tvVSRagI9f2
iXQslmBPaptvLrtHjqHaXjETIYgnwmvTc9hEyuU1nRTZq9klGUfwhxRLQNrkNOGn
pEp9+CvRxfMCdvraauQtM1fRwWqs2nmRLnBa/DN/kPpqi5y5zhhO9rT8jCfF3ton
u6jpv+8FF9UQUZsCgIwknCM8GSzJ8Ouwpvatp4I8T+mbqMJ9YNS4VGMGR6md6NDU
meHzGIl6x2UNPXn+YA4dfo9wE3Qdjh2RRp8b30xEvfRzt/QkaME0Awb/t7ZcJzYZ
o2pwtKvaaAISHCOsSkoZ6+6Lq97eN68GKjRPb0k0qkn3Ofij8ycfSt1um0F+ygBh
iRmpUcEjjEDj7yVfQ1xNFKD4yzQdHxSd9HMQicH1ARihXH7QfvNSFlruNi01ke2I
XkNVpDlj+ZxelWYb/wyRntyhXEUbXU/QdKE9to+dy8U+RqsoBCJGkh3EaFTLi5lB
aeSDDEUCZ7oLIqyVucYl7rGLj5inDmhAHeWvylzm4i6X+ujnElsi9Ar69JWV2RZs
VF8V/B5oR649GAPBzZDHyvB+QtTc5rIzzO5bxO4A9GS+PRki8/yEeT894pMCin69
S6EMHJVpCyJtu4KAo1ajyY7/38X8gbmT1JytsWI8BzSazJJPA14/LwVzBe3SCkiO
SrtkVH/p7V1yvRB4dByevL26DRQmy3RGBH5Ett7L+efo4RPlHBvD+OZcpEAWpbAH
A/gV+3RE/04LpzII7UVLXxvPBfoxEDjJ4wqSoApGo8gsx0sG7erZCwIJI5zXh73Y
ulkRHRKDx2Zx+iVj+HPMB8SEz3yVpu1jmc1siFvlbTs8GvGeZm1Yxri9gfytuuZQ
1M0UEl77jGLzctcgdvKPHlKKjSTauX5xN/pFjm6aJ9yr8jhLFTy+1BtGjjkQY+KS
JbJOXakGzIonaTennhSwISM+bhX1opbtVuM2+GmGHHdB0LHKzYEQpJmSh0zLfRCp
By6bWdP9eOFsZUz9R1AzYM3L7C5phN2HWifHmZAs/iYE8P3I35+dlnTBddpJFRBW
eEusxKqoIsDT+aiIYnfgSu2ZXQu/nb7/cHzynwbVVWMN2aoL9Y3Ia9VY1Os2I/wb
07wsJMob6Y4Qf65WGyRUcO67v6lsppf5qg0fDAKe1SaOQorR/RRRV6drpase78jk
mlPwzYXjZ72ryFIATr0ELj4myR9sjsiCjOvLbWy+uG8t5QM5d7hzrTAV3136UtJv
5DCDhXJzm1DTt4pDndOx1YZNpRmkEWzBipY1Ed86rPUbebxstfe6v5P2nTN4XWxY
9QdbceUJyPfQ3m7QFXahfqXgLQVHC1E2FnBLj1sUowmC3KeZLf3r7vwLk9NlkqMH
uw+mJenCVP1LEjbWLlsj0TCxxV5EXLnkT0lG8E3FNavkz5eqhO8qucaKj91k84YI
a2mFqTgXyIZ2sFbepU14W5QGrOSi8pUKrjF/7jy75hYD7Dd/h88WYIWoUwQGOtH/
ET5ONvCYM4uFQ/S5UH9Y5l1/kgoKVsHIBNRQeo/e9XOu4UxLRP7iGQYIBLMsy69K
48H1KSkdhviQJqpmw8Bhy8jFCkO9OV2RxSNqm9JDj4DeLkkfUbn5HUXtBZHrTXEQ
IKYnxTQdKmco48YSg7LSbI+La6NY642ugR9jthVREWSThIPpnRs+W+HYDHUMZviP
vbkVtu4eIxnd0g6B2FCoNZlmhj9mnAOSESWiUzxVS96HTgJD5O47diy2MrgmyHvA
kZBtyEz3hpFnx17+FrlZEgKrGOhl4fy8wNSH/sKgtaRwDLLoH4ENfRTJqm/JCpFA
Z2wuOoEEHXAYIrMAxFEba7VZoT4An/KXjLB1LV3WO+4eYJPa6FCVOqMOiEkrzcAZ
3xTvvTBop6XW8qbRSiAGrFyUg46WuGFCzasjsLM/a+u7BsAEaRgPz+7Lv5bi6XhX
K8rZDTi8g4JEvD0GMuA4V6LkeGLLNMYh70MvIcoFKw9VIL5mw9hoOCQxu7+3CmAR
O0oAwUVuspVQpxd0wnttjgDKjugyQPJ6orXX59JT9CneSA5I7DeRGswUe24ta5mQ
gwqKjhFyJPCk4sMgKFH55pCAofthgp7qkhDepJWr696WjVMCnW0J96V2vqzaObQx
1ftyZCtafJJDA12fVNT2xDIwCOEyPWHKL+jMZhVF01FHqAudWvjKWp2CiboAxplv
HVHi22g2cL+WiVB3PhJ7WQLUgonGFPYOSh/BTfADtE6hWDkVEw3Pz85IH5w0jZl/
l3Hk6MtDc2xs5ea4cR0CDA0mVoEEUmTR3SxPhuxxlWt3WpYc69GFNnzhYzRhqPQg
713whAAdu2UbApCkMmiVbXV4+s0AU+dTISIbIeVa1tQi/X9hPbtPvk4a1xQm/xgl
kR4mCV7M2KNftM923cN+dhWy6P/5OMdFyXef6XbrbYl3/tJxSshvTlS28qla/DsS
m4s6sRoNAiSKm/HzerowKNxtdrzCRnvGDjQY8+ySSE9enbMNu46rHQl2HWatwCzX
9SPrH7D3WU2rHLgkI8PLiHKqR1TSMM3zy0wRHVd7NSThh2HIuvztaY03ACDTUgu8
QfvMvUhX9uuYZ2bEqD6VycujS02nymHS5IObAkxVeLR+Cb/pVGZvi06Pu3EBFVdh
d+qS0Rmyb8YDp2EAhkROftV1axHvuLefzZQQZQ45pOnjsn2SK0sjDZPxr+Z1Zspv
pgu56XW1pqDrxzOvWRp+L2zxlvwMNcghGIKcmwAg8oZ+2oyUb9Wfb/oLqr2xpftP
aFbPplEq1Qj+uvt7F7Hxeqsljc5ym273JJ4l5vcyOH0AomgiJG/+/bSo4VeLdiyr
yWrPVpMchnM/MFB24bJXHGQsT1KFbBGbEHpvYLOMQ9+rrFJrbmwKPRXdWeqCcBhK
z0Yp5tN8WTrZKPNvBtIly2PgB9okYN1E9HUC32l6enP44HEJf5h8A6t0bkD8LlEi
2Iy4tfGSxfTEkabUJORLMHqASCDR2gfoWbikfOnKs6cDKHKvwFqV7TeZVy8bOCYq
XQB/4AMsM3piKRJB3S6BSSxdsmHHNrHio/9PCLP0S+FPX2gv/sWd2gHcol9PgkV0
fCGTcr4P7plwQFd9FBf3NBohi0vlz80e46Srfo4EyMqP9hh2d5XooE1vzgGElmSP
xrAp/3anzmr06ZrrdD/ueepPAUWKHPeqertmbJY8hbPeL0wLp/haauXZ2eJvcCI4
kTsGcrdgPWakA2EPxYZcQy6FanAaGzyI4fa9MTARTprgYXaGCCpx4StFLmit5ms3
pEthGged/iMsy0AD3u+bZoeHQCJcB6/M/Cq6j2+/7ov8hOLnTWSNSuFJcsH6YPlX
RYfExu5ym+yx4kHs30KwoEIrT8NbQwkDOce4adVkbzx3PYnacZzN7cyXwX3ca6VP
LvXQmBI+E+ky/RJ3biq/aqxU67eH/GYVZEEbkHo6fxdUiZpm2dVT2HBFJk3A9H8u
kb1v8I75HaFA43ca/kU9Av6ePorq55aHP5nFY1iq1MkhmfoBOjh24LgGIXOpHYrT
Rp3klreFQSeLWTwoLJgRMBhqfF2gUezAKz9sriJf3h7QcXQJJWFb6F5Dx6EIi6QD
Ss6GwOE/jLdokvdFYgK6HLa0DPsp56f62sc4JU39xp8DfcwRXeqdRkcbsdqgVCmg
0l8mzcfrrCsrAdej/YGZyXB59WbK4abngN9xN6IWstym9kmZE1aKWsoUxivgQjs0
LJy77CIWbC4AKSSBSb2AMoljTUy2JwxbrD2heq2W0jyckT18VMT3YUYtw0vd4U4Z
aUnPYde4bYMf305fIPo5u3uNcflthW9gfOMw61OWAs1A6Ob15m3ogwOC98tRlp3G
6lnaEvriB341igA403giem/VbA+3QRnZyHuIEQGKY9M8l+xYcd4bFnGgpeQN6Q6Q
x2Pum6UJmdyVTrKuAHrgl9YR7J0zheng8d3FR8bByRDJrAN02Vg1AfsOMJ6Fh93t
hBvwhlNmNMvrExJ8o+3Ne7otbG76RvKfPTeTX1RY0ptvdVHNMc5ji5PbQh+xwsM+
axAQMi+Y/2aZXXgbvBNpNX+U+n//KIMGmH1Quc1M+M8GNydMm+5m0nxb6/dwfv15
fNRT10CJD0W8iG4Xs/u8bLLLjwixzcdIIfkWH/0lTJ4Q7c1WhAIRku2/Hm3RjFp0
8aXj8BDIfXTjBIiBlMV62lX7IuBbOPHP48poOFc3laXiCKiIax9ouhBRFpganv8c
dk3cuznuqg6ntgDKH9yNnc/a9q/lFxRIjD65V+tnLGrX+pUMzI7iiCM/Y/ODBHe7
NcM7zKkK3tN6+ObGu4Vqz6PMqWQvGVETFTA2jDkgA6SR9diBXE6L8WqSMn+pgUOA
OZuIijjCbyPX6EvX2BSaKEl7L8hM8+RGD89zub7D+4Xtoc1qtUxE1Gfdp1G7wWs0
2JCAI2g02H/MT3OBgq0nz5mM07rhNTD64kyWdZJ1B0Se5o3iYJgg+fgqtBvI/ezr
I79tHZHhZATZOSULbQJncrm8prFzxDqaMuoJ5TiX1U7yMXXib94PvjsdxKIEfGT2
xxs7VlTI4/Q893UigRgmxLU5uZaFvIZa8+vp8KDMDhTQE+YJkvN4qhvVFe4vKdmq
zm4RRBGwJ97dab0/NU8gJucmFPGSkn50MmWsA6EOT+R9SXVCvG93HAHIgKs9+SOQ
ubPyvf/PWohlxSkkDLstNlW8yDA//ZlbdfwskfVnCfmQHKO2RB3rvJGNGMmLY5kV
7yKNvfjykeFgEywzg3+oV3BP6vpatdMaw6E2AuZIv72ZMcnRZDwr0B8wWtOFmMxp
TFM7R8N5+gRU1jZwzg5FSjhgf4CTG2/KabSMoj8QBY1Y7wTkZXgriZbbwOArmdVa
/5XyPwwYuwjnI4TfPt05czOZFKb56H2hgr15TRFDda/BmLeR6SLQWesef184YgCd
ZvUW3FXxtCVzFq1eopfAX4ht3ulik/H4x4xK40imLu9IZxRksh8/epLllEfNyEKS
hrDCVyISUg3HodwrD4tlJ2IvnAAPpgf3cj/AtP8s8Qs0Pr8fxds1aL4NHfOylCBt
EjFhB5P7WRvYqZofZD/b+CEOAke1YyQ/4IKXfXd8MHgzp9nbluxawAadn/CKcuWr
jVtfoqpR2NfF11V8UQOL7uAwJ8XJcqaz3pn28yKIbsCLwdvZCNzQPW1AI9Doo/gn
JesAB0etv6z6QsHB3NQYgA54Q4AXSWeGvG8JWjdCnMNj1LDtss1IiPOWa41m1VrN
DapcNZqjJwu/LSFXACSO2P1WXMgIxY2LgMXnCRXRPAE3DbvYtvt4lJKhkVOn/Bg/
VYFdg20TbqsQLQzZX4ysCJR+rw3WL2JFZVo8zaIbaYPPjTDGNHoJqNQHbw1/jK13
7QrkKlOmbUE7OvYAaPw4kDv9C8agfk0CksbuQzhR/6sunSwH+4UCIACz3NulKnaY
b4o/Xz1iu0V368ah9PNor29SwyZSfbJ7IcLjuKR0f2XH/yGjwoKzVYszOOTHwISX
N3Upfpx7wBly3EyYosCl9NZoXzsDiqRMo6VtN+got+PU+CbhmLkRkQRu+hqP5B3B
83e4xDs1O/1qgN6oTnFvm0zbZzXPEQjZl8S02KfytgFAt35Uupfce5dzJFQvmgEL
R6Oy6QV0F+UHnU3mg8p/mTnD8W1hou9aacNiG07ykRFOaC1mewTkCAdymXm7gpVA
/CBL4YhavsFZbFop1JS4QizA69J5L4K5JNbCD1UilyV0ZQwYgCxZC+wdUhdJv/JT
n+kiE+MdISnoZ8fZ6YbK2dD3eqRhJIaclzo+s1YKX/pIHO4JvBJVZvf0EzuLD55O
Ux5344k3cYyRkvEbH6y6gIzCqFYlcH125WnwUvrz12nJy92xkVg6j0Z8iEdsYCO8
jXlcpYhLhE/xh8AFTar6+KM8nKeIQv1VSbZ/+GwZ8DyzlVV28jf/CvZdclOh+wfJ
pMQ99Zrk5f0RrH5rzFtefGruAtRxNG5qJ+W3PPtu0M8tNMvE37Cwn6qxk9RW+Y+n
30H08wTWj5sRlQ+Vfh3ALZ88Ty3wxa9fkIITK2QxK+hKTZ3MG61MlB7i9r7GaVlQ
PnL8fEkiR3bl9Y7qcaRqnmHAFUN6SLEnSkjPrMgZ4CqBmHP0NDeTLYYVX2E/bkgh
dKjesUmFTQMMOCmw9fX28GBpjkv2kGdZPyJSLCq9pYwGSixsDMr3dKeYE6ley9XA
mOU53lijAZzqjSEI5OXEGqawXE6djxCWNxdHV07BoEm9apXhHpe7SHGKHLQFazys
T1XGV/2AndtclBXNXbERgBiCVDuj39dIUES3mvpuNVSeztTAYQUImhhgAIO5SqYF
aITE/OJy6Ef5MUKL/D+u0HeGwKOnzEvupd5txYvjQGCAnq3fUYB1NTkX4hsNenOz
FnYP44aIOj+fn8a6QVIirnCtXwBqxdKkNSkiF0j/jow1cciZ0jNzFw4a/bwVqroD
Gh47oZJBgTY/gdg1BBWjpgUFAWjFFU0KXbdFECzYZ31XKZR04zCERVf6njOlnJbw
f9UqeoJ2vMfVDf2awyx3klbqaRojpRPb4KhMBovxQiqzvQXr6djb1/3e/osPFlLY
Ho0vUWkbR2PHBcacqvx7fyTovHWYhEe+lO3r5/Le22TTlM0+EhHzv8Ay/TPGz5du
rxJmLsM/ukv5XAyFL5bZtRtjHjiPISHnp/MyajCljpfDrCe9lnXTI0y6iZcwnsKg
r2u2G7JqBzcQ8vKb8BrRtF7cuXVt2NmA/EJICoUHRj6M7YkH7QdiSoSm1e71Y149
+O1qQa5zwr/YBrRF6yDJ2z8TIY6oVWtMVq7WqV7lnu21IQes+woQJYpvb9swmbRM
azaka68nL6euzzhTcX4UjsEaioSyFSZsSJyY/fGpMM3eZXv0DThXt2Gwj7i22pX9
7VOAMP09Y0ThSYJ6VFqnM5qUWvY9x8dkXo9134wMSDvq7bd0TTP1SPBpg5WK/B/A
pHFXVJ0Tn8ZiRTW7rX40EpVKAhRKGBnm4XSok1HCR4VLoa0QlJpCs3iLX7SiwB3u
U0l8+qLfWPsuBTilZoXeW0IXw4MbEHGbhLLZkZBLfDZyhkHJX9/i5vQw+q57NChW
aaCspdSvPH27av1+pYNOCuMKqTXaYkbyn5/dDFquYpleLkimVbOSwXUuC2RGaQb9
XsYeU5YFdqflwOC8kEOrwTQJ6svxELQH9IlzXsuHGW/OAD50zm03F2GrpgH/dJ5B
m5nO3n2Jk4zr4VYNV1jmz2iq1lAry/T8wWSd9mfRTDmOYzwBqAbDO1Xhx/e0o924
qhjgvIQwlMqkXhek18P+U9RbB+7UWHP+x+92LgSVsmfGfQp3vXcRUiZz3LlYPJY8
e1pxDtvO1qxsxuxbRJO1fAwXAJzXjKB9vKUzvvKxA1Ukioxu/gkGKuHc8hHsLuZW
BLgMXaIdabKyua0+qFNtSCWuZmBBamkX43HTQCJhO5MaNqrFvyrx09jmxk25VWxY
YY3/C9ZM0lQ0JBzVklNUn4qp47ZcpFptGnggVmsg4AUWFO7QFzxHt/Xq0SzHI22g
anya2fCLH6IW5pjoj0jCMLbJFWK7bOzuNXPetS5oDVvzU8NEx4gM74zFdg6Qjs1p
kWcoLuqgL39AM4wZHswBWIkC0iKZ0PBAwjd84XRP78K3mN21rsrOz+cA6WTPJEAK
riq/8HKDnjQ+a311e/154AyaW1O3Mwm+dA1KkzJOv66w6TlKIvjYiSn18WJluTpA
jiPxEV7nLCeEm6LpNOae375Cj2iyLd0k2xZKgKSzZpEDScdWTKxT62Mjrl8HWsWH
pMYPAYYD+yJk+2FyRF87Jobo409M0EHHKZQYuNWUzzl5H2vO29/S/y7ZX7GttVLw
wGxO06fZrtlRqsl2xA+fVca2LB6DiEyvMA1QeQBCW4+uAI719zbOuiJRyEbXbeXj
nYv3oNGsVb0vEiP89gXUDcL/VV49XBQcT/+pgtUvnZISfXc2eratrY3ONpjXeX9I
ruJNtqVtNBYZNpyARPqwN2F5rCE+k4LkikSbwFAAMhKFnKAi7+YI0JJcYly1n1HS
9CMx9sYViCXLSawSRw5KFoFXaVrapjEgzUpLosBmYqodBefQZVKJJwX+3bpn84sy
fFia4GdPmHkHHdoQmdojDlja+uB9hRpI8Q7fQex6wxxJeH1ulSS8oow0NFInJjuT
M89Ik+DNWsJ3kqNYK79a+z7E2zgNbVceUAlmntKYEvcgODCgZH+4FQM556/yzcz8
4LhZz1HbVLG9AxdGYL11DFz2EN8t8q9RDuOkbgSaEWBcc1Jm3hHN4jTq4P8fB0ia
1r8SdmE86+3UBYsMb1q+35fgP03p3qFMMX5JqDzzvjV/164PBRYV4jD9zoCAAWjb
43Wx7CQyR9T/1Qibqm687QM3+9rtzQ7lHL5uMZtZLgUAyHLbK4F0j3pCorYweXnd
QSj2MGH12Pfh0v/LQ1BNsHUcbW3NGaJo1KnrygVk6xGxT/+YT+xjlMU7IGuAu4Pv
iI3zkMsWBzM+kxtL9sBp1P14qoS51yrbzqgxy8xTwPpMGJrxYio5vehVHuvIzYPZ
K/m0a3t1CxoC/aJzm8d9NGvfe7lygfrLM9LVwvfOih0u6H0fby7uqnaKglRJjz3d
CW/Db+S379e1+iFIbsvKws8G5105+83RXuZc6p4X22UTyqhMfuQck+ROvAK5A6ay
6wAFDx7nMTomUPAJziWhJrbhyuI4PEZXu+LnxpdiJ9A4fGvkFn4VrDiHYBh6IGa6
mTwUUe7TVFsJcV0S7rRjEHgjuOaeQh3jQR/tGMfixD0O9h9OaVvCpe0cbe3DMXHk
vvn0EVEwDuAYuf7a8PwbQImIqMsNqjHbJNema4KrYZAmpv8cB5bHOECtrgpKoYvn
a1OI4MfSClaanaAJGmu+KLexjMBJGtXTzkq35fgJkihH7NTcc1YxYHCaPhrLjuYa
lFO+yKfLXoKnrRHGf2DZ+nsSABYOyEpSH0HNAvqppSTuOGOB2bS0KC8R5upazcYB
6WuvZIkusInKpBGhtn8WglEQ4hmIMD9wIEAxfRblewEo/tF2auHzkWo6NvR9tmAY
I9QWoasLJRyxX+dvMKnUVldTEKsdqCsb3v4yXOXkLixlG+sUF9Fom9W3EFgcQ+9/
m/EAtI+Vcyhsc0ihyROBLffti0RiGxK+d0Ipb5JxyOflIVmOrSFHi0LjagFBLN6T
bq1F46X8vQsaIj9ThYGEqzluBpjOwWdu9nRJF423RhfjEwCZOyIe9gVnU65gjy6k
aEZfergYyRxXOhtdJuWlkACMo/GlKpqcAz0J6W1Z0eldoWdz2HUVv1tTRJ54TVTe
3QsGjcZQFnSyRo0oxgr5iE5gL7JgFeaa+hNXEagyqmR74kDD9O3ZGTsgZ/Ur9cQq
M3REpP7krXtt3OIwQ+kqoTXj+9SCdandE+GClI3ekjgf637BRDSB1InrODFwIUVS
s7NrD1EfiUQ53rp6XSMyMWIcmHwKk/N5nSPN464N2RMa79ZRFf5I9tYgbnItXhSR
y8IiFDKBTzNBOL0X1bdtBhpa6+sRl3Wk373rOjxrggssboFtn+Q94YECidYUNoYA
P8PrH4ID0IvbIuKmnyhJZXeFHbHU8jz9UgDcrmoGwAVf2tw/FMBkw2JoUpjJSX2y
ZzOqcfKD0wcYUXB0Ey/ZK2h3C9/S0Oi3+7LyHBDIR2GD0+7LbzzDCDDfGUtetv/0
vSfkKEnlVkPvLo1dTaOBvnCEe5YwrR/qL75QhT2tXRcqXL/6LE4KT6Pqy1cexeuY
coCPGGvnisKm70TYrlu6qKnICuVXuYC7anDmImxiILCNb/UxTq/JaAkMAOKl2I1D
kziGdW3VEuah7h2ECAIS+MeVsMNMUwPAhRuEbrdG6l/H1DMSVnMwARBZJkYs6DBj
F7wODWFY0P27zuAQ7ht6XoAYUshBhH9TYZ2cMBgAyYZds43LseIiUzJ8mS8mzAse
aEI4ik353BX8vrjBZQCe0ZlwPEbu9gciNbvcVihSUzwAevnkitCqvE4uT1V15rRI
GkJpmvaHdshlZ1DxuhpcpOlGc+M26dMTrjPWSAC1ObNz+HtLOVnGNo1agglMruU9
wL8QYAqohwCSFcEze8zHac6z92ysZnziDE1vC9+6mcepScEDxQ/kvz2HtQ4LLv1o
LW1K9VU4Aft3wfWLyu1/gQUY3cv3pM57te8TehcRgMdVm3/sC6P8fldjw1HQPYKb
aIcQcRhXy8Fuf+A0RU04Zd9erj76NPOpwXv1mYqXJnVqqjFlibzB3JezO1fJP71J
2tJqz2FLm2wEj2VGFNl7O15KfbF98X5og5qifaRtR56EXcTcN/c16foHWT8V6d+9
S+uZDMDK0mCHL4BuJR+/IsMKCvuFGJgszy1YfowWAV+5CihWsOZ0doKkY5In3ETt
mNO3ZKIbqF6meLyd2LtKVIeiyS1vy1AqBMWkTlzAgfi+ejtLHU1nHYmCMJPlUUjg
BNEKQ/ywU5C7Mh/mMwRdV+KUnvGRE8N2kSz0nXzRrpPoymOr5MH+L4QKxn3QEOcV
kNlUzkBJ93giPUtSY0iZlLLEomIJZWJAo1NO2cBSnyW5CCjmHvWEX+sy0WxtqVI9
+2T1CoyKWpaFbGMl7l43ZbdTXWSld0S8nhgd8G/ogWORNQS3F5et+3+0RcnFWUyT
bEQDKheFTtBPIasOATE9+Q9E48GsigIqWmarEwzeWoLINNnYM58+YacepI2Z3puN
aimIk6uKW9aaHcwKmXfvSFD3SXWXk6WknlXNTSn+444p3TbLOQxQDDTBDvkhVa1v
qGF6NHpGp4kMMtHHsJIQzVD6Cy2/81hnVQmEwXUMAj+83WwAMzLXD68yRjmZAGkK
oFpSBGrsgfZPEqjkR7VuGP24urkitUS9Ze+YFB/tft7vro8fi3f2dShJE5rgIdQq
xRl08I2RXtZkb3LWIWOFV8AIrRhk10ejpFK42ivi64A4fv1SM8oSkPnpwJKsTvD9
Nx51hiVrjtJQWLn36hTKicnn6dJK/SiODIs1WXtN8MzLTahQd+olSvx59X9zP7Uf
7cvqHyiXXCUGI5O+zT72UAmw8kMflPgakd1ydd2LGNE50KJa/HMih2NRBcSSkxKo
f9O+GexHvRJcQ3+1MoPadg+vk3FfFOxPdO3ldRR6N6P2EPBTlYZZcdwWYtKOqpSa
/IHte4xyn1rqxSAPGMch6Qsg/l0gKvQfZ9szBgWUN5XfOrM1HDx90RdAZxW027Rs
LVr0l/PNGvrszqdppb6lwvSJBl/iiQydmEOE6iEvFeX3W0EnnIO0wgWLlNwuNVMY
YUp6iOJ6hC0REaEGCW+fCF5LdXBK1RBVslIELD4P9miWVfzUbHjsoeY3cHNNS61A
ywP0e+DUt27Q6t6h1XDi1VY+rh8pLFvR6VTSgXdINIZJq+C8zxn/Dew40330RdA7
HlSd/G7AAw7qfi5bm5fNlzzycrBF33gQtQ1/rz3HdzK5WRd7rO0Sy3SVF7I2Ad5H
rtrUe9wYJbIiC9PiKZlkVeARNVoeXSg11lrRUZIu/VOH/R3tEwiFXDmaDa2V7iVG
I1MDON0dBvA5JAbQ9B1mW35NDKZZp86fJcSxhXGSy9LCfX2+Y4wRrxPjbcvAjaD3
5lYkNC5OepaK3q1ZL09/emP6zkcJ3pfazc3rQAZQTaBD54kKmdTnIi2kS5wSzwnd
99rr8tqHl6reC/nsOXAIDMK1w++nQgZjOuNPHlX+LPiDSWuwwm1BJRv1z16zVbm7
UQNhHuBjWNE925rwLyMV2b6WboCrVACWe6N7vdGpTyvzBsRKfp31T1n7dd/jdeOH
yvLAPGdIZ3r0b1BhU5Rfn6O21nJt9m/L6sGXMEpH9seVNImlbuOMbisODqnDTMF6
e/62Ee5Ik4R7qeprI9WusFRKK53qpovw+pmmQl2AoMHqard4QhME2Adwa6p7ky+I
H/X62eUvC40FInS/IUDYa31C+0Fj2toSDe/OVxfPpK11E0eM78mJwBp7REPPL1yx
K8wSl6tj/NZc+tSapp7+GDwzUE7qLAJOTtgqmzUK/ulBstllFSQ9SB93pM9DS8G9
2tFi7BfxQnsT9LFjdYarVuFaOJgvAd8CBwJCTtXH/+9JI1mt0Rc5UfAMIMLy1SZZ
Iy+c4946sEO+OEBM8GSaky/KgRfj6c+4wZ1LxFv8Zlb4dXT86gcWcX3Isz1tL+kp
aDwB9DrKLddS/jmbivZEya0oNxcrsOA9G6g/RIApl4G5pa3OiOI4jUTYqwiMmozj
CgUG3/6aRGkepPD8IQDZsX6DQN2N8WN38rn44j5bg5Cznu1ji4c9DOIVd43MbWVO
dB3DqWkcyLWshvli9YVLB9Ucx9oA8rBSsIW/wucQt77wuSdGGRT8BhWl/dP9or8B
txPI3hg/5GZk3TtgT8tidzbryBZtVUaBIIbiBhllXoBmcDjw+4dbCpmKuQifSjVM
B0GVHzbyzgzQdlWeFrHlXErzCJ558Bqt4HCVjN1K887Qher4KdGjTtb2rl+tMUZZ
3npQUB4vZYv7xI9LryBhzlCSDWZeNruLKB/3mPyc94+FEIfDl99sv8TpwHhYY2TW
i1/ZAiOjcDPUrlpb4Foc6z6cxnUD27+z3In5bQpqU230KoxWnmqB/C3FAsFXXezH
5PGa8vsXLHxxTpV8Sbv0cYusPGmbiLeZKh3xJrOMVf3v6OPQBowgPMbubN63xd6V
LkiPthod5eh4VfhjlvQgxT2TF5wRDCHxvPd1IYK9QH0mhzpyWbmvqSJMDT7O7Oci
MXyIG02QMKZFExJC0KlkvJK9WovDhuywX0s0NQWlW4Wv7DZ94DuyrwsbBDoqRr6F
p5sh14Lbkg/CwPpftocRb+3CbCwuJIJP7KY1s4Bc7lHjCdTlxLj4iwF/Hfze03OA
tiDoZhgfL88EVM1achIfLI8WAXOQYwvX8ehDLeBVCd6BhSepQT0zlXuSA10YhQnx
9zFS+xiN8EoIOVCjlCpqhxe69oylQPZHMEHFXw5FZgxqUtxkgKNpDJSb0gCB8oHR
ZMmCX0oq4YyxZLi/Cb26xuZoOW65vtsV6ahuXwBpikd9FEGBRX34TJMyHX+DxMFh
SELAF2GKiUN0xrfbvrGS6vyaRvhAmUZ6zj0kMADqnhG5hqWfjWjJ7bQmABTz7zJt
aFhRyZEBl6sY67bNDG+bSUNMGxa8P+jqZ4w2pZLzSKK+N8Avrq9R+dLfVq03CdUY
Q3rXPewRx1QCXIzs8O3bXKWKbMBA/P9iKlkZN2eJ1Ztm5rIL2H04M+Wyhcfj2O4U
WYs7DWhPL7eGALdw6hS1fjptKqKnhSSc5H3Ii4OTowaZVVz9KeW62z+sKXqxjUBK
lzIu32tbEsLh/xZixGEJfh+Ku3s5jbLoa3pUN4ZTCwIu6N/W2I2vJJGRKejIDIGe
3E19lkAp2Basc1FHcob33byBKYaXOmVgXAtl1i5qYNyQ1loTZRLJawh0aSmxx9rQ
8tMRPt27ToGn88KQeEML/pcXp7S371fBU1Ti21bqCjKHOB37EsTiysH0WYZujBV+
L/K2PpShUXqefo+mS0SrpeFtv/abSRly1vIywY+Dba21d8nTIyCbvZnxcU/dNP+Y
iGm4uQ9cJ73gcBaXSvodnvIzO5TwN+jElKT9/Qawyf55/WjBmu/R/MsfPAXg93FV
/TNkybfA0KGtCYbljAs+N4fB9CF3tqjQC6R2GvVNy0GSj9nw82Nb6tjzsyQUu4gB
dNC68XTCr0xAjFfy36eCAXARbvpDMS0JQ5UMpDTQ64UaD7NM1a51pbHwMf4E8dwf
Bv2DLqvePu71g5FiJ7DaCSxIiynUYGqeI/U5xiAuZ4mKTDS2nR4RtwCdCb7NVChK
y3zOhGt1H3J0GzmmNlr8oIzopwsYDyErrND1jQ9hhsj1wZ1Y/KMX4Gmfwirq0d0l
/izoIK5z7/8rwOJLs7evZYrFOXULDtnd1EceLjtnl7EN9XLTpqWS77kv+m0MZzmb
RqQQCQ0rHCQaNCmUILa0aeMurCHMWbkiHVM2YjC27fUMXHBakvf3eUsvpHCzaMri
p3IgURuDdpt7LXPgQbbuSDdUJ7YDoZYQRW6zQudYAthPl2Kin0K+W8t4LER24PMl
vptNEk6jJDG2Ct5vLRt66j5xFn0hDPZPnqYG+4i6lJiRhoeDu/OE/nLo5K9B3STh
MikIYucMfSdfva5D3x3ek9jI8hv1zxmAqmhmkrhMdXM65bPlifrGrIalzNyyl1Dc
gg10LwAjLKggWyb41CGOOiiTBkIwco6tAHcZbK+fpGhvHX9JIDYMOQbRPPIJjW0/
HGqrwCWWle6VACETu4z0DfifpEFgn1GELV7ugZgmtlnrloTUgfg+Sjv//4mHXqx3
Y5MSyni6H4FnA/s32936pJ6RN15DU50CW49Hlb6TUP1c/TM0Yp1w4XKcpAcbMkVS
FbHpu+cjKWZxSRyD7zYVSFjqSpNCLG2/3Qm1dpieOwe4MmI4rfgbhcbgnvQTEqg/
P29eCuhS6sdFVCxN7KGwxpe8OW63qxy+wDO+nw00+y0B106YymdmDsf1ue5LY85P
WmuL86jjdMFdfOdlqDqoHNYXNu9cwhuUZXyDbt+iNcOmO1Vw13jxTk9xURpp2Wc7
hUvAbaQP9JxHUQ0lDz3qdwG+tYG7q2EHt8Pm4L0w6dssiY6wykt52/qf+JQ6nslh
/vgxll658nJ2lZNFdbkiVd9IxeHFFKPN5aRatn0LZm93WAU7MDGeKeKTqqOgKuX8
jGbWNCWpb1IWDMvnE44gWBSFn8Vvk83OOVqkNGEK2+Rh9AfjfXxtofGsF6um3V8X
ZO7edX2luzJqp2kQHFQQWzeed1UcYP7JF2g7CY5k9GVAAPa17EdMpErPjfJzRgZC
njPBJhY9h+u365va8d9wuCiazPMI7Dm4XC6rjgJGqbL56HM9G9JiuJ4QKIC3gjLN
o0xmjEwJnJNkPdqkG+6dfTpJWY5osu7xt0H3nIoPLMfcrIN5hp6fJ1sSu9Di+5m8
3uSWvrthzunltYIooQcALdsImc6UpoyRClLMPfuqT7V5KrRAqkuCkLRTbF/OrOxx
NGdnq9XwCT9uDEKz3h7zq6pr6QpuEkysFCxJ2lgoudY9H9PA3LAj4OLFJAxYZ+10
FGF5SqoyWvFrAgCHcXU5gKEDKRKzZiH7GREPeOlLgzksZ7CIl6FscEA7ddvaAqyJ
5KhwPi6FeTJQdA3JgKFajR7E4ovkberWytCeLwOLK7UXpSWA3ySOlNgMLiGV19q2
M5AhajWvfR/aB4o3H/4fCrfQ1eD4OsRlnnMsX1Zg22X8bY3pLUuMlnl0bnF0/UHl
M6nY76RtuJqA/nTSyGdzwiQEB+woPT5bSwZFcXaMfRzn3VgrX72oD/bFZwvYiQRS
UQYp7/JDNCsI+LWa+fZpthFDL5Cf+LiJy8qvZxQb39bsDKLOfd2AaBendzsLxMbo
R1dXMZ7oLjNPHmVUTnzl0I5+3jo02QTTO9OuxcBavBUmeuFSRuoKBPkM12MPJvPl
j7makTt3W1h7DjxIymA3H71okdB6+/+AXPrCZYXbtoUAUOjN+sOS0XW7iLzugY6b
EXCBL9l1VgIRiQSQiXnjRKkoHy0wBABrpBWZQ8aXCgXdGYhNtSbC7oLQ82vafVGZ
Esz3irlaBP11YE395zEpc2kei7bJC9xPcz8ZPG0YS8Dv0mORVODr7nFUGJz/rL9d
TaQHTAjpvhcJNDCQn5z8zFtAEG3jTUXmxEPtRusvOlMIs7pNOwmzO1hZ1/F6iPSW
jPKK5GBMpHdLKI4pTcv7ZaKouBTzOr8RJZbMt5KPOUJsPsB0clxzbPfActCiAedj
zqEVJN9varQlnHbfMti5j0fe3KOtHw4zivYJ6o+heSNf8oRTQVvvVgoOpvSGBcmB
Vzde6+Ck+cZ5uEmgMSp0It+VZJQPSf6hivuTnEkPGPdS+1JyGlEc3Ifi1sjifjII
QM7gP7tdLQyTPH/PI8AzFrNHmvREj5V4ZmM2Uj6slTNjs5tP/hyHay+PlWHRRkXX
nEVevCjMz0slQAZk6k9ePtyltdEJPt2xHdl6Oed4KatkKcQ3UDIgeoAhYRzglxUn
JIOaLNnzMqtVOPJGwzVNIhAFFg11jbHeoup1z3DDDCeoxQHzbgTBuyMivphlZd5X
ZbpsN/9GPAVo3qyDf+dC86NMP0nRvFHq/r253ja/wUBXqid192IOfiDIEITwhQX3
bMDY2qgLvbRVIwos7hiWXIyDk7fa+6PCqs8jWX4AwHSG3hmVYUWzCKe2TO5eyLI5
q0mbQzaXN+15NVHE3ciQ/AtOiecq/vIzbTI6VpWpKCChy+da0HIhbADzEU9YHpr7
QTq+kJvXzfFPxMKRwXgsfOtKLEvWPfEkObzLMwBGH/WQu8tmJVuNeTb5XJU0K42E
zFczLSz+YqLw23oxmQwGf154AAdMn1KlhDb10RjzK7n8lJBTA2ruoeS06f0/tG68
4PieHXkxNL8dABOGGHYt/FqnvKyXpLIZxl8YzfRY/CeoeAesFBo2lvL029Vwpl37
EbnSLklDP+3rHkZuQDrDW70jIEpov62/uZqk+VWgZZ+Ahq5JVpDLHYLCRfLl8Aac
cDmnzQlZBkA/Rd4FYYQDJ02KrFLvpOJOPOGR4QWlpnLonxNz4fUfRYaeWHT10Gq/
lmrAX2K5X46/Gkal1MVle3uuWP3AjTjdzdHeB5sB4mN8hky5PudaXs4mk86OTHO1
wt4m9/Lc0dM1WQrbHBWxWQj3xuCVppFinW8VHdiFCUfDb+BHZhSeA8w3ro+zoPoy
SFWt63BM7byQFQ1JsOmcKHvf4BdGyN/ZrhUOLR6Koi8ZKNmE6ZO47th+zWdB3hkO
RLRPkjWXLihLbSnNDwjN9YztcqrSvYehkP5fS9Xvdn2rLgWQXiOyqrIBIM5kdu32
D9lyljfMmkk12FGVNQQdRMVtV9lSWCrCOK9ml43iySs1QW7txMl26+1Lmwji8EGG
s8JqYUD6KUZSuDyHiaPvJQAHDRWo2bbpRzF06kd/3FLZ7OADQJd4okYpnGxVz6U6
Y4ZAuBWYnOGHUhtr/BXy9Zh9a7C4Fj3QIGlt4eVwKcQkuvOS5Lj8pBUKO+KyLIF/
O4uXjKWonICMd6f3KBsaeVWw8NE/o2zGdMZdpcln64z0TirP0pTregfM+ef0I5HP
8S3ldhXQXYmk8EqP/3xkleZmrl6DwiOXDrRRYcPrBHZ726TNb1oPnwG+sOcFPxBe
i5PNytrw9iKcOwn1KQfyFZJPgKRrE2VzeVU8Z8YnryDCeFI4buAe3mGsaQ8jIEl6
H8R6TSUqY9ExHe420nsOuVfEw/f5pBY1a47uPsqaY150hxGrPzc8lnzgd5ft7bYz
QIcX9lHiiuE/7UzLkTkIiAiQjxDJsUF/+wM2+M9+tjZF6WRIbGNWI5dM1AhFH1HL
yFng299FGE5U7ZcqERe5BlNwcTpITaLJ46J9idCYywmJkZoNCLym2NEG8DGVwsiy
3Aze8DJcRoeZuT44v42nbUwE76UduBkRb0QaQuG3Bmw3W855k5BgDiu2B1vNmlRZ
mIkTVgwRwT3bfGTwHMxYICRtOe3OtlX3nbz5yjPgovuOQ0xx/KbqvofppT5ZegjD
rqqAuS0dOcWp3R0Ao8LM6/m0VBB5JZzrQ0pAPkrDzccaZa8COKpkb/HOhEiCh4qp
sRC3qbF2+VS+zjfgmOjGRNkw1S1aBBtNtKAzeEnydzYyQsyscdhSAN2vBXyWO332
DDu13utzKXTwG4qp4Gh79XaNjqk4ZC+7EAps0/zC8c7XRwljIhsWTvob4WUKk4mi
56RVluW3bNNULdGDp+IQL+ktLwuI2BohHIOM7m3TInxb0+ktNVHQKEsolsXAWq6d
D6UFhi9heXuzRsHIxn26dAZnQoM9gp4butfiRftf3lHLebbRwCJvmsAiKQMPKKh8
rpB5PUKqbWPjeqqx3TYdhJnHr0GpAzNrfIR6nwF6GL0ytSMUhUYt8nSZWQ/kTNMI
2GcbchGYypssvs6H67Q8tn+7BpGUrn+Whx/mDV6U+J9hfbuFkGTG4S1Wk/sj3gkc
wquwOAlSVWoKEs4yQDGsvQmx6xy2xfxjrDdCCsXMvJcsae+JsBj4ClpcCswZR02C
9LZcvT4wsW3KMMKt9K8iRX9Oli34kH9Y779pTV77V/8HNi/fBUOo8FBuM0d2nzQ1
zeIXD8YdN43vczl5cHmvqHJxIYx7BNQhSCC8PFh4QDJNh2kPU4AXR9ILmWHfVR1X
e3iztRXcEc2QleGZwpcgGqgFQKefqnVcGOT0jjGjanG7lNKTxFqPHt29gxI+a+Q/
PNe3oki3Hzt6mC1uT5oEkbex6MS1pK50xBVnNkY8qpDDNdYMpthCw9HKmiqrboB0
c4ToHZrvn9XHgouz4U4U5iaFqbRhdpRYBdeA/FlUIAxvYdLgfVC01oyHTKbpIhSv
h46CJmCwy4CSbwV9TRkYRH0nIOcWJEbyEuE2ZPWM2TvBKZyq5ol+X7Sc/Sz3JswG
UutAsi2jBJEPlZ5syyGhFfHrMzx90+E/HyrArvl6fbHLMh80OWcJVl4TTtbUCq3b
WsELALgtXAlx01J6iDSapya/bl3ZI55aN20GDRBtVpCrTZztIGX7XubNbps0yUxv
pr7HA2hTb25NXARISEBN0iRCyqGbzvqrxJOPDzIum84e1A2OOCstdiGSNw8+KNzB
5YxBINx6jmI0tEEIspsC0Kz+RKUchSj5IHdpaJyrD62pvmRChb17ODHidhwsEhky
erU9xiyCMg+ebchmK8t9hl6fBsQLwxqlH58M1IBRiQesWvvd3j7iD5qfrx1Okh7O
o3aDad9PfPBHhD+6xo+VjVVigOfgJ3QnlP/ujOEGVQ1gxd7WQ+ZjrFRzEjRraI0M
Uen8ST94i6LhfX+j+qLJgWy8dXwZjDvxk0RPrWdjc114+SvIDSW1FD+x85eFyGn6
ioR8R+GMxvfyC1mBVmo3vR8X7cwvHOBgL4MEbN4lCkbXC9+fFCcmNKH2d4I/BlUA
lHhcXtt8z9fqjs6JcNG2l/wAT+knAXYx7KA/AfQNe77DPjXadQEP2+ThMREnftah
lbHEP3/klXgHcrhFyG1KK0/SbcUtcBB192lFnJb+dCNqx7m12htkqtqT0pgZsl4B
DvDFw4Cg7Sb6sw1XlH6fMVehDp7u1A6U4yX9IQTbQSJTDCE9/FmJgAerCCudmgfX
eSmx2eX0FB7hOnP8ADhXT0Hqlq4oTNFC98QWAVVMM3ods1HE6DXTkPA2B6xs5ck7
Q3O1nC2/i5TqVeaYGkHVdobA4TXmoU0oi3Udkpf5ovjX9LTdG/+vfEDev31F+4kr
81uEUHJZqPdcw540EW2kbBHbJ+HQQaVI0VvjLWZSzVmoIU/hmwHh1u07O2xdL3ni
jTtp+WAkj/Vy5e5296JZZdVQXGJR8kJ3KvrcfflMY/AE0sbhHQ1JGS6opdtzmwsK
lAgpTCr8xtdhlNYnOKRYCA/j9rwKfRNnJr41AWcBYgJ7ooawLdrF9fY4JQIo2UXj
9iDyrtWc1ptAC8dIYK02/g9oNMxb4lJ6+ZDJpnJpV9/N/T1T+KuecuWH/arWqc6W
6675e4U+2qQLj7lgEuGOA3XhOuj50Iu1lErSuEshIwG2NJDTE5QhZb9iMfHaez3E
ZBO0CDyt0qBSFIYSxbUwOQEleL+wovWBYvEwvGf8M2U+8wMW/Qeb70HdkUC1aOAf
ewlDBlEzddvyRP4P50Yw5P4VFiMMjyH1a+24INZLNiw3SJHZLwcLIyBavOU1x0mD
Thh+RK5z8ivlvIFUkRUba4ggpEEPhXwOQrHHhVKXXa9XVV4fW4Ek15uv24p6Xg+z
7C12I/3NgjLDroN+RCGhNqZ2XS6PXiGpNNBS92D13PevIFTpLETV0x+DzoR38Lvu
SOauE0xFK9RCrR9gHEFYUh8KYbcC670L3TBVgEAS1HKWSOYpYoKZWwsqcNEDsMwk
OJ+cCR+aah0l25hX5P1TmOlNueRqAHIPCMOSSEnvT5jW0zEmjJEhv0wwbeplnPDE
cv1HXrK8/5Mz5eWacNGbWJx/aPr7Mqzh+jtV0UMLPxt+KBEsdYfQUU/KGA91qoh5
33V9CGBV3ODaKhIc8Gyr2CNUSB6DpcWhpNmegsDVp77WW72Ho8qR2gVSaqYA5cok
85w52QlEgakua1rC/jEvXV6Dp7Xq1jf4h8d5wJap22lKZz/PwCuRaP7vL+2pdPH6
pIKH3wFQsuKhoB4coptRSAy45dTC5ZP0XoWRyl+Ul3ZDt9gjr/LPrYLXwFjJzduQ
qvOlF5SQ7hvgW2Zhaap4zLCZesdFs1FB8KHTaWOD7Ogg+CwDWw9UwX9Kbt1NyXxX
plcpixnznigkizWf/W437s8tk7j6qjLRp7gn5L0xHpQFtR71HraXL6LDdTPN7BvL
JEju0PAS49qXoTWSb4s2acWhfk1jznpqrLoQicwIQojo8lBWGYShg+t0Kbp+jbDu
owxQuMtHQfEX3sGMx2BZzRaVKIF2db4k7Gu67knwuOTGGlIFsAbzIg2dQp89h2+S
OJxyVfYo0SAc8zEBX9lw44kPOcBMtkfU4O8Hf+7+F7IjLZNIo7XIIMU/oAxQoNyF
4KYfZqz5w0eTBmDmGKqeGFdZcjbrzuv7n4WpswPQFjGeryVKuPsOuP3JBn1TPWSW
Vv+FunrcQEdDOSOMV+FJBa/rLatj8F2lb+iD6yhyLM6GS66pK2ZdQGW4ff1M6yaA
RfKff2ne3ZLbkSF2SBFZV09Miu+g8enqC2qkRbd48ITRZGBFCaPTXzqaoBrSTbsa
JkoO60jvoumcxnwUnWqJAm76kMUMZiZVuBNiqnMs5ZwF32QOawGVrUnb7iWuUd3C
ivt+dKxwmOzouNWG4vlmnsVjeF1phUvp4EaMwaplCa/SHOfTBcHmcCOhdqDI3tgh
f8nCl5wugB9vplSf9QmpbbLtqy+bGpoJLOrFreq2aTQvPLk569yZ/FNFx5ifrpQX
WL/Cs/Cr1hpoWHO5nJUs3rURp2rg1f40hlVJkwdbVF//S62pRzs57ZE81MGrerrS
dM9wxi4HWyo4uwL+xkfvrO0LujlkXDzQMI9iG/oqeifMbm16pzPjj8geUPcq/Fbx
ZHcXle+wj8UjdBceCbLxbrMUvw31DMfQDLBKEnhIc6NkFx/RGfd15KYTjQolCene
KkqPBJAbBeF7S8pat1S76Rfi/RoPWpW9MaqdvTEzU8a87t8QMS3CxcXrCmN76FrE
+1jz2ZJ8h8Vdj+8limWAnR6IKJZhX2djYYSoe4XBejBniXuVrPpICFaT9etrcaY1
bCPak9Wda0RSYODwnNyv+uSXB76/nr1/CVlI+kk+B0BsXGGTiFQF1wJw9bLRrKei
RJvngymvRjEY5QEaBDQzFdb2KUK6/RxO0nwbjZIp8N6t31DFkT3YsV1oDWyRTKV1
MFNJDlgXGwbRLAXqjjXpbnt0pbn+wd/yovrmxvB33q7CWhrz2UPwAQHrRsmC/92a
dTC7e2exJtIOw4cJwJKjOfBxGBLA41wi0OFFvdL0KCB0XeWKbstBVgc4lpSf3FAb
ZajF6vkKX6IJuaNfyGY6/8Ir7cPaO7Z6t/GezQYTdwyHkE+ZjugJotB63Xl8Jqdi
6Yud4HNXUB71BAaHzg4WShyrup8pdvBbM8vt7+pab66d3wPPdo66KcK6sLNbM0jH
OG0cGM6OCLMC5lf8LbUcfgAQHAhEsa1RclAGVtlCbngLcsIl+HTnaTNeH4VhlWTt
jdWJqbbI42653p8yOzG7G94fKS2lNEIUlrb3xuj3tS39h3GZVQDrYuRvmle71WLU
zaCsPOlTMGoVS0XLsyxB6p3cqgQ3/YxWmdmo7BXdm6C+/3o06HY4erhuuqckXVNW
N9lZepqbtUxAOUwqLzBF9QSIfan8vfKrRMARASUk4BmQnm7KrHZ8ppr/xQ8qveJ0
kQYqyq+yM/i8KyD1A3iBucOzi/wC2Mh1nmHQGCy8r3Llfn41GEGBbGAndYaWkY65
F6BIt2KapHGB25Zs1HuCrzBOxGArtuIL900dipdBxQJbLluqf+ePdiXxwCse8VmX
5jggZbclVNtqV74QPFzYE07yQ1r0tVEGymcl899ZNPbMRJ39EDsXivVS4yrNeB6G
RMZRA/VQkKPgDZBj/IaRETIRXjTOVglhwitI+lZ1ztOnZmllMpNOxMtztADtCYN1
RCJEs80tEGIYKoMbTvguPmIkn05/+il6JYfnlGkva3hYiHmrkFjIoKVbAWOeisw8
wTULivqWYImDW91SFbjgJHm3QyhC05DHZkuh4QO0fNeYwJcDiMuDsmlGIc4JJFEz
mSfLl3JrdEES5h4os/NeLLrSyUtK7bPe0DRIrGQxRHmBJeVBp1mCAwJlM38L4RU2
33swE59PqdzWGBKO9Ula9pVbgGmNx8929AfqjQJXhA9iBUtig0K/7omDvzgYzest
W1BeKRn+uod38O+I+ZNcdYiL9m3OlZbJZe0DNiWa8rCG+n1iBZUAUGZWfcW3ky9m
wGiSJb6A9tOIAkgwUPdD/GxZlDi1Fg2pHADD6e0KLFxukNhxdPDXh3NuAShNO2GX
otOLL0Kb3TQ9uGrImW6VuwLlnevWBeuralVxUhHvjyiNe7uX/rBe0n82UwLmd9yf
3UfPGhkJ9jkTuf7R8NEhqcrG6whBJJ4eMNHxjMILZPmshpdcVJqyDIWHx3OTrqFu
Bvmtz9YxLboR+LYNsm+XpJO5+qd2M4lqROI4VXQkQxxJUAWsTrmqFN1vKe6NFwBb
4ln0Zmymv9jXEQzz4xXyWR/fWZt8eA+AplEK/qYSj7DRx/xInnMeZ/SmHlXjXjUG
yGePRlXkmMWX42YnMtm6dNn8EYo80MiVHkAtINRLMTAGsqkAfqelnMBgcFRjugHl
qrUt3CcBy+uxlDQPNy8Dg2N6JtqVbCMciaSAHys9th3WS11XzEpKRbkMFJlsiUkh
1sMS3m8nXtOyV28z/P1L3Gnl+IrONpEScDAxvA7hDOk2wMufHHLr0Fr52+fHggHp
n1VMVHZnMj6EBNQTP5pAzYNfNVy57GRKkpGsFYVlLV08T/jR6hD61H7z5e9I1PbI
pmyoCf3pcqzUW6i+RI9h5BGgug9DisaJkzpf4Mg0Thtlm536sHZBI+7KEUH9GSdK
GHZFWkRA3RRAMW7jcaYdtCBuCy9kohFmuuGI0xkdPyQb5Or2q4eHb9hJ8lKRhUvz
7a+dsj03etpEDJJfngJmqCv9C1Jwle44brPts4dD/fMFvADIN/IPRYoKRy5AMVgi
qbn1N5i+06P2VE3HrXxk5UiUHOzG8UYSr+0Nf8FU58hofpxL8S4C2ZLRglsi2gNq
lOJjo3S5oOcmbgaoYj9fMCGf9ODUGh+D8lIOmFmKopdzMaCt8Y+DjB5DjoM7t14h
c4L9PxL0KPVOY140VJqhkRNRN8VY6k18hdQeRJ9llgVtI85ezZwYlhipGOjRh4gQ
D0WxRhONoU+t+Sn5mwshCmjmdGsH1lR4E2cOUvE6FVEuDoc6rO2BuN5svgCFEaOs
rIHSKPnqFVSbdp8uY6tJUXJl/vurUppYqt9HaI3SICymO3uKQ9ktX/aF+pKo16eP
PgHQaxO4ex+r/sFAMAzQUignLFHXyVSlZtjBwKJnoW0H4CIxlKnY52yTjH6cQgFE
A8P6bx6lWFsn8qsoeTGaS0uXGsONkrX1JmCW5PGM5r+SQxyIJx7bzORUpoKKfstq
YCTzCJ5TLsjXoi85kR0bCqLbO7I0Cw/KlXIH7xMG5lc1YMpc7Xoh0wU6N+dCYo1c
dJheimQuDqWilH8cgrbFhZRbZ9FHZdlH9xkG7AmF7MG0buRUHfFxnFUEt150pNho
GS8G6ndZc4RL0nRhaFx6lV2JybBpFFiXw2UGcM782LwEnunstKYvxjzc0VdQk306
lWWFGAnET00Q4DXFiuflKF2H1GIAQ0y6OtlMw/cTCjYxR6d4sRCj+UNXxez/KU25
cKats0WBr0YPJA/jzAaIGFy2K0YPL58FuFTi+hQxPAzRlXvNcMTDzp/nvTzYfHbM
3a7gz1bWbwljgkoZBMBaFfkn4GKJszW/xY0bhJcy8elscULPjbQMpUzoamJGlH3P
gN4D0ThwFzwXz7zWuQhe2JZ4LSZ3DVa+SbONq6AZXJY/uyegY1+Tkh0RHFSZKuZl
RysntmpQYVFmsY2iQOLfHU1UCO+RgnKSFU6lPUk9tkFmDnmyYN/FmGqtwuM37XSy
gMpyTMk8zVJ/0bosDVaTzitZgPPqpfSymE+gDJ2lscuODsoE6zAbmoQRbeuwqVbZ
fzPA+zcdkL4GECmJrptHyw9y1gE1B1KiCDIm+onuUzEucrqbMoNq7t3QFiHEL+8A
S9c3mStYLJa4USddL5xaFutPKkMtn9oJ90kujYRl+5yONDL8kCq9r1S93TjqFbHB
h/xQENUm1SSQIZFvurRclSyKLoD2WoONnvoMngJKVQvEWgI0WQOoT4vU42B/3aSC
jRc9uFEJa4HhpiDYZriRtqsiOJPW2670Rhn61rjfAeC7eDhH28nftnmDGbOo9klx
P92F6xkjXLocoi3y8AkJ4h1PKalrM7K7nC0Dj0jeodI1S9N+pqbmM4Z2zuIJ1PMw
xtqiJGOTf7TIlwZzhGlCzm7x9HclOVLBqXJBwg0k9zClbCd0f8Y3AWGoapQZ2gK2
q/WLuhjLzwTFsLIpdvGJCnxw5+3u/ILbz01uhvYJ8aRYfBQODMN/i3aUhq6f4P0g
S1kAJd/ZTv8b0o72eTYwnZL4sTRIAfiubrhzztFFLb6/XOP4ESAJ9fyKWgCduT61
1PKVD2cKqJY6yJ/QYjnur4SqEDcXBhOO834hXcsveu4sb3Ftjr9sYgqcZPDUsu+D
gIuC9wYdECvFvUgECq5GaoYX5QnP0UofRyjmyGzTpXsKd4tNHdPn9wXiamBm9Lpe
lXrwRpEawJVUUff9FRfKqKrz6/UVNNGOxBUPLCmjI3avS6uJ7LhNeiN98Tl5WHYK
2wEepk7ivMfCRuUjeQCvNueSj+MbSGPI4H6c6kNsJekfaVce4Z4WJmPnjJM/d5Oc
nQG16aynMwgmAUx4ht1D9Sd+esrYCEQJtKqVaGmMl2Goc47ryB7HaOP3kFQhJtsZ
ODu11jkcSAF15gXarna/S3VvV6FztGZXKvZ91+h+yegMUTIxXzCe5PYeknUGbY36
o6Cjb83Hg34YpA/IBa++Gji3yz7fr1rQElIvdjdtsfwNPQ03UiGaxXomL21c745+
GmSrrkMehPOxdMwm5WxR6GJYl4IT6+W1u5SGBEeGRDNEKWJFOsV5DAyu8l7FK4bD
7k9nonxGgZCS5o48eC08J67PWEN6XuaZhrOhGvz/bHYLKXwfV3jsSpdST++kT4ah
omiIeyt7tDvAJazmN+MCuOGTPaWdlSETq2gbrJNpRJ4FAhx+F/hxUKb+rHBz6o8K
dIk897clQtbGnLX4PC7zR46MXnzuQGiIvG0NmqvuOYf7WNNeXv7YCyY/MGAxkLNq
PuQSDRnHU5w0u7M8q/SUEolp5eWituBxzNfi+H/jiIitl+tE4kYr/WJSMgbrTW24
DKBBWJpW2F14nb/X4pPyJI9VuQxgV+W/lP0csrGx3wTpr+s6XX4K5lPMeKNjSEoR
ShJU9T0Xen+dJ9zW1FqIyjHRNXkgYAqnuSiM09+DzNVyqRw5iZSD2t+CmYknJibB
hoNBlMTadT/chzy/oHy87mqQKyrKx1eBI1dpLvEirgzGNf0ioYqJ2LNjvyApBMlv
Zy1sTo8ZsB1erk77xzMr5TIecgQMGNp24kMTbbtRsJs1pPeNY0RwoEgq5T9/7YZq
hroYKQpKxL9XHyzu3+wc8gl6oydbIpryfv3gzsxfbRwR/5pGkyHk7F/kyJfMfVCm
arfMF5jxX3lT8CTdCCvZZ0p1Yloq6fNifXc2IrLDbd5jj1DUqA01fPQjqRwVxmDH
jrtZnbubqcLiltz8WsepHAax6+DNInvOYvQy6kFofhpBCUqBpvxLm/v72NmqBhlB
+vCsqks7Nps4OIKfzATfp5q8VNXzcnZCeYFpOhb9T6aEvFuAJfikdNsc26Jb9f39
FwZuZPcGCM3mbSlPDcfdP7EKBq6ShUPQG75+PY9N0m1eYthJxOuuj6JExU2rKXA7
wXSpskzMDEZtBp7i1eO7Dde1mSPeHcpJbb41dIjfnTCJoGJEewRMoSMUaWQ4DD1w
x8OwouoEB3Z20h2ODLODocqDx4aGsqVMYqup0IIQznudxW5e7ys0bVD/jz/bXKzJ
Gg6TsIYD7RtHbBrc6xyQDXt4vygJ5MnecG4O5QepulIhojWn/w2C/61RVg0RLzyP
VipQNVuA4UJsNq0RExXWVhGYp/E70S51mZblme8uA/vpJNWRwSr1oufjWJrsKXba
9QWkkg7K5M59iRbyHQxbjjoCDvdiintIb8lc72GpCdfeEM7WtKRODmk1dc3jH42u
/HXUCmzZTj5tbydiQG4qhY+VNOmagaNZXkjY9zIUP01RkqFfAOktEu3ANfyhpd1c
BcF2Fts0vP19TTTbpR56vqqE7wPi+8+86UfNstsfNBx0U4jA6o3A1uUAggZqV3fC
Js+eTQa+08syOVCQJjUJLwfqDSK4dgJjO0cy5yfb3gO4MQW1VYC5ptSMUQGlMsRT
81RunWFBjwwm4kGXWz1aUjYSVunE11ENLSxPQXaiGAhz8Xu+Y7oR6R59WBYveiRW
9oDbRwVzKFV/LGuqPyntcPoL4wkDld6rXuDCFjbtA1CZllo81DwArRkgSYlwnRol
Yi0BhVOY4MRL6usGZ5eLqV0lxK04x2riVT3MaY4E50XbnoVopwVOnsIkV9Dgw2ua
GUg1++QTXSMm1IlUR3HbXvIduQOScwyqYAE39YRkYMTxU/I09aVsSe5QjqndommW
2TWBGNNzfCA+Ztd2BQVfUkLsglKHxhkY0Lop4ZrsGLpUmjKClUe59VzDYQg/DAmx
7Bn2MLys+Q1gw6El8kKL6Xq4+hz0ctMDWBn6HzrEaYkIDPXpSW6yeDfIndqj9sjl
2FMM5YpSe9wmglbQPNd+lhlR0g/d7SKFMGr/DDFoerXOOHzZD8dfxjnhVkcxzVLS
2EA7jtiAdYbXQEKrQSfx8EBFKasSgj+RDj8T4/n+1UsA0xsHGUexiDMWJPJtlGFY
Xky0K1d7uIMk1PS4ljI4ML7P8vws1HKgNCHFHLCnDL3ZjJBWJMsue6b7eB7J5yaZ
IS8KSey/RBEO1T5KtpW24qqYOlCaY3n/1Ricg7Dfhpbmqxh3iQXobH+ISyC//Asx
qJv0SjT2xAkwQpc+w5J//VkZte7ak/jQTJY/G7sKbSRmwSXTTSrZFa/RR8xe7QMo
8B/+HPqYBmxMR4Az/K9riM6+81BOmxxoRW8Vt30rfT5uQhr1vDjxhid4WQ2qLWzb
RlIYp5QybPKC+yo+QlrumYOGx0HBcRV9SMPhty/GHE5bcr9bnTi+1EEHBYXY1hx2
W3qwF0GbbyXKnuCYIsPyZ3rkcaP1aVKi4/gwv56C6i5dWdsWrCw1S8r67rU1cxZf
H9hxpPfjzUPmi46mjWRvZ2hqXjJ2rzCaHEXqBt+zaQwN/3kY+PfWO2YGgxb0wXny
U7pwMQoe/HCdN7PgdVs6leR3cB2+8BBRUbb8JWCvCNmFnjImKESROVkKSUkFV2BQ
moqFb5WP0/yIm6DWL3N92Lhs3ls9vjaXEzl/tYdW7C1WHIj817nRy4c+KUiVvG6m
VDSWTYtHB8pDmZ+sHp1ljY/Q+kiKjJU/cSCS1vm0Lca315pLrcHivmmu5/WGNvpP
PjXwPCE3gv/YUWQwjG7uGZ79T3H7N61IIUskThh7BRC4SdWQDCkXKuwHc4ykQl+b
x+erz7Al0xrikQGODl0xC8eeeQG6OwpV14fEIibuqfVlqU1AoVQ15bzoVEqr8t+Z
a+hv+psM0RK4RXeaIDaDtMN9r5JubK2PDXc6ENwZJZTVGfHoHE2JAlljp2u3u5FC
uJc9NHtm0eyl53Jfb3FS3DqBPyEGred1+mREXh7imj8TMTZJwwHwiYFN0nfQZot0
k/pA0kNX2PFn1FDLS/GMLONCAQSwEBo/ohxiniDAaKbtZMyZbqA8YR86+rW7+V68
E8Wjk585DUHpKNLek/ch6eog8MBzlcXEvK1dXPBVddmIyroWvWQikFfAgpo1uDLj
uV9gyE9khxHJ7BSM3U2LwEEvorB1cWK7hnZUdgdmnDqAgcVPJXsYWRMTszNO3A1/
PBmyp/2oRh1X4aG/HE2bUk8iqtkUBN4FKUg2MIHDH0YWqo7/WkcTF4/tE12d4HDi
i3biYScd7zSDR+HY7PpDDJjhJZ+RavN+lLbpuvGvyCNKmgoJCNEY7sH7qA+AnuTi
YwbzdWG/PH5qK4+DlYAxWYWyvvZjXsdM6HuIhZZm5oPFsDkdUo+JkixAaKBK4YHZ
s38jdefG1JNdZgCQ58zz2oXHi4xeMP5k0GO9kwaFnxBYSvYZMhIDRY0uxRTQe8PC
ys8BQ8FjWvZdqlIOZWvpGeDJgPcKlYUknDi9XA7pwwwbF/6j9RtLVJwpxDnlT+KH
roHwu9FI/+jdDJMJs8j+N7haP8MgBqG/uvRgmrFafHeH9NHxtpQZk2U4STVreRJu
I/JE5olSh5XRPwL3WO8tcRUVWaDF+rTM2eeunB2FOnj64P3seYfx607n6Mpy43zS
Mzn5g6hIRrS64YixsXtJ5yuHmFRdH9gOiybKG96O2Qnpyb9xIsEWQI0xHDzXn478
RRdv8/M2q7gsvsOaiyqUzNU8BSrRh6kaCYokS7Fnkz13EJZMm5pSE5LbLSCWU5DI
OvZvF/T2OPfhnziwxRvvoAdNRRtAtoKczELehCRwqVPdsiF5UWjr/fXgkAxRZRrQ
Eu0IrR3xQNkY2HzYjqhJWNipEUA/EaCQli6s9mui6kbdO0a15Zk+l53hin6Xg3h+
EXuVPBWvvO8ssdF5an8Gsnx3xKAxN4HYq4rlNlOGW05NgKbyM7ijpKzQu8qwEDnJ
UONv9cUFMe0Jn2AgagKUd3dlpQq7u0GE0d4LaaBZ/YXBufFLnv8p3Un6eNh0Bqjp
BsQk3fZOZIleE4MChn/XORx/i/gECCcnvFTPTNZgnlUnO1PUBOKNtzrWhFvsC0uu
zYVdlM8t0aVB8HPgeg45R+riWveTy57bnPQ3YGc4/mm3CU9zjd9iIYXETiHIelaG
gwyGAxaG7bBzGqkgwcIzpAeAAOZL3hdtdcbBw2rmEjowKdRUJb/e7/+wZK8Vc7Lz
DfuSaMPQtAZvTo1BMQg7BVFZMKdhi4+ny8BSFEZzfLkY9+UlBg9pbpLuvFVBWx0U
EaFx0tpM5x72S3w4Z7ymLP60nr1fO7L/SmnCdh8CLzPoJbL36ng/T9AHektcordl
+pus3iBx/bIQl88Z4L8xSPVD9NqvLBFepFKUzHK5lS6y4xOB7ePkBuUlsM1qDqxN
7hrU7uh95+piMpTN7Cpx/xdHZZEi0YJ5KmHL5poTwLVIWfALdFlhtjdOpEFEAyQB
yFLWonYdKJ2vNdFUj42bAOaUKCWGVQu/zvOzLiP6e2Po/wucSsi/Hcn9DqFOE6hN
mBQpQNB+Nxe1kOsqS0zkUEdD7ua1iEuOe3Q5v5oxtAx3EZK0sD+LTFIpyg0NzUIW
ILORyXy47P4nKf7JK12btQFZxxEGUliekqYsuFF+2xpg0do83a2Wk7GrEgfjSt24
6OJw0BBl5+bIN43Lz2U3MHEFsixePSCRugb8K7gV3yGy+J92LOxS88Ac614HRbvr
avKrWqqWlI3IcnRHgSpqEAlfc+DtXgZH4XYdD0gReivbsIH05qm3x+stngbg1BN2
LmSXQrJsrQxVM2SklBTShmrfc4mkGB6rroFuUEpFCmHXl0CBza/dEBCOzKeD7s4b
VdtZ2f3QJuWOeft0kO+zBKHtD0N6Lv1wxwkZxn/mHq/67shWXWsaMxElEGpBq5/H
rZMZ682Pr+BzPLu6s/4Us/X2eZ1t6uh7mcRBEvIu7sGbb/65QwoiE8jrO8Y8ZZVS
Iy0wh6NuL3+BF9oLejpQe8J9ZmDP5zblh+R+GV/IQaig8RUuoaCTkC7rh92OnDzY
fn7+wkWy6qPMNWcm5sM6kwqI10N0ews8RFWolRiaYlWDmoixAPLVJjAERZND9x/p
zU29mRhvzRysHZLZ+HqO1Euw8IhcJc83lJMk01KojtfDH8VmFId3JQSootUXVpzL
P/eQVeUXnaZC/2/NvtLEotnpxvRJml138AXP77H8zSp37rneDUEAngt67oQJr/Cm
5LU8Pxy6p+/T3cAPZmWAmQWkKRiCXLDJ1iCVy93RfbWMOnH9nYegSyIHej3tsESm
CsK3YYmQofcCg3mthRgmYLfDPKx91mDH0BMPaBMuTc+439dM3eWjQZvUPIL86dAe
tCFfCodDJz6QcAuY12EpdYk+9+7WnTNYq74RYTcp1/EmaN0GZ2QYhVopcBxbGn+H
xeDGo3gcJ9YWiSOvxrPYlvVYGgxxVJEc592dKImEVB2JZg25dKNI0yelMeh0ithJ
TGGFMw65hn0aHiw7EsZe1g4DiroN+M0BrRkq55z/C4rIP/z5KpnGWcM4Y95/y0ZO
7MFL/wVSQIpOjor6Spx3o0pdaDhD//bHJCgupXhE2blHKBdGNYBReqkA3QactoqR
vi8387OCuCruvC6Mib6NmGSGc/GF2bPmGiLQJD09ZJdNdMl5vVmXvd6+Y300WyM6
DXHwpBiQw1aTENQrqfQPycAPztiSHhX4bMb7rQI1bvv6QWK5eNPbbDK+Lv53Nbcn
7XKDTeeHNIUMjLEHkdjdJnAcnjqdxW5KeEjp91JJdfwtcGfvm8MlT1NEZLaag0FN
0lki+ghABWjWwQR+IAy1CodLgnqV2LHi+DzSQnQbF6l0jGKlwi6DgNG8ytYCG+HJ
Ua+Eb4jeMZ1AsyLLxVLtgHa0lj35jnSvwTkGRX46n2e69JD0SXyNBCaI70zpmArV
hW0+N6E4d1z9CdZb3vJVLs8W8JWPk46DdFsFpIynEGwdVTpH2wGR/QWJJDRQqgBL
0MIBwSOjDsAa/EDzldbHdclsyF6OMoHZCpCXRiYvib98JbroJQmicRT91OkEDrfU
u0dZiBC7ofX4ZiMwONElFPA4KVRovyWAhfZvI6t9wHdWIOcbsgcDxM644OWCmfF+
NzNftb9Hqz5o4sp6wBXJTiYpJb/prDcGoculC2zsEe6YpQg1acDlHN9GPKVrUpXu
LnKbegPsSyE0o1UVJUxEt6IRuN/kUujF1DUlrYpeaTfDzA4Vv8+bOSkhsdBBXt6y
hK9kTbrsPvmj9qeQpty+nzi6OW+ATVQh+immTxtxjJ7+RvkargCtJwY6Umn9SET8
43CUIuwLpoYtigppZkvEsBZ1fSn9dkhT8Ee4ytGUEe+jru/dPPgD5c7lMxq59XUh
cNYc9fss4xqo/0zIe/fkQW/t5ht+HRNEBmRSd3eXMduj+ukEkQGkAezo/pYCnwj0
Bz2epp59xbRZj8te5CEL4UZZPIXerUuP33rqwEhHt90Jo8QJar5oyr0INqjOqKNo
aTfil11J6nUrN2Z+tET6QqKwqqqH8ynBGRcyWdsMKGuDpBmGrRhOyLMiQ/zgMBuK
sSevyy0UB7Q47SUumw/+O0bIHLa6miGE33LOWjxwAQomBV+Ybuxj4ZVCHYC8iQR3
IOVsWoSUmm9FYkdVDnbfh2kQrYp6vAyUpKJs59Z6iFEdpkNY2V63xO+3hkfQft47
NF+mBX/VwwQZJ81dXYc3KV1UpczaJyETwcOSKurxfgoKcCZmSRfcIENSdZ81hrGW
VD1R4e0vHzgIy5MS0xR6eKOkJ3ztW9e13O7D0bsdmQsv6HF5VX3yC1oZ7GjiNpgz
RzQye+OTRxEToZiN39tYGevPMTDyfml6crzUund9OfP/2A8tYwhOINc+9mFyVqQB
dd+pBHk5bbflRZ83N1H/DM5W36jfwwAUVCeoay5OEQyppXRcDhWLJvU72Smt0DDN
HfSR7YH0LD4XjwwKTfi7F09dfRlIX8SmYyOWsyAYIqR256SyUWg5KhKpO7hXFfcb
yYgJ8AXKlnTO9NHMJbjNxlGDRNYKpcEqtK587o1rujkmGuTzhJsqqqGKGF8uMugJ
/9xUtExcZsI0b3RWoCa3kfpXwk3dkaG8gHLWIfYih4ODX2CGDafH0sDVbPqZGa4Z
LBAUC24xX+vbDKzt5z1D+unS6Zzbjgzhc5zdh4b4IZ104kgSHstnkUqdJhb6Rbl5
gWyzmONOf+zyg6lBcpD8Lt6wP3c+ccT0S2uPk6zrDNopcsSTt5wVVIYKHG+c+raO
PRmNIi9Ux3KtmAHpr4YhGVID0ZV2SK/VoZcD1kJA/s59c/aREXeFcLP0Wxl5febF
RiY3jR8su1c2rCY0+PgBdlG3tRJQ127geioS8gX3jydYGi1z25WMfrG6HmJb+9G8
b8gkZpHphBSwx+JlSIErYy5x2YIPUTLCP9ORlx3i0eeGZAAHRS8yLreelRihdnaM
qlOx007NSTXDR8fdVtMBeCH0rdjs9DvM8EuMkypJmTEM6IxikKLdtoMlWNxLEp0Q
lle7XTjEJkqtnSC+8WnIYV+5K96JBT4tSF5xAnNVGfkORLEeAXmcKbzYqZ8goPYz
j5El0xqCt2Ik8NmYsBemkaiNRxyjtksGNu1HR5M2hFxwS286vKDqGJNZq3qgYwXm
OflGdzKPFXg+U3mFiv+oaY6Aqd4Kc8ViHrlnAuPZh6h+YoSbzSmhpcBnlqbJ+W3o
Vbrq/EopR47m6zZDETs7ues6Mojm5TUWYsWuvg0dMts4O8aVx8WH+Qh7x2/98car
6t/OFPtwNUUEsnjQa6ZAViAqwM0EtNP+7vUqlHQoyhhH3mCovcetgfiHJLJQ+wCx
UEKiaB2fkg+vS5aYFsI4D+z0igskhpapt8b3PHhobMCzc3/HxTNEe/hdB+CPPR/s
OwkxmAngfjfhHVjwQWtq3atzf55LCflFBRwo3DwcS7GX8KKeP4yRa1NHCGD/U6pb
er+o+Ytgk/TjZCkDqZguSlTl+ScaOw7xltBNwbnzsQS3GPMvJGVf/WO45gaSAHJn
6+CVJUq3rCA9z+uunMdzgdNGlyvK/InduPskALEqvh/0YipxR5abuvZ51/+sbZoR
yOzXymA8BB/d1oM+lQG+0Mf4vfE6Qlfsi0XQSSMsN8NRkPc0ZMnSuYl4gRI4SDM2
K9xQtqQt9u4xKSUvT80nW3NaTKTgMvrtaXD/V1kTi50vym8LmiKcpTP3xdeEbfC/
Zqho82a6h/gJXMMbzcgb4+kaxXNmNgHzdZ98VbpVvKlp0W2fGWqho8kftOjkG9La
j764B/w2i8tYudo4ouxA19glnxJQ30HMzyQQZkNO6KHMfn6gvdPccqFhl9bHT4or
G8CiGIXc03tOTPBfIqTLL4NYTR5ljv8lAijluK9GXaRb1XFfOi8BN+dBtGis3z2b
WWMBHn39AoroUXHiaRK/Y2F9+1tJXz0uFbX8TQxyA2awECgQ8XvIWrT9SBPWXVTa
s1aYjapu6cBAURMpziing63ZrEkFjon2SeYL+rupW28VM3+MJZj+WXq2he3D5L0s
69PnYQXPJjRtaRXr+iFREE3ruSAwRyF0EJJGe0MHytqzZtQ5Dl1BsXObD1fnZVl+
uroHdu+0zymfga/IZMFKEafG77wuy6cvIeW4PpfCElR9AaOejZ2glf91VGg+mA2D
qVyCdZTUNxtvXwgkS2MR2hqyaFPTM4EBT1JuBiry3KO2RYQQWjmicv0VKcra+Xdf
oS5pV7J1Ln+NfwdPoRogds+TiOhZ8RXA5zx6+y/jKnX+nd0A34Xi6bQAfWAPJU5z
CKduDkSPkGJJWZkoW2lYBpTBM/eg3Y5hXTNPusTPOTqFGZwQOpvaqQAnLUJ8Gfx7
BJQ/WkmrCK1AVwzAvGAgIwO0oWc9m3QfiEhyFnOQAnk1QnZbLRAaDVkQIvYiWe86
FthbAu453pGo8ll666zERgjrDApm2bcM8xa9XT9RqIyc5KzXnW9rR3VvxCwGdpWt
C2NH+63XYOPUQNM6pMB3iSRxWddTPbGhusgYItfjqrGXQj1RdAjuxuo/tRXkfP33
327yZncsfGYeGVgTj4h6slZR8x2sSwdAVIbEWHO+3SdXS4Cqvx+XJK3NIxlMI/sD
SjfpGSdmKtiy1N25z9y/CLZ010t5mgfexWBPISDp2CsBg1hiq+O6Gldp4qFbb+zR
noAe6Ne1ZbALBIhBYYOTyqwidkR6KNM6PKQ0qV98Y0590kTK/QgyePhufgvK/hMc
68QWBZABAq8EMSu41gpnFyb5+l9p944CBNysvy6h/Zph9CB0U9vpGqJ+X9yQHgiq
KjsCrcmKhFB2kPj87xzeYhFSyKe6gS2hjI2pgK2RUi+k1V3bG4CINrTcwoXStlji
aYlIWJSk1v6EYPEO8VIhB223Lq/HnemDeCfhP0tdZo7kI9lfTPk1GCWPG01N3vhn
5z3djRQMVim77za6GtOUv3lIiJsLNQ/p0DUv5m/1B427loUY2t9uW4ZszhO4PQeS
kwvpxTjs1d9hOe7ZXYt9NfHxMGN2Og45SQSpp374YrI5zoVpDHh3Dv/yh9yyaeSI
CAEFAzCJNIhB44uD5xynYrnzgcXWzeHMfRmnJ+g7PwLHLh6KKBRRKXVMvP1HQTLz
05r6sGdPGNisSjvWJOyTdTS7BAZu7W4162PwhJ8IqONcXWARoRosywSuaI1axjBS
8cGoxWfOwWXm+B5vBX4i7SdWlMSW/brwTBT/u4s108trmiU42fkma09XOuw3aWOA
euaDEzCdCiyH50lLbP0Fg4QAXUlWXLLmd2fDAvVlMuBI9Ho3zUbkT4asjjyxA5tj
fjmsTKbGOdYXKYips07IENz1oI/LHfIhcmVe74TmtzQgoYNW2VTsWUoAlggm5HbV
lV8KYg+BfAJlPHLDlWEW9RJ4NuQm/ru9yUvJsgQ+g0FXLna0vQEJYTHK89pC20fl
8qtJa5BHf3hrd/gzsPDCGTphmRGC8WPV/Bs3Mk3w/8bUen1bynaNcr0xt4vE5VyU
6UvLfR+dgUDJFuISKNXIl3JYYiDwK1zwse7KFTCcJ2q4aLHlpXB3v3nMUJvqNP01
3bQjBeFQKHVwb30l9PNQSO7sWHbpzTArO15IBH7vlHVgcGEW34KJ2S6HbS/JnkAD
apwIxkgslwxPt4a5ShlQYPaMpRs43O5m2RPTMLrWey7mGGGaqtJQOd+R5tZc4BQi
6+fT5mh+wfYXwvZleas+Z7BaIGO50uPy4EbL0cuKp4n9WU4S6usaUoDVRW6XHBQW
jKjy1rOafOlpfz69ab6qQZF32m5cY2XEMu6daSdvoNQnOws0MhYZp5VK3RBS7eM5
iIA7GvxGdJPXefiqNiWxYuAywRBKqiOcYB0FAfWvY1pFJH+zMZ+dGlZXvpWYkvLr
FftzsQ0xuyg5jOeIrY2pDswHNsO/SV84ACq0FSq+lcpjmT+zzxWW9Vmdxf8wjKtG
ogGFnyKS1Bmmc4VNhp43bWZBvmQX8Dezf2CoEhK1o8JST5iQNLQg9LfqRcZu6O1J
P2qCLuC5Sb4Dvrv1o9XFMzqSDcxUvCXKUz9JU8wdApTdBF/Zj4hdfuoMmCB7UMSQ
BnP2flfW/7QADfLd0Up+HfO4NIBlE8bQQKpY64omlKj+VDWcDW2qQ6JC93slJ20d
Il0/dtY3jnH4Rrr6ATndJ9JYv/OegGwPyXQvm2gAgTm5n7jCmIMVyrlaP2/M4cIE
9bbAgYfwwT28bztAyI9ZyZAg7hUs08MRzRnTbmIrM5MIot2n0dlahEI7kFKrNMWQ
Vwd8CmJ9WI8acBrnc0QZaPVOZ8ckzULzJCM8I3B8KfLTlZwpNUMztRfbSXD50BLP
O0MNnriei/GGmVf7WAt9jmVlkub9IQibr1zmZ2l3ZZxm2eDC1ybLvbhYNi6dHFj+
hnyoaEzac1xfxDmmb6wdSySEjIyCyoHaJttrNEMs4F61Sb+FQoRXhKSFQJQ3QD5E
VD8p07PYXXI6G4u88cBPOazyALzpJDghBGZLcWydzjJleZW4Gnrffm+GCPZs4pYO
MJy385JnJLf4E5t7GT+VFMVimhel+CvTF0YWjKRW1LwmxCcvUM9wvl34PX8kTMhN
v9OVGKys8IDWGsOADG8JeRoMfld3yDj3IHVjDkyoxCKIE1JjT/lNLmafLauV6lay
DOfTcp018LCLvDnOe8ceROyVtd3hqRQ1uPXsbkcJdCTamMSaGTxY6B7qaMaj6hW6
ZddoWpQd/hJ6vW1Uiot/BejnDONN8ZtvpTxZsZ23vikGEK21xm6QszIC+KsSzTkN
dCGD7lbfK21vvxQKvVHx0IKXKdVNRXEYYlqHMMj9AWALCifF8Q2P+Bt9IvXsJr4k
SnCWlhh6DkMzMlSlyZSS3I5Rp4u0J8ff4hGJ+tERNZkUItbaE2das7ixFNkP4QmH
P0+GtHtTtgm7R3OzZlnAVZtzL2qx8Vb2xD6VfWFYurCwseskKwA9CtJDhBI8ePcS
ovQ5+j3MAgrIdBaT7v/xqmqKwllTid0mOiJsgNtanDLbky43p16qCbjvEP4hXQt8
AOSEBe84FwVJ+FzG2HL7CfXEyg+6IndWr3cPOETKv3cHUYWYCn4kcXGRbq5kX3C9
FfjboP6LDZZEz2yFIo2D+5i8q7KhGBpJG3Qxk+I8NlcuRJMnHdp3aOwxeCUET7zF
wxBOUDQAJoRg+auzy9GBjtjHmMJkti5u8ZnkrNzEYHUegf5+QIWADqwwV6QI1ASH
4DU8X/Xt0p/LNHeroQC86MqO1cWWV+ZO8Bat/+NOs5Upr56IG/Ccse89p3yoqNb2
xjamWEMbof1Gn9AY1dPxFluow9/WCIuozGEohty30GhtPcQkgMimM4tKB3B5RER3
nu9YSpn501JSUo5zy4RTWBp3EUYHZAI5E7FGbbhPTWt55mwb9ctXKjllztbk8z/U
alFpiFeoVLfmazgsXN5j8bUzExiSTD3INCMbZxb5h3yDe6CXxYoJ1OkDWpyf5Bqm
MuPLFepKrCZ5pohAm64x0zGD6JQlO+Xfp207episNJMxaaUm3+asMlI+y2EjTtyq
kx8vJ1j8tfbio2ZWYmKCuBb1ook7v5nD497G88iB+rCIp+4uWBMEdkEH4apnrEsL
VdjKEsxdyCSSiPNdaq4lFl3qhDnYhO671rfxBtUJdPCUl8GzVtrlMZEDtpRn4ljs
ppMoz4oI+orVz3z4p3M5a/g24FNoI7lhyIakTVAxvQTJn4zZiHjoSrCBSQ6WIt8o
zG26wd9JdvOWIEqJWiHDXij9Ms5n/GcgtskhgQpAJfjZtm5EOuG9R8wJOjZl+s+6
cd9VrnvTFafxLM9q5C/mczpcnry9uT5HFwbo3DdUPaYn5MJ5Hg8bSu3ldNH6HjQt
OGjzKSMRo3iydlYfrAfwNy80HKtCzXGKUhq3tEW2iERD7d40HsCmL5xNPtf59SaL
YxHDQ5ojjoVM73PNYeFscjsIwGmQz+U6o4G3Lqp6zCsfb2kK2jlU0im0NRUXN8h/
Ve3QpmUnJtcUvttPVITNNeEssqjeH7zWSIyvrLR8Kq5Q5oQjuKlhoZUDL5VciqYk
LdO2GRemxrXYRA5YnC3H1r2bZL6TPYRNDrk1RU/pid94CqYQ7LuZfRf3/UzZMzrE
jvNf6o9XwihR42CfK2LFNVSHHX7blueiH1tepVmUDFfM9EbOBLKLo3TSfBgztjtK
PgSAfx8wUFfxMGfm6JpkoR14LFlHhxRUzdWnWuIofrPAHdD/AOwsFLBGrckC85nw
nD0dEuek2XOXamiwr9XuNEDBytxnmuLcIyeNo6N2OV+XCvj4r3N/9j/wCxpr8T5V
iDCjJt9wBXaQZ1qXI17s6RAZslAh6zNXjKEpQhxI8FxkDfaoo26vzWRruU5ZsHmq
cn01JX5GzZ3ZtBJgnNuYcKY800w0RuCoXGbqTMxhuogSySUoocA/Q18T+lDR2IcO
VCWZfrHOXAwUWnkByht74r/rnqmeZidYnj309ZwE2wgyzex6M/PcU2BP0+HRbyOe
xqPwjVJ0Z+I/OiWloGGppY8+kbOvKUfdb/dBMVvc9jM3stJsCVVxQgydeD3xQZUr
PzSGKh3QPu72CPOvpsZhJvLWKBIalKO51qLCnmeJV/5s6L45w9g1VN8fpBdpSjSD
yTEir3sGC/izpUyHKrwcDIN9+eeBdeDzHXij6pvYDIgZ/3dmRZaZMsdvFIZM0DKy
0xNwWyY4Xf0rl6awOdfH16SKPh8ozIIbQAtVJFuzEZ83rNxi1g9ShwV4V8dOBB2I
pg5szdJdk364JIVwUqaC0mVppi2b5nHGV9uHptvpGSBOS2TtdioMNsfMkpz3BHyE
9uTJZULkaxKNF9obVpOgSIudMgS2uprFXGZ3dLPQHgdpYf6rG/Ya4vVE8UpJhCi+
/N5Yj2YAoj7rClTBaq1lLA4AJRT+EFvKCwcG4MgeU53TaKKSvifGN3rgd4Hao0HE
Yu275qkdDVs1uaIqpUZeIolD4rT6dRYErdnttG9BPTpaRNTxHvevH9Zt3LjnxNqp
btgWwjoVzFBHB9yCO3qA0eqzC2+qkdPseobkQjhKCm39/9vZg/hwjeHeD3JqkPrF
9hz1HumPjeV52e0/Ls0TQnhCVcPCE+4NhKx88ClDTCrYY+b12CIj+iKXF66vMYMK
G3Su5DbZzqJ/xxANYo7yDmNyHgROL7X55Wgz04zxuvdysfyiv1PL7hlEZCDTuG1H
0i4TsdLhUuItq0aC2o/02ThLgV62i36aLjYLeSiGoUFy25OKA02w9MKG16atM4d6
1briP1YF1GmdoL8gMRRJxKS8tqFOan0ia9Z9NX4rhmr8Lyk6csaCaQlOdsCiH6G8
4T8jYmwsPqfEsRLsxl6VChixX7w74MC9AtdRh0mxFfHYKW0NDPnW2df209bIsL50
vo3lnCD59tkYHupFFqFq/J8Po0PziVRtlGUlTD0MMAL0G6F2x74Zo8r755AtPhcK
pmYawVac90RLakSrRiUIwYnMVnBlKGnO2ATAh4rrvvdV/TiBof01XqTww20Bl87f
yIynTDqRbFmD36kONhe1c7PIPWOmPrtfCxrvddIx738TPphP9z4ZHN08swS7FsLE
7dNYmK83KP1E1ki5/tBPCkCklnxQFGEv3qooiaEgvzygOsDU2dBIgHiGb2wBz5Tl
ivLMFC4/sSMBA+8JNTO60csUP1kxyAb//bUhBRtnroli+WNZL5xODXnqtOud0fMX
FhSOWZaJelB4ZztRQ8tMfCtQz0uzzexaU+/HYggHAnGaHlD7ZvskGgOcP/vlEfsD
n3mMNbb4gdz3EPnsRFX7qr8G3vf+2XB+hF26cjPInMovhC4Xt5yr9n7vHL9Shw/c
FkWS36EblxgZS3mwJ23g+aDDFYFPXo65F9rKmdxMeSL7j7XgExsXqa13udy3Mozb
DoYRXhg2c/y4PnEFMax+FgX3YInqHirA0rN2efzaH2cnJ3cmAflWhmqTpyybMrAB
XqmmnqKu10AN0eRTN8VB4uDX8RmZU92BMfuk7Llga1FLmN2KhlaWg81dxP8JaSma
okOqs40EEhv2S86G4Ncc4j0LlwyLVqUMb8VtkrfwAvApKas6aeZBvNuKP+kxNHq4
hfxfgveQXKUwhmgSzRi5tkeEnnWDzbxa5D+Rz/12Gpeqdb1BuLogw4nuKPUS8onK
YO19/6S2zMO1dC9GpyoxzlxkQVHfb1Um0WhmJ8r22Q6qmtlxLplGW206a6qzjCTL
d7ZoyKhu9qwXUkkV7tJmV3jDLW2YLhnU4V2HX4Z0IOkiAeqyMb/89yw++zpD4gx/
aZvGPcO20y5wv5xdT+2pgbW9xonjjuZW+V5gRN/JBPoY/uU8uckn6B6rFByqrRNW
HAgK8kOmAFSwL21was3j+LHE0aP1+o5KjPK1Amt6qxMZ5mDmCmfeUrfxKsN7auH3
y04mgb0iOjJG4jTyitOubT1nzClXhDt55DyXtELOI70UrD7Uq1VYsjnwCyxE7hQg
M6TufHvpLoGwDwUEI9L3wsuucMAs+r1WTgh0vjmiUFn6cBtMpJZ33k8xUis8xRAY
zpEPQd9YuJ/m1A0dSZ4V3jjh8Ooa2pY7FK+wqx5bFVaSl6pmC/NkbaT3TdQvJ/pl
l6W7F27dx67kvvoSdkBtNa43Wf7uAJjpU+KgOhrcN0CAQ7YXN7/lUyZUwoWna+2Y
sszciBsRkRvWz0IMCPrU+XdxOieKpwPwwX1sxpmybAq7NB3pI+rDQiXAnXyNFZa9
Z+KQpT5TPWaRcv8vp2rUifshV+ykpIjgPPXOazzyI5EfZmJm5XjIwwoZtMAaROok
Mpx5aNmQ4Zhf3j20LKne/+t0dXjvHBNSYyBT3lhk9yLa/Ch28KTnq3u7Ccgc2NHv
7lZkU/owiyEnRvMMDR3TcmYfHg1csup/v8Sz9vjSpmEVkx6Y7sINW9LriPa8j0Yu
5sMcUI/w0MltZro5PRytmI3LXoN9JXUaEV31jvFKRrdg7vLrhb/NXXfRiNXFgdz9
Gb1YJLdlGOibmZRfZn7KYPGKeT6O60RuRjzAjTmmWX4z5jfbiIhzvJBhruS/0JmZ
oJZqvcsiZCAPawEfh5TbfsZ3LJeswSnh4CuXNwyGufur9bzkLnJchHAHLRzQlDRU
EQ5MX4qyTUO2k3MWTh/+mSZDkyAuS3XUWJI5za1ii3mAGGTMVq+1W0tbWPuQXKGD
OzDQQuYnia7aUDsXGWT7nkyJmT303eKJZWeRfEMnkxmsfWfp4Nxg8q6fDc/RDaZ0
pz0huOqayY64a20JxeHYXc4jAytrJE8CxL+kNll1Qb5LEvirEJXU2zkMAfQw0FIx
Z+X6q8lLLSe5iW02n1yCtbzoxckAXQrmoVIa94QS1qHY8qd7WT0qGXIQdl97dHtz
zNAUr08RZmdSRLf8J1YhuAwDWeWf0sZAAuuoovhZBkOZ427L/hlTP5aJweEQ0nek
fD1DXO6p2Aj+9W/HGz9fLvquJYiM2Q8iKlpfNSUXxi7stkMFEZ0MMkJ/pqd77ihC
Yy78JlgQjmNuq+mUzTA7YHktoiuwAo9wwvkiBXRjqVuLdD/eGZbxhNqmTysMfQB/
Q/dVrUyDb1d8KJqAk7opEcpeGwAWwuUTT6u4GKQjRtrdRSIlyi4Io2vJlWhSr2fw
J6Bk+zgQwQYniZ/QgSos/LCnEQo6x90hKmAzPbyB3iEhC8hCnfXwHXIkhMV/tPoa
J37sdYCkK5W6yEM0nn1MGRbtQ9bCNhCJnA22Di9A14wkW0tdOWacbHixDwm/1UOY
YVKhjpEvjJAFQTDQW7+beZiI4seakziepw+d2EcZ+bz8syVdTsoICRT/ZNQCV2Q4
cXR4IqyMOhGioISpoNuwtPcNIKf/Vu4SeisB9tsOMQDHNn+JitJ5HlCHHGfsVjFV
/YFwaU6fa8/6WnchR4EFuPhCXMOByAvlbWqnCGFt9m1AAHMXE/orQE1E7p65bGR/
scW5QE4JRJ2k6R/F+c2PBd+qNjZk2cIQ5xMgzP/ejB4xrBJBgL3oaV4MBYnYVTtz
mPr3JKrm7ObizWoJeA9SGzf5PGGNyEl+JxJUiX77Ned4C4kvyUgFYKSdvx7NYrT+
3joRJwOToWviIhcYr39cE7LlQEN275xijKiDZUuugP5HBLHQg/nQcSaAFagWG0dd
IrkTmS3/jjrXmNYBrw085VxZ43YY6aBDXi1KyrXKZ3cDFVK3qO/neRUJAX+Q5kpx
aU1lPDOLDbbgJnO6+RjDKgzrKjbEc5sEmDuVE7T477eeVAJ3t88XYsIf/Tkn4ttA
joRF19CtSoKOzurE9xVE6jpwu0nF12BaHZX26Wfv8s0YauvxW35BpkN2QXhrtx/o
38ZkhbhEhBUSmDe3xEnDxrUqOIb/WYIuRxI9QXmfr8wwVXE+xI5wkvM8HmBuM0TS
gxP9L/mMgZDEGxQ6XVXj0Ma0CQd5oemkyzWU4BHGK0VhwAxWIj6tNHvECrMAY6Ts
nebWyTLM7HIfp9kRgdN3vntJWr3rHRzmj/2NphPyBKy6rGbWaeolh7aGzQQr2BZk
GJn82JZHyTZUN5POeMIagp+5v7Ad3FsuDAk03d2TkgOqZxwAjlmi3haEcQWqZXqf
Ly/8oFaL/1p2FWyYpC2adJgEqXpYr44+cIIdvPbWeTJeVcRGneBek46MbTgH3RTZ
WDltO8DBYekVQdC50WBaQQ5ogKFwATz+g1zXUyW+NbeptTlj5CyHWdTdW8Q43vo6
zGe0Gj3raQ6/ME7i9SN9lw6RrCR/hbGGfjPIrZofkfQIl9ZMuVKObi5yNUNG1xAJ
FSIQsufwJ9O/lcv8Pdtd43XlcqdomAlDJMPrYx3e9d6EvXebWsW8lpBl/PJq5A7r
SQt20RunO2VYlnOLO8tokMK24OmXdsqQWeRgDkKTg0GtzqaDiA7RlfT0/ZBXvf/u
sMoF8nYNVxsLB4yMp1MLnzd/+tXLNu+dJI7CFweLO4dzCrwKb6pK8UFd9STc6UVs
hUtLEeJh49IeqY0ihE5q92WX9dfNvd9dquaFVNDDtVsNvav00STGmghgCeyshYYS
G24IWiqXF91su5RdyDDnY7GTa5kyvXTFbQ6kwtLDmaJn2/U05tUOKGaqXBqa5BeW
EuT48o9wX+T3oWB+Xr5T7AMVWCf/YZflupzuBy74af22XSKHGkRiqGZNjmHINE/i
URpP5T077sOvGjb3xNHYwtbAlkKEG+xgNnf8EhdYgL010woRMIpaFT8xmSCHIRot
tBSc0GioAO2s7jDE0zCNBmMwnkx1JGonPr2a+73vVwv1Zn7JOJ7cv1zugp8WpKis
r1TCVIuRzxV3/VuFwRsyBGkVkk3NkbDkY650J53QMstsxYMBJnFOI/gp1zgQNa1j
W0tGFXPAw0sueZ3m0U2wVcwUbuXtwaosDT67F9ZuVRGW570uu1Z4y6+NGjuBVO7B
xmalpGmugBeLTy6lWUI4b7nFd9vm6nQ7MRuBdUVmIcCQRfpXCbT4B0PhsLQBcE/N
jdrdmPNXr5zHPF0zRyp3OqdWkow59YL1Cqsyq5pmZwFJyEojcgyR7koqVlyHgyTW
fCc3qfxy7ab0IYG9Tovi//PZIXhojnWbOYN3iWmNvO00ds9ikyZFea2ho9ejvkut
UBaUnZqyuTB4fB5mJ9EP7wc24+0RijDTwIIxoPgIH/PW2x0ralG4fIlAYvt/ZLAX
9sgP0R8ZOeB2QGBUFIVoSNP+31Yd0362FSIkH+xEl9gY9L1unVmHtxdlF5xQH67J
X27tEazgBUd2j7kU4bkSCasr0QrYCyDoBZze5PLoh4VyK7pRIOeTCG8XdsXKfHZq
6jUMrsTDJ49NgQX64RleOF9iKdm4I3JeHv1jhSJ8qKdl1UpwScZTQXTxuYaO61z2
fu3+Qh96/tz6RRmaridpebruFWOsBeZjTcJIzjF/tPytWfzajwhDq1vklQP8rQjk
jM0LC6wH1Z5de6W8sb3v9SAHnAcRH3dmpZzIfk9ap3cZpVCPyTWEFbx/3ZiF4OVU
0xyfaqBDga4yff3UeyxLALLKOwlDis1wLgnuoK/E5rRutcuyuFVS696CyPwAB6XD
kzWD5JPrcZcUqhsKJd/AYLjozMJo6NPhOnjCuoikdH8/dGHwx6AF0fsask/rhM+V
omXj+oTM+KI540q6MGaZtuhvoPPBoz6JrmIq/qxcHgGe4PkDMsEprRMKi7IdEnU2
6mZEVlOiSK+nOkybWVLzj6fejhKFU1tS560Inpg5bQgpWx+lyUJbHzopKIcht1X5
+ff/zz0jJ21NE24CjRbvxKO5hnlH/T94GF4xkCSc3Ui/QI52nLi5kVjKgk93Q7/q
coVHIT5YCGZP9Ht559c0Cj5oF6q+HCOQoYcbpDoDljPi3StjP52HweKDnDf4QvB3
gZac9pCxJftuRlsyfhA/If8Xl1IDoDZr83nJFcHda9dT/klvMtU1bU4BNg9bOX8X
nUeST+jtVtFYmPhTqKv7Ox71E5oo3dUtXQm1LGcdWCMEVBogen2K+H79ztyeCpz0
v47BWBJ82Y3P7qo8adTqt1mEOZjt7srpojju4NSSTdhjbva1JguEcyaefv6QPIPD
82JLP97yjz4JMbpBkUjLeXj7CHgPzp/Y+xvQmBrp8va/2CaASOMfLKTUT/40YRUJ
mVCTyIAZjJzlnp/gVLGDZa0rX45jcijjqe5qVUNysbLT9JwZ0UnRUYyWqwFA2TWN
/tdQIElp8WQFn7bnPsebLpcuI70z15ES4mf++weje9UtJVRmAooS9FtHdxGVVxPA
jsn9PyM1Gq1NHdK9dBbjGb5Gk9/2C4jWQrBcz9VjnHNLYZfRCuFM3cg7hOHaJIpW
j8jvaHSSf/4FIKwDgqBhturLk7MH4YTJADnZhEJKjla7dEpSenhQaZRqXqwrOlhg
7IyBuD3KWsDngollgHylAGclJ0hEry1sWTY9Eo1GH5EaWz09qClR++SmNR0THNFb
D0t7TqU4E43AJtH1mXa8BprfVL2WcV+/n2RTXNe1K0xiJ3jn6+idAOOpX8T4k3XM
mdgcSAt7VyhvE1sScfOfzvyWKNSW26jklZnBVdumoQFT4lHkhWq3JrGfA0T36X9U
TEmQ41zKf/JRcUUFOPG/MwLfgQ9wgpgzAi9l/FXWBvfna6KgHpiJw3iWCuw6NO23
8RdnlOze2R3pnOKF8uTAhiqBIh2EtuXOd39L+H06gaHmRiDC6qKJZrPmDxWzposv
LjeMQSLKo9l6Amr3oDYflwe6uQmXv4wtMz6sx9Wt7d77zlOV2xvSQWYVh9AYX6hx
fIEsjQ9Z7STnE1EpFG+Mb8O5BiZkqs/p6W9Ot+yqy8BarSB8X6Bkv/0ynK72C3/0
sa1BgLPVMrR40UFvSQL6MucDjxvUO59VQs+Lk/eQDcAOe1spSVs3kfC9E5WMRuL7
X3xCgcm656Xv81oK7hPXJC0EQrpT64DkBwjWFjD7JtGbpFuoe17XG2Uu5MZ3mIbF
VHQQO49+cugt1W/5OwtKV9zHcOe7wXigi9qXlV2I7nzFzGswBMDCjPDEOoxmUBPn
k9zzIUExh3XtLaE+VKiCycJp94Mcuphct2enqT7/LOLKfoIhcBJZjti9zd3Sw/wE
epwBbN0yjVMVmw5rbdOY2NafL4csJRiBpMR2MCVVB5IjYka8/bzSfpSF113+Ftkd
t4Lp+OmRrciqtJcHKxikvXJeskX5lbekznI2azCnMn1nswoxDs4pl/deadSKKG8X
7tB1SkZXT5LRSLhieyw7eRucTmDhuajJGRYTMfBhhIfRqzFZI1L93mkxGtGcTxUa
SjoAw3vCrAKAuKEl38/6q+80Kt29lN2apUrqK4Q5mHzp69I4Cd4DCeevm4IP4n0j
iQrKcFDBs9vIpGcs+Av1USrUVRVuuTplPpyFpjxYQsLwFlIWBBUU/reuU+7oyFN1
MAjcHgV1zXsh325ZC4BdvXdVG60JE+/ZF9HAPJj0WQjPUCMBvIipnNiQOwa6xKGX
X+uh4G5MDWqpZlvao8J5UtC9aBQ8XgcpJRtYbihJegoKUTa9JIv7XC0Bxmi6FG0J
8j5ZyN4f6BARmMn9W4wm8yFa7o5nX/HauH9SCgPSBKH8gdr0zRu0BF+nZX7jfGyW
yjHQ2sxIrLlvQD0g1LI0MH9l2e5RyLOswfwEEHtU7df1Ai0k4rtdfLSHypsxL1rG
TdqGXgMxYoWD6Lq2m0w1wbKkDlccnf6t6V4GeDYoCCEzYWhdAoYfuYcHL/TwwD90
OkC8dVx1a5rfxeWpBokvDSjhisouyLfRxrwzRvsjE5oGDesuNFFZNbVem77gQJLs
604lQ3qg3FwUD6lnPtHWkIU+4jEp79SnQeLZrlYkQY2BP+Fmkg+XH5cgAKbPNvwV
qpTzMRrlIwS2pjkX1dZ4HrEISt9A+iS7/DPyEJMT8j9weRRX3Y5d7eZ6WspgQSb9
eLX/Yr+XlUrvaDKpnVDyAID/8ewD4/pkEHVLVMc93YHABqGXLvvw/R+AatO3fKrs
DrjP3OPrJspjLvmZwMRx4jQ2xSyYFuop75fkl1v6+1nwV0Un4qZz3ZyttkvtPk4q
r6/oVd8yG8vbGA+TuuBavQzvhvHNo4epLppiTZYrqw39XnMuh9pd85E4Ttcf669K
lNWTUOEG9JBM9fJZXXTvZnwhlhMsOvcdYZD69Lfc+mLTxeiEp99rnC0nxCTCBY8U
HsE8gv9uUAEPSMjpn7EGri2JhATI6vixuz+n9T264atSk4g/OmrhotlAAVNXg5h3
1jboU1cG4FCBmTX+ZDllni/KpkFDBdnO349BTYtj+rrzdjXWVy/ewump03UJz/WH
YgPUTFCbKjLJNXfxPrjaFOSJDPjJ5glNevvnIgnJyWiSmY1tTK2fOEuBVKsn7+V0
Ce097LLybjf+FO+OAn+kHWd51qrICDq1WU8pc9huof42IAfH3x6f3PrsjWGVQR64
pUtD6wiei5wZ956w9Sm8EeG46L5RniYequ9l0Jqj/btUH1/Q0GGiIEg/1AB/qXsq
IH2Gw0bY23PjvpCQ0aiSCV/sMczPRQ3jReeayGZCwWZgMYC7538hF0xzA/QIWrxv
QBFO5jursRLzII9Lnv9X2YoolIK+vCZx/75TvkRgWQX/jRXl4GvvefKQS59o6xzO
pWelPmBAtaRQfGrbPpjeFtrTwCYR1RCMG98YhxjyfL2RuSXU809MdXZ465Tofn3l
W6MN8RMytfZipi2dvGh5uIFjdsDi6hoEIO4udselvouM5lcgCvnURkvnnIHb7P9S
Wb/PykK5n3JZ0eEZVBlhBUSjwtSE48yOymxfl2KtZEGQSkUBb0/JGvgAFwSFcTxI
aviL63upHmkri8BAfk+mpuVlWEA23k8bieAPWNmzBt11AgIF0tRMecd8F8YTS8yL
qd4KyPCiWjI+deRLp7kN+s9pqVmTwipUOL8clCttRZUzIPfA8KhtfH79xgyJc3/2
n2ajmoF51L/D+lS9qjaOU2mEpPn1ndRglk77mbamT0qXMgV9zeW6k8i2h361G4Y7
3Tm0aFQV/fqyOH84bAtli0AGjwSHoT5enkWHoGaNsjcI5KubF6/PdyAWzxTYJ2A7
CMF9I86i2nU17btmBd1oDcSvWw8+QK6p4/ihgxym4Tu2ehwc3E1ZFmAd/RRzgnqO
Q3AmTcUgZElAdLkFLrlq7ho1ZL/X0Z6bBqN0bJO0XoDBTh/JYnWfH/H6rpbxOfpe
QnSZNJU9N3MsG0pn3U2YoZXu7aIY7de3+4iND81hcyINhvrRD0FQHqNN/miBd0uQ
CIqy09IFqSzVcprOkD1zTjNc00vMk1MXHpVBTdpgqB2YJgUFBu1eSpgJWlbFCdTA
4W2+LKuzOIAPY9KjDLA+bTbqxbfu8dBWJbPkdijujNi7di0s8MqFltZD+ZYaAGg/
vMGqtux2Bz/cyx4VxAqUS4My3cURcxFNlN8gBNyfO64pNRsNWxRffiKVDox/HwWO
POVDhh2qjNjsKDwP5zAIfQ4nKi2pbtfS+N+2DfJNcx/uUzlNpg/djxJv8PF8CeDn
HuxFW+SidqE26VYSvwq6yaMy5P3yIVZ+dA9hhhyPWQDwV1S9KTPI2qBCvl7ayS4q
Fsaee7PCK0a6wsT2FvyWIKmWVUEd5XkbPJlcmjzCkuk/hzvm4sTfdNP8Dq4orSfm
HL3ab+/uCzKuTXm8QuGkEvHmh9vg9MhihrE1UNlOHmpsk1RWJsy6g3hAzQKyX0YV
RqchwsXzlJ0yX3dv1JHeqNfOHfE4nGeTwyUQEXFl6i5T9ROtuJmXs8TlD2FRjIQ+
HXNLeeZHFiElKetFYkdspPLivvgXUYV7YVakl3QjSSJWa7h4CXiLjm6oAAHYc39+
F4Ux0m5ItxjBUAaZPnc40n+fLVM1VzDKWjquXURHfSwNs6GaQFSosTi7ZGZbZYy6
BeAZaDMsLziu1ufQ9v/8g0LHwbl83nJMJo16Da4xMl1U/TOnKJFmlZY7e1oEOtRu
epBBgK5J16QBajl+8nEaJ0DyQUsjFrR1WCS1ibAtEZqhUap/3EFzgQ1QfJvftcLq
OifDKNAuCBgvglIYceTIzhMQMNqWUK/B5n+n6NoAFlhKcaml2tGuxI3YiIcC33yv
68wKZz70dRDD60/lojzjw5sGfW4t6WqikSfeLms5Oae5iquU1Mv4o+vf9cpGRP2/
LQ+j+5dLeoCJQFkJ/UI9Pu+lEn2NzF8Q3AZ4E2+cOnL7P7ogkNbCsypLla8CW2VK
6NxtNtidVGrJwknipV0TwNxzWug7OMXOfpOYsL/xXNh80Lcux5+1joxLwfj8Gqrw
DYY2nra8w86QMCvCHMk86aiKCptYmikVwd2ID9JG3C+cRAHaZKXVQO5esXcLqtDf
jD2po/jliXfzG23SXa8eRbNh4Fr5/W9mfd6R791BPbrQNAGbujqiK2Z/LliTLCUe
Xg0uBlcGgCI/SotHrb8QFP/UgV+aBTVrjTS/VUO8zJtxWS976J0CDWoc1FA2NPAk
kJdkyULdyP5p2Fsd+TES+kSuhZ850LLJ58r8baG6edUQVGirpAFyYHpXeAYorE8C
xpQw/xTyll1QKEykyat5Ncg6Sj3HSRsWZClajgzThITGjAekZYHIY8rbxNSYDxZS
qPeoT2l3PPgjD8mANqvfwXgTEYNEiHnWfMVs3tfr2t+7Cm8Wib2WDpWyTRj7nQIM
s7iNoNtH0Ww5VAO91bjW+evn3wbWlOkktd9upa/lZhInoCgPbFb+vn8V6kkIGpcP
5GkmUok0zxU6lRZRZ6RZAWKMRKDwBNCWBhn2KD3xy9VAgrmmF622CFIIXx6HsiTR
Vp1scls7HbUPREo4WYCMJmfHqWaGzlgW2P6fSGNy1TtxR46PgxRF99sc0L58oFH8
4cBgK4gn+CfQqYczJmN1TBt5eTbcDGkrfK4ZXOne9J3zbjt06pz40Dkza7IEtNpc
diRmPDnDQqt8F9qci5pF2/rjfXb3X+dV3SVgAN3xxFj5/lL7buN9ITEEKWfD6mVg
iMCAiebGa6ZNduy/TYZ5uA1D+l/s8eEbyYvj2Q2d0Za01fY6Oh9zp3f2B+de2aan
LqSI4793DrhCL+0fAvmUoMsM1+QGtA6wEfTmggX0//SQbo+pnwuXyrRyATI7nKfe
7rKYTeX2J3Mn0bUIzRsMAV3mR94QGY8+2mqWV7aVc8JmfHoKHaeKjC/szuJJRPCI
0D302hQxekTB5X87gYjQCrEPy2K/Ciz0O6waJGeKKkxOkWkIGVDwzy79qRhyt2ka
Dd774yvI0GFUeLqmmIX5dRvqycI+NOkPB/Qc+ao3dhh00pQu/tUVvzCJM5ROCuJS
EJENQcj0aOol55SL2lfcQCCVeaAVZKPVaqNpNF1TvWWYD9znWVPfgi/DXb8QYe8o
73IF9iCeKI1me0R4pQ5d1qQy5wwHDLEk+J+pxzPq+rVkCwDsQ6IjVANwqJJQtanM
Gw0d3wES3z+jqnoXl6LQiuYfi3BYSq85lEZJC2nFLctAr/BwlzNxVWSJcQccDFkj
FHm5Xc2KyXrotPDKvXCPWefaAAeVJzzn4Ywhm3gnh6TxaNylap6f2jofZaCt5drZ
8Q5rLa9ZOKvJSlnqZzXO5+xj4CkhSNTsFC8zpPOm64P9aUVhzs5k/oXIjC+NoJ/5
Swl2q7jj0cr5skeqxwMaK7nqD8qxSuUDzkD4QX0SGAkrbQqWzWElfGoVFlquaXoo
o6okSBNrQdOt3WIk5yOhGyOsgnHZ3apsNegUQuY6oVGHTmgpg+NcHy/RUuDAphOL
1cX0ugk+Y55StS7imlI05h/JkghLbzpX34w3RWwaQhxsFkuiOZXpENyKIqImdKvQ
5KN54Z75kEGh9gmLiGqMdN9SLUXneI9utNqtSvGErGfz0FSth1rwQXRGa5Bu1O6+
3DWTciiio2VNpSNxlHL+fe4DF8A9EXecF4/kSIgHde/J/P464xVWc0yhVVimofnl
swx8wV6IEu2dmElx3tEShTvdVssvi0BI0rRkr40tpcew6h1oOtBTU2UUJ880T9jx
sZj2ypPc8bcXy/a07wayyaNUpYxTTVTcNOp+0RSq04N1ivlSauV6B0/eZW18ZLcz
zG2SSudfEGRZ5pZv3feGdnN6mWQMB7m3BCi4Nm8xMri0013KBkInkaGTsGkgkZ4T
i0EhXODMCwT7VE1iu3exdn4hFayfujYHt5VsE4HJ4VRgyU3U55PbjJGFQokBOgEW
j0ha8IkCf6JEOiSM774BiaQHuG6tsQKhZLwTuBvSGjMzOaukEPLDxtuI9Zoosm2L
fOxc3KDGEgt/tcg4X2zZQB34Fv57WUvkC3aRKQeDS95QG3wUWvEKhRNf57qeqaTr
MdUInsDZ/V7q/7NGoHfVREXYfX6jKo8muCxoMFPYGzEhSXfKxUl84yFa8qLwOmim
uAdvfAnI99DtIZitN/r2DOVDPuZfWHk2IElPk1RUGWFxF20dfmlEXNaVXV28WbSt
c5JxmUFxLSxS8xrxpHd6/4tpY9R7lynXLN/8Nx5X4wT+yiknBSsq1slQo1C04ZKN
NdbiUCjLCUpIwz0BD6trn5OTTWAuF8p/gmiTVJX4++K7os3dTg6YDbrH/pdtVtWr
39m9cgxniKSMwAvrVG/IlTFg0aDoliVMjgfUomOGL6kilbP9j6UR3Whb4XtYnEst
ESYpdZ5WNbGypfAyHXtBAPWVXb+mLyrfQmZEOzet1R/0KJur3IAlJw1RJN6Fqtd+
dMe1Ao1fSuL24kWFVdd4L3i4Nss3fotm9zuRMqImVgBoagdjB3zUL9HmaaUMi1SD
YCuM4DXi7n+eB+nHubqsu/I9w5sEviroG1lybNG19vBp7kfmEEDMKRM95N7SW6/A
sFYDZ7nLfl6+8TqXIygw+L1AMEOBhpzaO6CD3/v2RKl++ib6IrM5AACrKkyHRPcz
y1DyLaFDkNDDcxzju8ltLfUif94Gr5rLsXqMJBa2UpZeTbNfelWU4FziNjOEHTXK
8B7sSDfgQ3BObxYX3xu1jXAyN3+AUTNBC4ikCbKukU9EKJ2TTOLHHl9AyGI86wnm
uuDsSgRSFlyQMCqXmX2HFCS1j0/EgQ0LuEUKZCc97NWeKjHmr2NQY8NQR/cWSrNu
Cwbnb79YN64A7CYn6gIevV6AOfhLI5fQ6W9WtmPPL2WbhDQl9yH+A+/5swgmlG3J
FMKdz2eSp0WCBVvc5or28yNcKg6xbndkuF6wciE/npz89jXji9UbPG/1C8skIl56
QhTleP4rnqLOGH3KPl9O25mVulQeoY4FCWhpbEGK4REdASNPv2FKx2U5W1oZSieM
hcSq6ydPhJJTKQPMQfiXMepPQi5wewMgMHOjfvqouzWSbzVqeouAAPfBn5Dgxbbg
KzxF4F52bDbKYOMZHx5pj6r4ncuYELQphVgxLLc3YFoLs6icRAdoawnGC+n+IsQK
DpypaPkOXLuHnfDYrOBsOYkuP51Hnis5aXvA/sjf5Hu5eDocZbSYNgorJuuAIMDz
x5hvqvBJot3Z/tqkYsGgYpvlUhsCn2RNZIuLfvIOljD92aeYOVxYrTmujO3i/C8V
vPjbTEoEDYeAhZx8uMKYIOumx5BBMzWuKuQRPZCs36Oix3k9io+QDMsqM/J3LN3q
pWK9uiUcHQYyeeDJcRRIzezY26D/J3w3cVo86ARI98T+kwjssSEuMsPqllh4P7si
jJeZemhKe90+SQ4LxbEupRWIq8sjDs4e9X/2cYtluTi+gOqNUBKp+7WdjnMyl4dh
79k++1tRO0uxz8eNSNRUES9pmB9pOZsj/H2isedr3oQz/d+/ovcS9zLEZ2qdTSsE
CwTQcwhNDgSfougPqOUxVqj+KdnWIYWRMZHpVtr1b9YOs5YUlI+yjzo8D48D1cfu
qFH/pEUbh8HjREwkD3HdJa8BfebfRuhmETgCeXE8JIbPefZe6wSYrGf5CObjMcOg
ambZlO9iUQaIwnIdvgg9TwmUAcPWcOUo16KYZJBXf5A6SKDI+aDUv5PxlWpkB9Z8
vuBWPyQQcAiCtWzkb68qxweMqi9HwVyBVBM30j4tGAKZOpCwpWcAnJXB70AMNpzR
2WiugXoNgWg0CY1zFY25kNaesVwWI4gEfu06xp9EodgxAT5wDjGx3Bo3/hHXhjlj
F0LVId0dh2Knv6YDmN2zmp3mlbjam9TGsIL9nhvMXD/vtQWJXkvo7KdHHcyqTcFR
bKHVMaJF7zgrGC2eTdr0PTazIUwuhqOXXyR41NPQUBtFn6io50E0dSn8YPOYSZ3B
OWz0xyFUVCI4oeQc5IZ3zC6WHdzlQSMGKRjtDoxDNmNyYz0AeM6t/VZYjeREcdw+
DK1sgBJssdNypeWPes/rjmFaeOIsqCBvtNglr78wlyJdpRpjqPdfoszxgVh2pyeJ
RIvMSuHLRqtYPSv1dh5HvxCpUDHzkDMrcyxPEpzXp+/6TOsVJEtL+5V/E7aBEaae
yMiVXr9va/6QYpjDeRoWyAeaubZiQNsr0mcWXi0X4e3D/Va1KmFD6AeXW2qLhPZI
sW0WvgYoCWqFij0zrRP7Xy18gFAAop1p0xswa9dzus3dcAbTeGiaWcaHK54lp/9z
BEnrljynPQdmPEOnlxOFxG35cfckastJaxRn4HKmBPV98HBo7c8rW5G7bX20AFar
xCh22o1Ufe+Mp8loc0xJUWTtl5gOJ+X8qkERLzqzKdFMYNEfABeUjgDmvCkkPzjS
+ovvuLWUPWUmIPkCoR1/c+EkeKwPcjGYGY6Fg6rRaYC2xQrAPvRXu/tJ6dTvZ3uo
KKfGZvBux1soAUspoz9qwmJOnO5w8Xj9jiqogdHcYlSnx0V+NP6PVq+oUoAkD+e6
McBvfy/LQrof7V3IZFAT7SOtlNeJ+yi2Jv//BTRVOY8Ajzoy4TJaE6/EQRzAJRLr
Aha0Cnc3/v5Getr8UwOIyOGNIHNpNyy0bmqra7tdUwZzLmAP4k/wtRfGnKfsCuL+
xDBGnSfNq4P1Qbeh+KA0kuR36M2pSVQUrtj66lQNHTQhq4Im9H7DOHyQzhVzH3qB
E7V54CLhKVAH2cNSB8EfzgsZUA73bE3R/vfOZVyCxgYxYiUHrPRk7S+G68AtOFyx
0YABybF647ZxoEFEV+x+tocD9NfSdOcTUnU2HU2F4rVE0nQo5sIaddmau5kTNeDz
fzjIvnJcOUwvFk8sWkTlEYjbNc48gmVzHp7H2v6dxMnP0mT7cCCbX9hU+Egx7Eu9
fgdTDImQfxSH72nIHmX7e2vHLwCiVrZ3HW+OkP5tET68QjOun6DETy+jrM8rgvMd
O9umD7+tYHBnOW6IG1vAFt+uxs9YSUrT7BDCZDq5K23PLEXWqK6mZOks0cPNYEQo
QE9l5XKIVV3NHUeQbv0jaYI2rNIZVBLLLTbmW0fYV7m940yjuR4h2oTB5J5FFhPq
5RZSDF3GNwPgu9r+bdlchvs/zYyhculb/KpKd+YBYz9+RIjOvFvzd1YrtF+Ts2Wa
nkFCNHReuMDWT235nsNd9+hkQqOJ2My+aXGfZ5iSENiSjVYG7MB1ivxteP5YKlz1
BSREBc7arSZBofmPRvYblVzr2xcUDqjiC0DrmiiS/N4XOFmvnsHLNF+Z/4oEUim2
W+Bham10Rt0vsOQeAnwRpuhBWw1ypsocqjjUg5vZCW9tafhkZrsHLxdRfJGxQbQj
YjxyPSV3NOHk3yoDf/oInXPRnXPofQlOK7fFwo3XEPAIsdyZOtIUOTAlwV6E/2PS
AwmdnWaZmXIGO2V55+7Xb1Lnsab3Kf1pzV8lN79WA2MhEhjelKKiJgU58d1qlIDK
/IvMx/Yn9kfhnT93sgcpHAxz/Iw8vDwdOrWKtqYNkAZdowMwOptNGY2RQjPoKGTq
YcyZPmrXslSnADr7jgAnapFVPUNSrHrlD6jKl1stE+IcIsziRjTqizMTjJrOHPFt
d1NhhQMxChaSyoHrDDY+gkaoNGeCtYkpaXX7F22O5kotd7xi7RPyAcdnQ3scgyyW
3mg8GKJXpcL0BiAOl+PsHZh+4vreTR9WT1rzNADqRVNT8e7xqu+yWiFdGIKrr80j
EU7yOdJbsF199Y75V/zADs6adM+tDqiz4AS+NMlfNSDyCBHMBWStBx5GhRxXPBpG
Y4Zl2ND6r1GCTaJn4PeT0FwGRU0VVgDjqoAP2UZrIU23hHUgaOqNTMWIwuoNeXHM
BK6byhzwsml5HZPaj/WwbNIj9IQ/BKhCKBWuGi8v4V9Y55mrWpaQ6ArggszZl8Ck
kdYkRwVKFu1+t2et7DJhjSY5bqI0cjpEkkRw4yHpHe4dD7OsJdVJPpqnBfYc2SeK
peZZDrNs/Lm7pQzZKLZ2ozh2EC8WhlP0S2GFlZIgSisY0ZetzDVw7SABDR0RCvTl
BmNFOsZHN3N7J5TXR2tLaoFCVcuP+KS1RpdjPtK9vKvDQypOaNiy+YLuIGN2Sil0
5+N9luKjRnBUEUdIfbLIoczdmja6kv4mqPv6q6HS79qplP+1wCAW+2BBE8aLetPe
fxNmv10+mjeAce7Ur/YpM/tGaplMPMwpKTBtDhjH+LldiX2KLDc20LHgD3r7xynW
SkqLoLlh6LKRd6ar4t+QdZZMs5ze2RPsUcV+P6cwDiVGG99d/jRSOBMhO96Ur7yS
BY0heORPxjYQvCp2FR3M+HtFxkjTDtsQ5SMBiqMUaHUK98MkZKbirWOjK/mtsv7G
9I3N1iuUOdWJKhaQW5trB7UJ1cHm/ZlstL4nFZMTQvmadHzlfaeoTP/isHFHVKNc
WGviKGtEUzKWePuqy/QZqrdN7DJvujNJYEiP4s7FoOpOhKlGFws14bGjra237AZV
IWqPfUl16S5OIll8dICi7cYGaWUku3H6BoLa3Mebpk74e7h/kixEokutnZarIO/1
mIzGv2saG7tGnf+DrZYP+Z1d96UovhD2CWZaHF8uOHeGELMGLJaOr1MaQEXpqQmc
JUCu08wk/al/7UFjF0wA3jrP6oD1d5KWYJb51s3Eil7aXKCLx8Ik+cQusON/by62
dagoMpGzYiIIT8inksoUMawGw11qJS0lbqWC5sTHYOF0dEFWFwuGOkU7WAzJILJJ
beuUrD89XJKe9db2tSuKjWnb09iHH6sDI1JpcGSSyYImXBLyZvExzY2Ye5Th3iF6
PL5Y1KYNOz/OhNnpn2XW/vpcKocZ+uBMwvv5MDWBUwHRtyz0p1SXHqoPJg8rNMwA
8HkGqGZ6reGWg0U1rhVOchRhV6n9zxZy1h/UTtPkz7mv0ENHeVAI7aHo2BNe0+br
y13OcKk2BoNiUbYNomDQ79fqJFWwdkY44WPsGWzi1r6hoHXMznCR/8RuMAHrxhTq
JPkK0j9SS3AJlx1E0QAkuRhkwwCBQuhbvVqIT/YnY9reIPF+ojXQqNjqbwhnUkqF
s/udA9d6YqcZiLR3649u/TwcABNoqeoIsYAFtfLQx4lejgJ8RYURL5v+nMDNQSvD
aF6/AmJsV4eC66OXaW2mukfFyJgVIDn+e65LaS8kSA/cUHokMJQXmIhFuBzsBC3l
mAEvxB+QLBElkdmjsNEGfl4NVTCaJOK/xEUJf9Bn6jrThqe+UZu6+ZXOruC48kuM
QiD99l8Vi3EcsjGiX2xh6scz83u1SnugNRvMD3EJq9dIdf9UHMsLM4fkzZO5l0PN
wc0wKEHVfLyZfn1U3yze9+N4SJYzSPnzM1sO8S5OZYN478If6RVjrH6J6+0gPiUK
z1OBR/h1uueTiaG3fIHnhjV/a+youU+j6pR5z94aFOBXvv5A3idW9KlonhS1tKEY
NZuiFrOjcCa9yBWhI7N7yGpIvjvqgT/+mArbE5yD7K9/GTK72HvKtgnSAXconS3v
1bBT0uNkf432gD1qEoQwCR3hHJXCF4SZCuzcfeyvlwh+QZYMFjiGllMOr6a4DsV7
NAeT98p+TOlTnFiJFqpRf5XKg/F9GLCTYkdkmc6aiI+O5goOyu8tWl+8d79LPNX8
FVCq1A6bJ/LJH6Zhe8lD3nxlMhAy315PADvRcongbNK3Bw4RjztPwzzw0oV5YW/P
wBohiVa2ISOvcoeR0mzOoS8qwMDCVV9QnuGFKJmwwz33bdQgycfhOEsqr6qbjo+H
ejxyKogvRNPGWVVQ5BUqBKLKkUk6PiKkOkVi66uxyVUFfchN1IFGID1zWN8PWfjt
L8+WGmwfjoPLtQP2p7+WoVNBVDhmEwIkS3ekPjHQPO0XkC2XWXf7scpSJo5e11IS
exQCNxoazlVDa11q8r2HXBh8MblhdnnY8HsKTnJO4760xj9am0d1Bs86J0UpzCW1
Q4p92TiMN5WNVw0DvVmBXKqq8IWBoqN9sggraUFUeJ/kEo+W/mSOgmq/Bo9f9WP4
TsBQkSs9y+foAqgbY/et0o3voyOGyHZNNb04XAb2734QAoU5OwL//n47dYUmSyUe
Pxe6kxAAtDZQrx5bnv+96LKC8piK4v1r5weVdaxVzcozP+YSyRMLikMTsbli2zt5
AwavO130YaFAhRge5LmsiIWadPdt4kFB1R3phf5wT3jHE+j7dDT00y4ihD/8jApl
oP1ZyYAVs7LmPl93Brw9zzTOoYn5i7xm+t7RCGIL+XghkItAUKQmi7bG5d+0wztO
0pVVpYUyfYzn542wgVKrZUc0l07hQu7ljc3pzfw/9jyYS70ncTgLkck+WwLzkOHX
Lk6db6x5P7KpYs/kZCQWnJKv2kR5DCfJoSaJyOf/8ph76AiANm1qmFxhF4LqXl5p
P3/I649ZrlnsElvic/fjzQjnLiDge+GZS8XftEBn1WrR/0BLTN/mYzlq6KcVHgyT
OScEF2WGjMvhaN60FIhgeL00X0wvSofmJTSG4YgmnnoUyyKeI7aHYl76UlynyXrn
oQUvzEKQypfb+atXpWgRw77CWgBzV0p1MylLRD3CHWEcoWtkZofGWUp2wwsXEWnY
vULxRQely99SQdYKIbwZpS7USdZJL5WgmmxJIQK7moOZRtXT+eH705QkscOoTZdr
BPY2bTqCv62j5xjehLYcW/V+sMhdvu1BD0dcqHdp5ETfHPXZbGkQbkx4uQ4EayHM
AOO/0aJv4J3pqnaPMXyRr2tD2EfmcQm0ETOi6S5kCP/RLlR2bU1zmfUED9RGnGbx
xOvgLGkjTqH5dqZILTaF33SdF9DLvQ4+o+g2nHholPTHVohEXGSxMncrNN1QC0y1
youLlqCf90mx+jbdK0Y0QtIeSs+FBBmPM873usXAcrz25wNb1f8OfM65yItKE9jD
4unrwFv0SxK0Hy5AwwUzRHTVbfUmqCJcCcO0que9CKX8K7tgTInvU6KEqlXeydC2
RlaQjt6CF9bldu0N6IRJYAb7Wcx82/2cXQMCiC5AweY3zPs/xgZ1ji6hHN9xqpCP
kGcKSs/72SWyD3yRq6O0SfuZqPywGbEHJoXgdC9Cb46PTeCOYrnlTUo/skzb21xW
r7JjcBz/zGFsh293yabr672gUQVdjBwMXwn0gifvmg5zMr9ox2gWFfX58zPX162t
+6tzLLmufWGvBsgiXxxJN8ofZ3x7+r0/qe9P2IyZ8NvX8aasOdDZR4rxBZxfyvaE
fBQUTFr8xijW/xe3J/sAcjZjtjQgstK2hz0bbTwavBAg54t1WSu2v8C9XeFJ2QSk
PsdFzcUurcNaEFGvpza4GaCwmAUxplCkj+VufyUBtubSgdYVXjxyO+tDZc35Zh6k
WlY5/9W0s8hEqcKD3ZEoZQm/vjnQAHM2RXkg2kMbYcmakT+dQIRTY7eqlFGxD/67
9w0vcD30hOv22Kc85Q0rbGIzsQB6DUwkAphph0Onf5Gj/4zln58V+EKZhrCfqB2E
/XHkTHRrANy5AJWabLy3/lA0DGzYGXhMs093aULv8xDJ6P04dAyxi4dxEJkN69Sw
wjzCqqPU86HSzDh5P3OhslLEeuwh+Ojp+nYtj22gvDTGDoz9rK5eCbCm2pJECoaa
JwQqGKbWADm4Nx6xyL8YsqcRKwJrpHAGg2l1lTfXRYmpxhrPw7HIN9jt/uS6uOvv
7LyM2PvOYVS34tdlYm5o5z+Rs/cxYQ4WVrQTCNdXnUm5kkWuv51w6dFUywEgcQm+
zQuiSlLf4MCrtW8bILRb6oVLUd8cGVw7jdGUpi6MdaGjo4a9C3PiaBJiqROD8PLu
Z3Kdvcf7TVFXiWFNGiT9j176oEW4RQZkXum4hCxIbSdpReTiZiCfUwpMuJbqZFA2
tvuUsktgVfaAXpYBeinBmtuLdiYeV7SbTY+pexB1gAprNJO883qpf/8j3OxU4r2f
RYn8kI1l8q9WH8yUZ3mnm3MTxbI6o3JrEJXzCatzsVnd572zxJm/ziX6cf6cCvdO
cUsQYKBGed1ajRLE8AyKneHGCY8lx3A0IwCxct6angbQtJAf7h8IxNY51acQHU7L
uVEaOObSOTviLoO5yNBECOtavDmfJtDc8QDNye/QVfzOExTA2iKBdR6xXe+feMQP
yS+PtF9xo7GqIuOWUVmV7m94zxOJ3N8WS0MIPPIa00VKvQHW/yC9lVx0I2Mp+pM/
DRpUFuFtCp5zt0Xwk/9+4a+Vp+8uS+ho/lj0n0we4qoDrcW5FN93piZjghUZcBeH
S1pm7Z3LYgwTxLcndryqT9LewZJsKPtMKbrBTPireMO4+qQ4RTcwV0S9U8ubF5Dw
QEp7ufdpReO+KS3JGyvYHQbFfN8buyoU+Pbt5wVSDQOFU/KtYkplBozBBAif2Jke
h05R6my8nltLRsNiM6D+VDW2tlbC5ux+lKX6stjOJhQuphheU7PsFmg2BdSOQN4p
1aQ2oiALR0iTdVrFzS3a2Q/jN5xF91lIlHUjfgo/NKp9vmP59x9RD9HgoEW37xtN
GYL2BWBZlykCJ4OEa1lRiezQAmAVSR1m0juXZ4iZpX74bPvO5jHQvwc4H0SPyuKs
jCm6Ix66jwKRfjk7KTe6vbEvHj6UPyi9D20t0GabNPyNpt5cuyH2dUPWenmxQ8Qn
NDjOfYaR+EimxiGbHiNfSWNt7SE+icbSW+u/FAzzNiyo0aPRVYLuK4l0EEk4Cvk9
pNtTLbI0VhX9RXVOLVbViJKqcxilJ8HAI6/W5wpetc9jDkWxp56ekenhdzgb7Yzh
0C4sUmuozZAtZddhRQKO5ocNMfiVlPk3CkHs4m90LU2YbiPvocYeAh6v2QVC1eYO
MzGbP6K5WZX3sC90edbhov5S1BLLeeqPs4SMbXv4BF5fBAn93p43xugTLJic3NcA
v0geS79Qa32B8zMcpANkGxarcp3TXZ7f6RsjwmCSuleXq4bhGiD5GLKeiAbp8nzu
jzx1fOBln/m8JUHVs08p2htoVDKYRq8yojQH3YJLGJwcYjlflE4tBD/IMKcreksY
KdjJnZ1GquyjuZi1uIdw3V4ZIDij+iRh/rB+3m4z7A7rN25gd7kJ3WL+EphI51PH
1cgCk7fwJ+d7hYoUf1b2TSZNUZcGyPqhZsbeqxuOVk17LXXsPXzMgDO9LFpLqjzF
zsKKNsdonu6idpwnDEarn5ahB6k+p50OwYkmF/oEpQhYydFzgEQ1qo+RCvhMV79W
am15icC1wRUDmtE/V8gIBXisfP0nprJWRyXr6n96s/G12xXw231BxqePVs8iCDQs
7qvuZ5fFMw/C1PsBtF5QbA4zQ40CJTMAjTR8mYgaovTkBBPzLniNHIc+IdGw7V6W
ElD7pJgUNvGcxS/enaZQp4VqYE/GyaSumQcfbV/Nud2oJqHVcnDLw/ZHzfNe6yGB
qk+GgasXWyMzII3MZ8RL0nCr5HKZwaHwrhcYd0rtO7dSzf3IsfK5LgTcT+1s1u73
Z4y8HUIaKnTXE+wyRqllaKzrtBQGLIarFPGQLCIRyE6YDLLECGqjfx0YcbD2Ywj/
cICAC3XZaVm+VQMcXAOIX7SleYNAGh8CsSuqovuQ4tjIvkU+e15jzOV8qLYNzYD8
0e1v/HegvskG3nJJ+d3o5mClLNp5GAj0BF1zaIFJnv6VI+CgyT3WID4ru5Usvpwn
hij4FteeVtQNzwjoZBiyRzC3At3dU/cJmO/Wb0qAJp9RLQFO4V9ApxNhFA+84d0g
afMKvq4TFcY141/Zj8hKQ4Z+KKaNG74EugRb5oJYQlMzuQfsYtMLcVyjCQY4aUz5
9nx6uoZgYRJ60oXdxItjwE1NYm1N1MhVpy+fPe5fDNq90rWbii3zcivhUu30SqpK
3o2Xo9Mnm5iKEcNyjFv7qNGANGDulT7weNZDFRBbHDv3pPp6jgtGUFgilSGS01kC
7DLAhDTN7YXeH9C5L6L3j0JrpdVyP75A80f/q0cp+IrtV4/oiNkogfMiuU0euR/v
33kHutNK+/j7qnX5MwaTeVlfK119HLtk+obSgFKuTcPmgXzMEo9Xusw0yeN32AD2
4Uly9ylCi8kVsNktyy8r/3LP8oHb9r3Vul2gbtQDOIViFO6sCrq0r2u7rq/+vuu6
XN8A3QFlSwlrMDCceoTwmR+OPeoWMGu/LfORQRHgMrYroxSI2at5oh1mkgsna8uH
KKbmcD9dEBbknM0KEBfVhsOODpWv4/b6RAZfWMUWGNmBvLsgEwmGetlJurSOERsU
4KIMWwvfQNHikjUaf8Zj2DuQpDBTbh24YJQYnJncH9uZvFTe3b5SBsNwPfLIDz/3
ymEFFSexD+gPzRe0gFrfHD95CYGrJ7qUeEnjz8GO2MScpN8217yHA4F3r24LLoD/
7IkJN4EuOMRwnNJ8Ml06dL0zRLU0+lUt/SD5j/AOooZEM8mL/MT9UhfoKSCJzrK0
it8XAm3QwIRnioHg1fRt2j7X9fgljcfkWp0W+R6ckikHTpMQqrS0y8u4WTZtar1p
3QYVYNkgRAxHb9iI9mlQTIN9O1n/imGKQeVMUkalNUgAfG3yTyMsoVvDdm39xE45
4mSatVxDyaDR5JK43yXh3vgVH6p2i7LXBflFIyS3qTPpAOf2qb90o2EPrj8+//hG
2FDSjHO8LbuLqlu3LgYTrKu32LEhs8hXv4QfPI3iz5+rY/SH4r/WQOioRzEzyHX2
WfWPZAv+JBXfq6hkq3QV0FR1u8o7CLy5pgkqu1MeD/lH09Jr9m562O59bNp91Oey
e66apBFsJx5bq45h0t/aZKtwr35TRo/OGj//+aG+92Hm1vwCrmQiURHOiN+PpaUG
6cDEMUgTfXrM3SG3MW7lef+MNm8mt64vfAd7BdErpXDW4+xvtxtbF+EXh5ADQMky
7V5Rlyn0bhP3PEZaRLW/6MvTa/sc533Fzk9CXDPrys1DUxEO17rsQOPfnGNlsqlG
EOkiyH9VVBizo/L9ZMx8z0Nvl+3ihxRQOw+jPMSdmaQl6v9ZvbxeT1A5gcNc4Ezw
ZherQ8z0TLiPkcQEfLdAM2WnN/LtOJqarIOcXUYXc7qCpZQp+dwZAu8KGZyot1vY
+kbEmYE6qC4X9eCv5BIV6hNk2CCYoYwoY+mGHYgqDDiWlrJJtAGo7j3ILWqGoaZI
VhaBE+HvzzxSBcAjQ9Hhw+71dnZm3Et24ugNDkLjONO/Ylh8vJJLu5RBKo74iLU/
58kKo36eXJ4vUAObUE75O7Fvaj31/8pSlqOFYNv0eWkbBJCdmgb+lH7JMtBOU6XZ
SnDQl3XPXwbpiyfG2fdHyZL5BC28y/wCEeF60O0NBaDFP+IHA5F1jf3MFkKvKAkV
GH/7kZw2QI3Lw9Ci0nktMpq/cgXuAJUQdRTKnDiOM05ioJ0q5KOaBZCb7Mx9J4if
x6oJc1PIRWHx0s433y1g9waCDloRi3p0eyECLO3Sv8Jg8wIo1MMI+QvJ8rrFHt7o
BMRuOZwoww1jv3JyMEIcq0IRd+MhHhXA8wrvoMd242lxscSYWr0Kee4WvYoRNPoF
mzhpDj5DKZYUUpoNZlvmfXUbNxG692sduFs7nHDdys9SWUQGAFNvPAO6QDWRvh2w
AMaXn+3uwdyDqgpHdJttseI7kt1wNqItt7kpokwJFJX6B5+XMqdllDUHojz493cy
UcOOrfqoy6LfCPTpldb+f2ny9mFY5zNYrUJIUJXI5H6T/xoTeIbUnOnsMkoVZDnu
/HiLV045aXy6sk0BdwNhTd3WHgAE4F6Wv7I4AWcbXOiCbwVHSIKCMFXAp/A7uM2Z
aveNm0Fno3/0BEjzP7QWg5+suFLPrhr8g5gCRcTw2ZConftTBcYAtAUjkvMMr+op
lDOR3GoEPP9MsRRcRGmAbkJvwQVfdoVmBhm2j/+zLrfh+UUl0ffVXcujYf7UQMl0
zOHFTZM2novuUGTbufEod4WHroag7m3pjVFlkukWBIwq5uTtfJVGkL0+vAcJXmOz
g1hUekzI3IKzIzcAr8W1dWjiGOcfuGWmVBF6goNOjb2hCE8XZg6A0CtwRKOYaSst
TVEZ4o6zc202pjxYyo700ZjIfNpVtb75cD3thBmvNWwRen7EYYyPzavpcXI55NXa
XuGsBsWqhkm6aCFOKbFV5fBhDX48BQoZQIDXqK8cqWWm+cQzmPsNqlbeVOpYrWJm
cSUUH0wQkS2j2wqrJ1bkb4YlGd1gffYpqOvucfac8LBF7EBf4wxaia3OXUgKp5QB
aj80UFw3TuFsmUR448b5z/CkVsOocfKTvN/7a2fDWH685mGX4HK3ZADViF5CUDai
jM4VJLMWw5qRqkHfaFTjG6S8bByKLBef/aPuflqIDk7UiLyZA8vkC5nr68qV3CQe
Qi6gHSakC5OH+3W4Y6PzwM2WhAYrZ8Z90ct0+j3yd32fyya1OKYzDa0/KrHF3KTA
2sliGxQ0PDDcqU+Kkbf2tcg2/5hoB0ZgerFMdLIWBFs54GI6zWslJ7d06gOiQ9s4
Q0LK4RyY7jQ3cSZnM+kwWWjewZhtwWcDaL8jsQwq4v7WAeHX00u3fRVoYplsJqYv
ao6ay+OiY6/t+ZLgD/5OgVc25xWuVfQM1crezt+Xf0cn+YkiaHspRxYDCZ6z83qb
e8X9c99QoeZzxp+tWqd8Or92z7jeQMlgUKs8BYc4UA6tYweqVs7Dii0Mj/tSVSCc
mI1Il5Bym6lHMYya1aBwcp4+gqH0AjxNR/3IbvQX1O+ajYCJ4KLisDpmGYblz+jZ
FG47DG4EtpX0jFq01AZmk9jY5aCnhNv6Ezb8UpglUmax6iNzvGetnIZ1NFW5/T3B
Enp8IzCJGZLdXCufSycgDIE+4Uvc7Y/xteydcTulKOYXbheM7tSEfurdTjwWGmne
SRuFdoFxDWttlDiP8PT0e/4SIdp2PV8rBBOiaQUrpWmiNQG5evgfQmnLZf6Cm+/N
K3Z8WkfSY8vmD6LP10qjqF1tKyd9gKUHs/3iikqpXYcY5SkgOwYlwxFwcrEKyMKj
nyg5NTzfsccgy3NVMSCq4CHTEaxrM1h+kXx7mU2Hz/UZLUDUd04iUin4G/iyoM9m
/9vAcmFnotvfHYFZQKS4w4BCGkuJbTehuh8aGbaK+3qM2pKRKNssnLKetu3gAWLW
nboj9NUyan3JTuTYj4DuyKGds0ekf4tOWvjgJiRyk4MCoUL5XuplFk7kw3H6jiUx
BhysHGgAIWlwoDjrojzqHbV2wt/UhBCMCHT9LMTDnS0ghyNNHAF5xutjFgWK5NZz
RmlYX1GPicSQoFpSBiJ8NcAUMBsxPB0QyxFKWPSEPq8zjpQ0QuV5YmkXq3U8jbPX
wz/zJyqoNFMxF8ksqX5jTBA+KNryGa/d/Qwq+Y+zVDZeoyvCh1uloYunzkOF1S2G
8CuQbQi+10p/49bG+TsIOcZOi4eVKn6ekBQjqfVhO0COjmWzlY+rZNy3i1ruDhza
JM2nf5OJG+3xBOe7d4OECCevRRv6wr1KMfqBdG++aVTAFyI0MeVIQw2I3gZkniW4
e8uG1kpfxzPO7ohfnf3lHFoCC9FJiJ3gjCESLC4yqjsFciqfq0SHdRordOosL2jb
LlOuRR3FclzKB26HDnnNnq1Zx5aL77v++Nu8TV4mQRxOiCZuv1/bVd0hsDF4u+yM
j4ls6szbtMmC6xpZSVu4GyVELjG6yg7qc1iwyR9ZidhObZunl/hidYxFNtWbiIC8
A2QYHjWhxDRzzaa4nF6x2rAsA+HFI65rX28pkmTIhXA0iZpUVqR+Lw4hq0ZwCf+J
WksqR/INrp5PG9iGHTfkRlrOBRz9mUXzRjdTmoNv9F3YgWEegei5xSRFOpsqnxra
TUIZsn9IqyQLA+0MSqlaNnlfFerpy01j8XxkYWH7cVUgZ4yNGsWHPbjknfo45GMo
6aWFMAHs6UXoVYrKdEwtVRYMLjPoLZDgErdS8U98061sLcTQ6k3MBBJaZmI8SsNz
8fwTJiPSGOjUS2fusfaOUyXfVgptyQGp16gsro9lkBueFOS7cCQmc69c1+QwEyXL
vMtYyRrKODV9ob7l8uqYCZPGPPx6YvP72ceVovk9zfqffMiUnsEpoX8InG8HLcLR
pLfJUr15opUcxgYPEKqkloG7xYiIsBUxKTBOr41yvi8ZKdFF6lF0mYp/3ekVer+S
DdJJn0XgwgPvEsZdQ3t3wAD+6+f9hct8e4fwUGfZomQXxrGBsmcdByTahWYs/J2p
pQbhqyPd9zlpRawI0Fn+AcX1D/xQHark6QLwQ71HE0yiu2nGTG2TFbNxL5bMQE4Q
G6iooB6wV6MDndI1x9mmzR3hUTFfL498tznS2MEpa5kRUAX2elcUFp46ZLZoSkiI
kPs0dcWxGyi+3Ii2n2XhJltyd4Y81/Y0nwIMMAXTF8ulwB7QLyABgQGHdIIRZCnW
hgRJB/+kCnQQHCys2BwZjtG+mLq2+YIP8Xt97KKbDQu3wrTvENiJ6GfqkBpIvDx/
7z+7BLIrhCbs3OvHeM645Je86kZISUMsfz2Ouf6fZ+zr1IFQdAor/ReXs/53B+Ry
jrzCRkfzEPITCdU/YyhoFrn72EZE9uscwGOoOSDk8yh0WGm3TJkl2TpY451lU0Di
hNOKJtQDdc2gO0ZE7f3zCOfpY95Mir9OJ64B4kQe70Wgmeu7YUXh23jBzP9FMSXs
7TnOBRBAchVsdiOPsU+9ALgWDSJvQ/Ugt9lt9aPfnMfp4agVW10WU0U3NCeUpkGK
NB7D9Sx93+jOf+4+Rkk628/0RXxd76i3xe5Y/4pjhReLF8tafKJBECn+77/f7UDj
KossMTWMK5aNSlDIro5zuCEMT6dkO+jIUtzazwaaV3TWIh3+KGiSlUcUhVXYr5px
g/PR3laRNE5CwK7QxA+jKUjs44/ffxvnORALHB5zZOd8R4Bn4JnNycKFfFmHo5Tr
ZuJyPkyGz7regFbWJ1Nw54oHM+DOm8A9GK+QSd6vqgV2gMSh3jjjtnyHMRpMh1ON
CGKDNDF3WnMYPHZUVLdFeCRlD/0UXY34JvrdOV/kTddeYR67t8XiwL/vfNAY8oKZ
dWjDhF2lBK1i663MsYzKvIozNXAKZzj4xboEsp45OAl/mwMeDohP5PwXhvyaKNC/
On9oNOLJ12nBYyX4GUQuDjYHhsmnVVJiOnAIdb5PETHVohnRKuGwC8rnw0BoTfa5
gfnHy8gnI9SwtuyADgz+Y6hlAil2VQt3SFDWd6hF1lBvfvHBpI+1u4OV7S9stElF
afNwKS3vWyF14k1RqZyAvPxuqmJYC9K6GJefVhsG91d5+8RRAyue2wcT3XBBHm3k
+eyr4fuUbs3uTsBoY8NUJ/4eLBkpimfi5Xu8RQarNNGR0qEdY+ScyYt/jsX5FwRw
QXgiRcrBBUvi6AkyzuvlU/ky7QPlHiZTO0e9BBoV/ereFBJQAZtrPGDMJxMpo/hj
5dQk42ox0O9pTL8YkdgZi/AVA0MYBCtZTm02F1ZohOy+C8ClBiqjSnnPYeYatR9T
UDxoKGYAiTmDKWO87w7g80qAWsnf51wu9kVjbO3njXAjOrKrx96hhaj+yerE760I
bxzHhsVu1JH14RT5+cm5HHN+QhPbJkJ+UWRH4Qsw4VPhoeTCI/vmaxE/3wiskiV9
mgljHdVpdZduEGqBjmegpc2U8EM7ZXO3GJfVsSZhYqYLzgasI02iu8OrsDaGBZS7
EAUJomI5eJ27gqglzuVNyIW9uwzRHBfSGkWNA3mRSPNfd8h+aTetLdxcTLG3pVj0
hcZC1PbR8cdhhzue3JVNR30/1Iyd2u9c9oww89TR5rKtMXv0RBOO3Q/2RKMlrk5T
nLzt9crC/DBDK58tcO0fFDv/zEsJLCrogI86b/nVjpIkKGEJl2bQ4NCwI5diQV11
kMohlthN8NwobS5+Wy+Ck+myBaV+zhjJCkRrVBtImTjrSwV3YMit4E+fEittTQWS
EM2fgdhQlPybDJsNy4EIPoS2tzl1Z8XwX1z/DR+57NHhQ5h9o0Y7DJGLWnxE2SDs
a7T+zD1xEV0FNgO9V6Mgfqhr90tDomqQxI83SvISQcawXSu6dr6aZyYJ2IY3jX0f
t4fNiczctygPrTNvUqS62zvT7ibZRZOOwXh8/ey4HPYQarF4LsydgjkyuB3yIeqB
HVx6qIEqq/JYdjo0nCwzgqKJSvkT+hY27kgg+ofWWTqiHJXWZUjBm1FvJEhyarBk
8Dwej0lZuagT44qB4Un8CTILDPiU0nooKlmg7h//rlH6Pu+xI6Q8qtKtQl2p9a/v
5wB0a9zm1PNO9eQ5eey94uDSe4aYoXfOEXZiHWSEQAjXl+Zz/fqkRwsMUcc+goED
gDohyJynbN1XAzr4rpKHj6tnGDGObjUFw5QqJYYehXX3e0+wtlVbb0dKUVyzqWH+
34VMCtzJPu+sEdD1L/VJnFAdzl/uHc5nMaYGj6PgewKI8bXeuqfX2n/iVGjcHZ0t
SP7PdbgfDx2IcLyuq7ae+zc6F6kBIoqRe8kkNU9u5VOVO1ewXDdwqBARl/gqOtri
9hYyxwar9JDuYJ3CTdAJ6XK9UgZFdQUYHGl9R4Fw3NQolheGirTRCoNPxu8jV3nK
bTjSIKBM3x1Mclp4stnuLCzz381lDQYEgqZaif0GLNDW1MgQazOGadnNui6pyUp+
aNR5uPCfHP4ZtttY1rZeuP0ZUun1LvcDq8z4pXhyAgD1x3UAI5Q03EJ0P3FigFTG
nuT8Y4WGlTOMHF56MPZzo7C0Us0g4F3LGGvCbRQIPdzEDy9NZVnKfYtYcWJ96XpR
6pZ30A1YdWqtCST6mRudAyYfyGSDuQ8jOLQTu0IJPj+y7Nh7okVDqvrbbFXiHYI+
gL4JSbuxIZHEo8ch8napjQkwvohaLS5ScRJYdbKneSxESw43lkYTxgO2YW2McBQg
AwVOKnScgla04dUDiO8ufYbXyWD7r61Tk4+QBvv4G9jt21yrDlNPi6SMMAQN0Msr
f98TcMaPX1gWeZ1X8AXLEl1HkaZ4vtu3hCLhLiprDw5Yj4A0GnX9NlGfofMy647P
Dx9eQ4pTFW5ius38k1LEh+OH0xhAzVUbqVCk0/vfKlhaEIpChtB3QSwmqsPLGiMx
GomE7zCnrKucYqgWUb5a199kdJVvC+L7fiGnLKEslxOgGHhkizDZeIVzMyVpLvOf
x7gurRVvR8Kh15LszDmOq96lpnQ4eTqgRcCHfMcRS3YjkGzs+4ch/Yqf9sYXJx+P
3GQuvmdyL3aolrQhNYcJWAEGIunWlVIGQp5jjcRTwSuhg6hGbbRiUwncij1QDw0r
gZKAgXJxkbW2m3a8Iy99Bv/XDc9HUtK5AKu6CuU5knIj0sT6gMoPgEjkwOkT+w6R
oC4acdCcyMtZn6cGPuqpfebj8+/3i+xlirYlnRCnqIAGBfcGVjKAIUhM24iL7fbm
zTL4eqA85Yhxqbs9MBZLdKwkex7Lbps2tUIQgdrpAun4/T7Sn1iRRso6CEb1+Hck
JRxJVR8v5xSvgottdXIDfG1Pt/zRuozIiZd359lDzPDMw3f/63uIax83ZC1TtH11
EgJhxv5StW4Dtfhhrd9NTMu5C1/l6PKqh/gh4pbHaXKT/fKZXVjNcTO9ZZSeQCWc
JfhWQL5/RDO92q4eJvjg9/3gZZ0AkW4YAxdP4+9AYfI9ZereftWhTZZDlbz8hjyz
CI6Y3dCK2FlOM3LWNcMgR4YZT+GpUIsKKE619djPhDwfwzhAEpfg3Mfx5uMRYFRO
hFid6DpGCQUL6NGCcp7bJIAXAlxam/6grOrQ8az9rhmI5uKhakFCnC9zK5YNHeKk
uBdR55xTyxM9Z8sazsEW0+ZwWNeUfON6bVFwYgPLM5kpn3BoQe9tUSMDvRrwaShH
/YKJmQraR5p6QBQWwdfgE8arWUEc67e+mZsOYyf/Ygz5QAg0t5WcXmO0hxHwrTNg
OBh1vHrdgZdfGI+Xst0OC4Q59HNQafkoGRxvILOrpf7xdU6dmjejOtkwq0YplIbt
kLYeW/T/EQ+CdX5P3uTkBCcFvQWATh3owmnV2GPg7xylv/oJm1nFhgvPOjbf/b5D
jzfduCvR2a9KjVWBm0PHy9w7tlXIM2kTeHqNbZ1LsGKUQ1BsMRMpgSMPDYcc/TBi
/S5cBAC8R0HTJCWNTayOP7+r1aWnxNj4PUlH9oAAVAAaGt2UbiaBtOPzAPSbZDwf
I6+8Wo2tDdhOJ+B91wjsm+IHlNLIj+dOjR3QCioRz6yECanhPOhwz5txqGYIN9WS
McgI/DkY+YUPK6W3nADa0VaCjctEALRQeKOPSGx+y+tvrmoGEX8DbrFzuzbkrwP/
GjtUfZ63+P2q3m1dg7faMWkcsqE+gosnp7rqAKEzmdfejh0F0p4pxLdEc1X26IyY
FRIwX7dO/WAHGStCrYoRHFFYXRnmWmad119O/y+xs24lUgKOdmQfUa9trIULs633
oViY4mvUN7Gic5Kg6iKG6FjAt5ERIQk5uscyrskVZUBnXG43GJPk5rBH6OeUndVW
ppGQKA2mU45DlNMZWcwGICWRciwfPAjZJrrkPzUTOGS/Yf46PYvdbmZ3aQB7KmIp
KseTIwe7/bm+YOCPd9Q12bMpRErTtA3sUTMTwZaUg90FQYDyj1XBtOzODayZmoDF
LpHyq6fRG2nKRrsw48V6sYcs8Lab5Zl9RXRT18wll40vCWz8MvzNGf/9zz3Od8sQ
+QjvceP0t50OYBTfS8xrBP+aF0Fjejx08vY09S1+V4LafEH21S/Q/zhbrxObPCKt
fs4WN8legm7z2igACz9jiGSwqoHkwLsRk6CIJu4hFiotY5eCr6E4nrcJXSexRy3I
YdkbbxlAN8iXPfGx4cIjj5ZjDUWPuoUve4tTyAEMVpfwxAQPqCDn+jIBqjah9+wC
9xL2hrZP/TOR6mFGQEdW4a5F6uA02Qx2XQ5byq1sWYVfGWfxUQHbFTvGgE8SQ1C6
gCSDZVM4NU+WZJ39uH2T+S+oFFT46bLg0vic6xQo43QfDyjSQdem4hRK41eLjrs8
YSpyzL6DMt3BgSrf2tqLMzBJ8ezM8S4OJIcClTqF1N4VN4K97hbWDl7oZi0ORA+n
vnF2c9DZrVtFD+65jut448zLnwXmcS2MpufgyGNMTDu3zw6ShzN7PkA25VSVCddh
2e5b3NkHNjnC0zPDX7vVDnSjh6Z9UiuAQ0O/mGpfm1OpXTEjP3SaWoV7TWk7LfJl
lgzagIAzYFkU/QfrqioEdxWG0Cc6TN7fC+O6LYcdrxNVmJi6ZpL5ED3H0tcq8dC7
25XarWS0+yAvGKXH8fRycUKhV6DRp57zNSsQAmGkhUR5dR3UQ1GAEdH9VoYaRnW8
DCz1ztJ5+ZYfofVtu3faDVZawUlRxQCtdhwFmI3sCbtotqsFa2stodIOfCc8nyI9
DvXYFK/5CmZJ4IshnzAYlaRfnEV5Q6YTzIDbq7y9gYJi16gFwWSp4c3tjI0I5b7t
XVkgURW1K5xFh2Es9B+icHoMc4/RTJrb9Nt1g8e5ZI9WURP2s84UV7qi9Pu7Gtoj
HZPBzdtg/5J+ktxB56zxgTJEf+Q0f7FeWct9m9mqejS0b7GhC1kBNGb0Ondo0Dfu
+8w8jkqJGxyAFRJR6ZOvn/PCRP+Qr/FtGW2X9Y14hEQAIJ+LoZ2M+FhN+06q759i
sXESfkb3fCEblvKFE9sHiQ2HJ2QwtOMiIUbJ5jziHGq1Y1NAvkQKNj+D7qJbRtwg
vHnhB2Dh6Ce5K41OZkYFyYiyynmxmOI8W6bTn4+F6EnKQbDC+7lbI8hBtKXbbe9A
3fDKj4ImiBiYgq66+NpSg4FJXMHhAiL5rpKvTu6vlhNsaNjvyo7eEj3/expUam8h
gvg5uw/PW1mHDZo7LqWxTYkXfZxr4BNxAhmKydPtERSLJxZmB1VwQg3ZvQNzADJH
SMBT+2xYGUqBJTwqRpfRKOF3Nyples6SiC00A6svaQhF8ZKrw2T5frLgpkbt0jmJ
ZXP910iOyHzeI/O8tRDoodL7/RuF4ZnqOezWFuQxehog4HQh0vIIZgWW9sp/daAq
mTrrJ4u90vLqsWHZv//ByKYIhdciMWEcv1liJ8bMUWEQDcdXT5FlPB2ows9axfzs
0neZKIg7/w7zpKw8efGCf/DSZqeXWheuaWwAAeU8s4wsBsSauJ6adrC07cake46t
RqPSJsytOH5FFqSjgXMV65W5ddxXsPnzTmKiQZRfUBeHVQuzKyvbvqZQXR0BUzLj
1KwOuxRq3UO9+r2DJcPgDod/JCeU3O0jc8gUAExuQX9g+PHycAfzuo2JgIjW4T/5
8sFJctrAeANHfzwHoSxc95TsHHrLXr+7FMBmA1gIkMqurVusU0m9gcJTW3VIuJHd
4CTLfu+3hfqazjBOl3DiGzEzLD7ncG6lBcrob2H68wCkXImOl9d4RtA7TVUtmVgF
w+4HVocTqmCtEiWrvTsyZrcF3nTiXJDurZ1quO+hpN1o1loPSjy5wfrE+dmf9Gwc
AR463nyDKiL0gFF6OnuanisaDoT+xquxJc8u1OSV58Waw+qrHMIIGis4BVAib0jg
dak2Q6hawP6HfXkNNimIPymwF2jMSrndj9GWkk92LDWVZOO+6cTNySiJ87/0AI71
XyGN/qhg2Opd+c9KjQzlan5nlqpx2mdUUHWhVjdNGC/p59kk3ihb5tq6QDfP/PD4
uV+MOF2ZhFshgcX2dnEYQdEnCtGwvlJ/UDesf6Oj/xHFXIUY33JNokOxDZPqXs69
bINzBUpcEoof9C82BKcnSSDb+IASqJJQFs9eTxmW9wIJUCrBLin0Pzausm1ujnSl
r3bzI6JHGO9R2jt9esIuBK42WFyMt+vC0aug4PxK3DGnScBOe/1VIgzTl28Zt93V
V4JSYV7Uxa18VnnXfxECVikTNXJM1C6dczmlFcTk12kokJl0fT0uEYUuyBtEuMj1
VXqKYwaFezIMiFTfzv7DdNE24wKTOZY3vWN0PdsS1huBbnfsd7gmYPIahXailK2N
ISdxfx6+ub0EU9hwRdmycRnGFHbyfZtL/gpTlgHrIgzZgzhKn8rFdM7EQDVJkOy0
xJXFLSR0zAq+Q42cndx4r+mxhK2MJc9v7D31m8OHF+TnNyFn6Oo4ipekd8fI49V4
Iz+EA7GJf2tbWTH8Cx0UhE5OUxY+IldGfp4367myI5Lm8tjGTPYIT4lPe6PmsEzA
sJ6+R1tJpvP7BqjNbPoXCl1rfjhZ+cT70HmT6ni/DuwZvw+q3zNSenBZtj59KZ9l
UVi1RX73ryvE5OmE84h8MsQ8Yc667T/6LfR9U0IjukOKcXTyX8bD2HjgbiMBDFzv
FA418/vXsgOmA0fpnupJPLFR77Jjw+UnL9OatJaS1oKUlK7VXApmJcKk22HLLjNT
/aaTlnPBziIWsAtRjZUSBP+Ay8wlKDcBJQXPIJmb+gJrj8jZD9vfYBvrVcr2+mDO
MBY+mgjHCmwn13sfmk/0j0ZMKdMZazy5FcFI6lOLoaPzmZ2h4YI/zL/4z8AEWSAL
JGgero4/113ANzf7IiVTp8+UP4RsoFvvaY14GacU6EwudwHBeZeh2pHpRuciRQGp
KVAVxlj44JE0WaSzluOW51+X0bspcJn6ABtQa07oR4P/XzuwS16ga0B6L0FtbpG5
sRo4vvSHceJuDgjJGNehAmfl05Kin23wdb7rQmbHtUCkQ1vO/tZSIIxamH09K5VV
xTWSBFE1WAsXIFxfBTPd5TXHT7pj+bRlvbL8g65BEeOqM+yX2tivAtpOp3Io5ceX
8Rk3VoTwXKPHnM69iOK3FLCC3gYlctTfRfiWbuAoWihmvVbqI6Z5SlKVIz6+AWe9
s1XynfQJUtFzu+FX6tIl94BQCdC3Q/UlQAr4+equRWU04qgzzKQggzHqxXTqlLUy
H8gudNvakletVGlc+2+TRTF9D9SRg/QurIZ/2/cBB56uawjX1Oiuw7L1rhl6C315
3bcLmnuKE00wqGvfoHkwxh9owKRT4JFZ+DxDyrTiqoy03XZ2eZ9bz+qhG5eJYP3I
9RU1lt907BOru+eqV4wvxIZcVoTHkwDbSF/EIPwIst4gCE6zaxHfj6MDB/IRq8XS
qIb2TMtvyJBlw0QbiDmhjztEjmFIlKRjedJonY/3k3nuyJ+F0AVCXm35UAr9d721
++A4od6/3URv2x/NCf32y81IQRcudvZUMq2WYdNDyNuuVzzpzKB35m5i+fBkHuiY
buuSAsgejuGNZYIGFs4L6SEBvReHVMvvsCiEGLLFHSmp2N4uIEniKrVYxpxSH18k
XDPaiOJe/8qVTXVkZhh40rvADgXxQbVF8hWzU/6MBYRhMz7PSrEBB0yUeykFjK+O
I+MgffJ//1Q3SL5MnLyWhRaJKhTwZBl5CkuVK5wzClKNSn9H4vw7pffZXCUknw7A
AyYhP/h9vSgZBev0l+YUk+rkFkBf5cKuWFK7MMUHz1ivP47nb5T7DeuS/C3mFF1y
sD0Gu8CP6zgtRC52YI5cHSvxBuY53wiRRl+zVTrJkZXE6kkcbmlswvbp9qCrZKLq
Rmavg45Qj7eqJhRls/2WmWhMtVwKesE+aOUt5o8IOqK8Rm0m16h6Y5IOlwWnT348
mEhwSJoeX74I39n6P0CoTDVfrDsR8GBkLDQNrw3dHfx9Q/WZmTzA+lzdLtk75MyB
dhehCAenbCZbXZo481kPXin5f3FFmaIgEb4XWKzANgTo96uuBCLI/7AbOiWUmsfZ
ovBbHbqw6+ssv5+6QynTFJB09aB8OLOmfV2qnYY8jtpAl0QMt7gjknc3QqqBE0Ka
5oaHl4SFW7hW9/bKnOrWFxwr6Brc+mR35WMc4cVleHDThqwPUv544Wl2sIgDSdFQ
pZEgd1jog42JIA1K7bpY4wDxNzuXBvtYzwhVYbLxxP+xTzI+1QM9L+9S2hWUB1/g
mdSQY3VVuI7fLXXnByds96wSO8mAFR5YcUdXzwoLcWaUY9R/xXm7bYq9MoJ2B+5W
41IiyzSocVV60sklAqpYC//pRbkx0pTFEFEE1O8S8ndeyae7QnBABswB4i92GrIF
WxNqJLMLGgq5gq77tHnOmHaca9IRj89MY9+Lk7+5QYGb+VS6ISkQH4oyth89E0Mk
qdg788byydEmE8Mvr3bAUY6j5OrV3IJyuraBjvwHAWox8p2sx84ouRNz8XHwlzPR
Z5JiA3X5uOgqiD8mkMPlZfzLlzDLDnsDLHsP3X4kQcOpUfGUyuMQ6bjOayh61D8c
HSCYUHIKbeRU+AnU5uW8hEvN5xeqHdRqH6tv82aPVECsUQe5hr6QziYgg0H2s0do
hcjDBE6Ss1FTRTnMlG5E3keDazU3W519W/KGS50dQ+JdRXxU36fQUxkmVcRftbF4
p34bJFFpY3XENBj45uQdI+jzNNPrvditkDtBJesDEURKpKzboiThGrnUddqseRBW
PLbvP8WolhsDBUc81n3ceCECDCvF3XftnHfjtjQogwPTb1T2vBgS0aIiIzKw+SRM
PWPMTRZI4whYQ/SyghgjMAm07sL8ys1XdX0HGXL1e4jX/XI4mspylxBynqAG3SSA
w3RNF+uBQE7cPkMX7Ofi8GO02Be5VaNS8wmLe76VWVS8+66rmH2b8KLho3z7NwQ5
kOKRAY8iAA5+tpkqJEA3tn7vB/0tR1BUeBZIVUV+q/UJN8D73Xz2DkgkQCNXI67N
C1+GS3FxgeQQu68pkICd+P/meDIpUaWYvtyfm2bOyeVLyvIzbI6I2G7MeEFNOh+E
e8dY9RFfjKiCDxa9BvDrn2kC5QcmdgOCjZLHm7xbaxKqdZSGcm6v1hfky6KaFDZD
/efce5oJRRWlOpUbmhpyehygmf9lib2tI+fivS9iyT0fA2TdE52F1P32mh2lzGNC
9DD6u2Ys7//z4iOQXCc3zIsErfTKSn0cKx7KgFvvM88wJkJIByIyJaES6EH5pa0w
hdteJuGyUG1cM9/PB2EhCSi6EvpEcw2jPDVIaBaW1prLMNF4GI9PjD6pIC3+qjtw
gVHssZKoAm9hfeik/EJL5U4gxLogZDhZqBj6Lhfm44Wbi99G1I0xt/Nv0NgSk/SV
iulRgaBm9W8AAECLGBgggttPd6Yj5LRqolYVWMsQMwUOmxtLm1vU8X5aX0XPsy0i
jkY01RUe30DrHdtgo5bVOy3Z6/qogRCSxePHo3yGTDagOuay+pNt36XLdfbkVah9
KT/TJ/fTkfsB0MgntbSh08kx/c+eTD+g16ybcGKSQ5pzUUHi8C/i41zSn5vcYtSf
gWhD+sOytNjRR7EcZzD/h1EReU4DvVVNob5flw3Y1oaCIQsH0+eUl5DIzIoV7yJG
UYNb2BKOs3EiIUZ4x812FtJfTcJTSgEAbnxyvazUWtRWO6/gLy5GIctPognyyto6
3TToiqjSWfiZkyDglXqNSvcFnKofuWc45cJpOmRO8l0P8fEb2dCTiFI8/vzAuBXo
xxgKJMekC88mx8fol0WlgMw2P+b+BUBWGpiRJ5ecWi5fL8s8yiPT/jvx9vhV5iGO
gpyZswz/uv6i+IgWfVg4t5j753s2hrapB6czkV83/He0i2fnc/zetGfozt1z6JIg
Q3bf++NJE7K94nAaKGA4wCrWJqABOXcfWquPpWypEiW7EvLBOGZIFrIHPvHwH/cD
A0IOrOHgimHKW/DaHdf7NvMsi5WtjUh4xU4qLWUYWAO4PTCWNpHFSclY3qczZLEl
7rHGUx+TlQXhpD8rxDHUq5rNzmCbZaUu1Zyv4CjxdF2AzQYFYeCo8A8bd9ygH0Ea
SqsmYbGPtIW89Yd/9oWk9SMNMW3vYHvHXCbtAfRfBUFGk1KXfQKnJjSI9htxcvAt
WRQ+xvFA2cPJeKNCqFArikMhMZlAHHMPjr6clC6H5OGd4lri3LRjsDKXvkP8ARRf
GEdRwB8PZquuDeQx6pyHP3hzC04VusOFIF8JbzSOy5KGMQ763MeQX82XL5C5lW+Q
XtgFO3QeaziP8/PMRXg5vHxKwNe+SnyEjG+W+UBV9y2uwoaq0OvugFjevUtQHSRc
QZ4UF2Lx0rhWugAfaeNFKr43Ls4cy4gaqeADRMjMdegiCZ/7A8JLj5SPy/fXBfDf
xXEyW8r2bQKh9fBiZV6cUU8b5a/khzxlQl7ukPq2ZPi3vSVdQDs8Mc4hBxAB8lm3
KuE6YYP6y1nlJaatwmlolPB1pPZwfz8sIMiwSMZZw3eHdjeSEimBZE3Kf0zk0zEg
EfX45+LYx//pF2qg/mW4Iccm1aSazVMygpYON7P4XkrFpgtrZ3uD5fQFubV0bFU/
MdtwdgKIhSfdQBEkD3k1F0uY9w72QJp8tAVhCBuh0zU+ug7gaeRdZslaeW9kXV43
HWggDIRPpj2b5Fsz9ZqdQYX1+4qHE5uzBVZG2qQl4H09NaHXcZ53aJiTuXgflnCx
5XztPQNYmL8IH73wn8xWzoyFqyTiFUcVCepddVRzdG9hNt16LLONCRHG0OOpWXGR
YWoFzx7Jwt+bZhMQUCkf++zUGpPyIGUJPvopZThV5071nqaIHFQN580FXF4dwDlb
pT6HuyQZ2FCeQ2Dk7oF8QPLh1W2gSCvwd+CgFE0Pjp4BuxjjBXyImli1CEaN/A3Y
rTkz+jm0MK0RfCZmFQUxrVvEOLfegtq+nbzlPCnY2tjUtZEfBpJZXMhKPhopBKUC
sFanZEmJ6PITwEVGr/4IE1QhTnANP0GzhhEPciM4XneSLkKMYSOOXnP3FtlUKFyA
q6hKVY9DH2n1mykzgBRHm6mlyx7mz9Il3J0tj0AmlQg9ryq/m1Z/L9JXhnmtv/eE
5K924Zir/95LIsJy+RvIdzVTGo5BvGwpy72eeiCc+gO+ah0gf9TemroXH4/QFtux
zqqdQALBmzfKVZ/QKNsW2eDtIuydt5ZOjeYDy7pXv7JyelJnsSE8eerb1ioANKsT
1qnPjMytDlVGdZanpEyEB1aPgXIn/D1/XEbZG8zMMuVm0EgAbd00w6VOtOOqYdBn
QDuNvCCZnn4IbWk3Vp1RZtIZ+J5/dp1DEC+PsEob9YWS0or4XtKUsazUKGKYiyxf
B5MqRFQbiIw9K+r0rHBl7+tMOWKmMrMFl7j2w7uo6D6p63PUq5gmi3EHkUfhwlSD
RHciMcGfL8+pjPX7mBhbDdmagkuU/9MRbq/N0giOvFzCSBNdv0E7hCM4vmxBw1dv
YGZhKcfE470fkVrkbJ7iay2qzoYWRIVSa6WC4lOtkzPr2xGPASOY19NLWkn2vGyG
Yfr2qI7/wtbtH03LIOquW+JB6KWFpZpSiAUbj+w9UmWbgnbxsrg7H5k2W0EeOkps
0v0cvv2P5Jmsww50OE940FrHJ11cgK21MfqAgQmzpHxL/YhpKPipAK+cxmokZw9s
wPiPtzbhaXYMLBU+8XsqXFNSKyG3/g8NwjV3NTkardjSjA7PAm8YwLyaUyTwdYRg
7WLqMs1Xk8NEGILuNunx1tZadcccLPVUJ9SOUX5E4ktRQlHT+/0mgZG/un1Ov7Vu
X0Fj3c+l8lhU/23VGNf9VM0RGk7k0bstvk/IUa7As0msxgOUUavyd4OILd/7eVEj
Z7UPXgxWU5/N2D8ctR9Cr7ZWETjOBsYYcQSYKv5KAHtK9LQwhObIQbN/GYvKNNSE
26PzzXFIYVvLtgtGSDd/t8j8ayJWyf5dLnDBcGTbZ8A+9ZP5NNZrmFbSLnC71qpC
7htZ52Q+pfvS131SGemHIhLXBNGFL1vZ0HgIerdTggHZO4a3DbF/glW6c5BAdtgs
2W+w/jw0yygzMSSjVbwNJjXrlkTP6hTaplIuPrJnoxfrJ8K7t8Iz5P5iikxkqS0q
d9HTTNJs5sOZkYQhmGHbsSLFyDtZiQYx3xxeyqy4PPXNZ1ChFM6t1aAUPxbvyUtU
5q2wXbu+m5Y9qb5f4Ds/O9nLn8o+0oGfkOJoIpBBi7gn+q/4+/G2DqfztFyfAGnI
keWAgyel9pjaxkMiFa0dhMuMKnxMMFPh5uOgAhvzCZqBPxqwMarojF2LWo7oXAbb
GBckOIhOkNqW76t5IJts7HkCp2rGTZCLimNGIC8QllEQ7Q454M5PFjm4dYrWyflq
FfxgYUiIcwzgLzqLzjQvfK8UaCATPDrCciCwqvJiDJX+bp7fXMM6pjR2G1NSreJe
JIHYdZ9s2cqfbGFKlpV/dR+VSXqJxZdX4cCJ9NGxAhsWvbBB/vUIzNT5gtxmsltm
Bv+Vcss3Ias59Hr3ozuyG+yCyxCHjJ6g1HckPS7yPb+yzTcMJ7LQP7UuxLErm2Lm
5KFC3uh0tPs9qq4iqZnDGkwWri1j9dCJg33M2GueYAlGfj7tzIg18g9TCX0IIYHI
PWZmfYQ5vGeYdVN9EtP581dvsdeLlIVMj3zn2U9eGL7w5bSMb559BCOgFsuPKxDT
lmRovHlULoIFoUFbtpb2EQe4z2V1WF9neCfJUGLVFWuHc/UFTgOkB8Do+376QsIg
hD2ijXP5BgZ3f+yjt6Z63otRczloA5Fr7nn3aN0LadkTgF9zFxi/P/YXnK2vX8YO
6Wx7jciRjgh08a30hxXsZsQXYfd2efPNMED8GSWn0i+b+LYlzqLtmxESzGgitkGO
jeLNQCcFAiNfQmi0D58Vy5bNhgn22H4zRZISp7/Ukaq9YEBAp+tZ2FyImZRKrx1z
oYLnq3J8o1zOkhnu6u82qTKjRe3fSupBPCz91jwLOpPLbrimn0tD2A8jJEEqnzku
awUPyjtgorNRsNz6Xx7RKqQ5F+6XAagEDQiSRxvrR7khOscGUzldIaGdQcflevGV
ZwaeoAXP5Mh8yR2GAMsSGqzZmNMX4bMhqVzHziMrUD3hslvbZigwDkMy2+adysol
SQOsQpvVSuXs3Ym2dcB7HrhKwMuBwi13RUP+H1aYcLuFpaXvEgXZ6p04FsaY7ryX
9FPglA3QFO9Omz+t7H+xln1uOhjr+xDs6e86dCaVhMolN6GRj2HPwBCFCMTRoltL
K5NX6i4k4QygVlf7BfNB88qDclb5JvzseoBjn5lLs3S0vlBjkivQ0e7F1HLYXGsN
tlWwbbj5tRAH9aW8Lv/m1jGxAGKYs1ZT/Qd+wW03GLN+E2hPnvK38F2pvXGH2MCE
hoWzO7Tg7xiLOtKUXcyo2LQoajpWso7oHnVR8/vkzExGYiN7jiU0cowcZ489tZlu
dV+rwLIk3RkyIgF5w98LboMuCoDsf+7dX4KqNTP71DNk6N1LpLVZxkrHWsMVi4O/
vVbvSd2yRP15GZ9QAz5KAl7+HxKNGWr0GZI8mBARg7cGHSd1nvgpRcNjfsLhr6MG
0BecX6PwIFmzARkeCet8BXYKZo5aO47gpDK/UCTCLF0ewNgq3ztIbfTgvWG54mR4
TxwtW8zCu6wnfFh+VMrHc1VzoVMGoAxcp97cbACf65PuVhCPhkV3YibY5wnfGYXF
KjHjsycP0NjDNeGISv9fyUK6kYYKsxH0+St/vlzU7/7+wftntB71XjudqmTssShH
4tFWcPu2zsXAvDvZKCKsHFj8x1fzm33CCGK3QgOIk1yd1OTxVzlEPV9IqVdlWk7D
9vTSOT0UpxVW+mR/rBcGX1WH6FTQ1x4TB04JDGlNz5VlJd2nqEt71k5q2Zv+9U82
CtqnPmxoymFrboZaYEZOKjQ+i6mm51/s2OzZP7ukM94spAuJhqjvTFdmsLeRI5Tq
QcJz7ZNmn19C7Kf2aqIdQKxv446kGS7boBqhghPLwwVABMRQrZekNA6kLqyAmwzd
gNbQiaL6Bht7IiE0vujlWar5QTrbk+PBZ+K+X4fRQMo7XInocXk0PxKWmA8aHCrO
17zPO5IclcFQmAzqKCOu/VDLllEpqMDD39vnMmooMwQWDNCAcL8eBJQOwBmnYn/7
JaAuksz9/amGzg1LuG4yjINicqZE2fcPuqjKa01pon6PDZSSUYaR+74lyN9rE5p0
ty2dxWMx9HPtie5Pqjebrj9PbuUXd9RoDj5G0RfJ99GRk0g5jMqBjmaBZhT0TmBE
4HYZGSA7o7nNE+gZN/PIC6mMahbEoGqzIR6WeZaE1JKmIe52baNXNO0FfTfzyUmA
n190m86OqEq1sfo6iVgWmHhvwqyDBn7h1BD5HtE2N2IqGnjjCnWL8PhTNUdCNCmc
Qcs7z5WSJRwYr+2JkfDOwVpUXKOF2Gl7Z0b/m+azWwQ+YZvf2pViBZ2Uz2C+8u2s
7zXyqKK68qES31BlQ+QHWaL52p2YHskcc2GqWvpn9MwVZNS3IkQsPylD0ByOi64n
iVieyOyk4eYmwhAJHYPFEui4uPXTGnjd07ZUHmFsnhTTMISbhRvP+TCGQZQNNY/r
CmZ6W0glrVTbjLbyOmQCaS39uNtp/4oIlXvdHUufn9dSIvmDTjbj05DEwNPWCjAu
ROscbR+FVfQ8KVecTR3uMOcTRCLNbXlJQNTIe/J1iZF12/QgfU2NWZqveZMV7Tjg
4K8iVZnVPZVgwaCq/SLf6qCxWxMjZ0Nm14WwIKG7SCE8ZTpOVlidhxEiV7Qajm6u
42q6qO13Jt0Kvx+300nbXsPWI4V+l/d0pehXtaK4mXXYtxxfQ83yE8t06RMrtPjX
FRVnLCNUhuAYQrYHIdNgMHaZpylbBIZkAEXledS+U33LzSs8/K3snrIMoZtTnqz6
B9EMu01VTDmWMPICBXQflGR8C7NLnCTx0So1tVf4x3yeUeb0WsYCUQhd85yDXYvP
ZEi43fh6k/fNf/eT6/8PwU4ww36OIapUnNjutqG5xqui9pg8+owv14xy+DubORTM
nmG/iYGwH9rskEclXnx9Q7oV+Rb+Qrf7/C/wYqzOljLyuuLByUc068p/NvRmoArl
`pragma protect end_protected
