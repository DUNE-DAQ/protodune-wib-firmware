// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qJ3io8RK3Lgorg4IjcuQC4H9wga6Yr+bdv4osSpXoxGaXtJoxgRIingSUdTKYmxr
BFYpBIb5xUDlaj+0YL6BI5Yow8eQBFvg3aG8vsicRv0n0Jh5XYGII18ZZCdDV8O/
G4lSs0vuSTRjORDsQlRymTmVDd/bG/SGsqC1BMOdnpc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30144)
ChCigIAfVXeCpOy95eNbRixVe95Q5JwSrSpJIHJ/yezhCnUXeWnsLKKxEV4+dp2R
ET/1V8czGArbGhzRhQXQ7Da644j/+B5PGa86+GTfUAR/aKi4yEwdRcQc/4roSkSD
7rglKM8jFIjZmqJoe/+5uCuW5dvXYUmIjwczVm+T2+rGUs1IR0SMxv0psgW23yOM
XPMHEaxtncYxbnN9dt0UNneIOeBF37Hv7YBUz0mAlQB+NZdkJJSFTWzdLBDF9BCN
PoeJBqrKLk5tFo57KiS+Dk6CcKbT9NqeeqCrLVMJeq/0tb6phUsNYKr3zkHzbene
00D+gv2flnUQ23Qz6KYOJdxK3GSP8ZLMlj3KuKT4Bi1kiVy7W5qCqo0K1eEBTMZj
c/yo0ipv2R517PMsBJpPxXzxNpNrmlH1fSBKtj9ot9vZ5tIqMeD+fffAihk1FtEl
0eNvgN7zmzlPXIgubaL6wt+2Fe++FYZwpDtmrjrnj82o9DfVy7OnFmqaHb8DqrZv
g7PobmNdCrDv6vkDE32mUrZs9WJtUVOzo4pMmqXjOj4Qz9akPLAUbjtembTAJV0U
xHScdSLwyqDrVZjFQjM8WUSz1vKSPMDAX/5pToXF5ycIqc3DYyIEpPNhUbpNvNfj
H8GimyUCeNSpg7nsMJq1OjB0uOW7eYm9l/biF4doDNAykKWz3fx/s5KahOWEDWUY
mZXwZpTNQVd+Ycsx4Dje924aTORpKFr2ewza+dBOa5flJ4sWt2u6EccU/Gy7P3bT
qsCvVmzxKleGOsSLvd7+UGafLBVrBC9bUipBF/LYW3xnR5uYObasl/g/LfY99Ntc
4/E56O9eXQ8GpF3bSNYbIfQTeh8UxjYzLqlvAVIbkrGoZJTJOLQp25XyqOgoB/1c
bIZBHigqCIJuCQJF9eZ01UvMctjvi7MBGXYPfXsEoJd08tb7q6J6IxAZGLU1bu5l
eyYM2lztDBi+qXEP700kI8kxQAo28tUttZpjuSMyzLr9+UubuIcVvTzNrgNHQahK
17kX09GuyO2E7Nmzm7reBznmboqb6lOc4vOaxBB5ke5/N/mNwGeh5KwB11Gkh7vS
D5dcQRAkgl/Mk18uwxRiu80B+WLwt2LlIrRRODGoRQkNrDVHmJQg13mHXhKK1lpR
QOKLUmZgi1ewwxTlTMpWywD6W/3NzdtX4Jy9K+ybjbNcdzwNzJmtkMst4whcXa0m
w92JJrfrsy+23v7sdMnUU0FidKXbmmBIhVkVBIpkATHXxO0RRuIftT+GfEs7cPq5
b3DHrd6fIHeX3BPqQenFJ88uMVJEeuirPSncYW+sJvQSAENH0y9/+aGzsciV9m9k
+U5O6LLMuP4X23TRhdyzCXCi4UKvj+n78TS4/y/J3DQEpHoVmlp15C6wbcTdibJF
muVm7LcVcHyJscJncpv4VgaGU1ky5CFCWwZMmQLg/A4r4GYZtKAeJsYxuENeKyEu
cw3/n6ymbzeIAkrogWZ43VjbeNiuidqeRQ+FELMPZ2g2nXyuaNezLuOFmcmj3yHe
XRqX+dGhcIlIAZkr8uo7k2Hni2HXR+ajdgpleM0D2o4wq1s49YF3eSUegxlchs4E
V61gpJPg9hvXnHlpenuQZQVHpAT5tYpWhV5y2+5OBhvQe9T1i5nlT9TIQWSyQT2U
5RlwKIQCcxkOXlUs3e6GptT3h+q1ISvk540K9dQZGMzo8o9bScWAXoJglZfh/8Fe
YuUyxCkNVFx18DhzTiEHnmxdPix9ktfuyeCFA+N0DC/nHhm+E/dU+nCDazHXIB0O
6vTD6GRAKEPF/Y8EbKXty5z2hpeVcWboOwjMyiwImRI1A0ogLXpZjpt29HT21XLu
9HxuYkaqlt6UMMu6xU0xHj3XepqAogpWNy6306q8+K1RGHYldD82qd6VW8ip8Xm+
rbUdpmF7fjWrgcBroNNfGXMsBRQtGuHAceXJmi9nec5KDOiLK++wDkJEo+2XLR8d
Ai2xXKyqdT4U2ftzqeHH5NRy5lAyOEx/yzUEj4vFhb16Vb9VZRuJWpF31lsCmqzP
P6f7HwOE6H+eaCN/ySCeCTDGtq99+BgYHTypdPI7Dt04oOUA9iWQNC8UClMzopxd
6NNWp1nmrNeUebCI+hzmhKoPlKsytgUb7q/h7ONGvygoRz42X+I59JqFVnq8Eo42
k9fJEg1C4sdgIUrO8st+pfC7lR/CH/5nfFDp9h3mCcKsgnULGy1UtBdmi9hMsRlc
2m7ovoBtDClxGO2ZHauF9WGH84Qw7PsvWUrCNNwN1b3jhlX2zuT4jjh/YlAjixAW
nuBhrIu0Zh+iBEUuRoUONuupEQovD2FT4WpdubzsEHAeFszlWlnuC5I0RtwKlumf
/aUl+9pI57mfn4CTXxba3gYBi1sJXQzf8Ndf7FXgvCkQZcN25eHuBhhF8IHpNE05
1zsuAdMW7V6CdXUkBJ47Ud9iam/HqJ/KU7kNAR0TNqrBt2Ym3BHuzxXYiXf0Aghn
pd4obfca+v1L/fRtHNaJeaDwsse1DzaB28xycuwp/Y+Q+gQy8cskRBNwExkH4r+p
a4OevX3GnsiPXTpcZhFUI019KPjZLCQcUE9Xjc1pl1waACXYjZVYDOR71hOI3oyW
g86q0NRHTnzeXlNsdzjKkvIZaVJbrAZCximQqUO6ezifQy3JASrfhFUjR8uM0J0j
wiKVkxeCi5CqdpeIbL+rLGP1O0Lu7HgUrL+uoX7d3fVlbdMdD3yB6HakR6mjQ8y/
tUA3EPGGRUB8ECyZin+j8D0GYuEfH389Wmo5VAGSF6diNy6rdOh4v3S7PxOo4jCa
BQ8T30yfsRv5N/yrGEqgPPQp7OBEsNernz7fTrAhO5dBVxUDG3eNzA7uNl4pIJMy
XSGTPa/T4CYoPluf+97fo1pZNhs8mwcS5iziBvazZyWJvkzcXEsHRoanR+4JOGZD
XIx1xotNJqR4N1J5zaFg9IsRi8wJ3+/i9BOupwxuhMQPNorj/EVxtd6K5TEUyyYL
XtObbVBajaZTsygGv6ecadMrvwMEpDc/Tqct8xSkZWOo3D3AqxlNRXOMVFUm0+bT
OnSMUsaUbxg2OeQLZ1KuH5zNCEsIq+fG/iYlitTTBjF1i7vUJmRHka7zGl2drsMA
9/0udCcTqJnWlb0URjVlwto346xzWpeTfc58nxaH6XCD/skeG5UmBX9ZxhWwVGE2
pnR+qZehksxWRCGPdZFfxAkAqvqcVYbEt46Dj4FPv4Ps8+PFuiVgZOayrmO2Udi1
Wdt3pyZS80CufvJCefzHNmYqPobzHn6CID5T2opFDK2YBcHcCiTRIMD2wQ44za6g
Lya/sPo8Cu2UTLl2Z67blDHqjrORXgeGNekV0h5HbLyT4X+8stYp2qUBeF3gFpLv
B8vUF3jMmHJOZEREuVbGqzQ0yaeGlPrTTVoSkuOXY/I8TYPREsLUj2zwf1oEC23z
HxdVHEgpbWsbODwUlUoCoKluozvwd7miMfHup8kjqC28S1MIB2mMHhGr0UjASLEv
h8pkDLXX+MPMf0FPc8Bao102/XmpWp6dakz9MyNnu1GL/MWnvL7Ce1qJXKIfu3I0
mBhxcHmcbIb3Q5S6zLW0iKOxz+kyg4JtXHMZwoRVpU4ADaNE7iEcuIr01HCtmGkp
vkjCYsDW8bmG48ZyCJQpTI+V/vD96yncv6L795oOTZpucxqygAEl7/jmkNwdruwQ
B4RNpzhTsFCSgCkTLlZd1xgYXO4V6AEepKglZKkNhJ1+8W4vdu2FGCqfY0pdZV1/
Eu2e2lxIrqLTGGxeQmfgchB/5zut8Y/nroHMAy8ZrPWZj9s+oHebjYvbDUID2IGG
cBUdPrFfYj7mZEsHPHar51wztRRuAGiKID8R93No+iRcEPd6wOKPbVSRPRbi8Bnb
2eBCu9LeAxZxMEIYsWdl4PIVNc0aPYMWPMNza7QF6MNauBU9cnFhE61CU2VkGFMg
HSC6mi+wANyRB3c+gVNya8WY5Z9E5MPPoOrJBCeTr5u0p6h6Re+CDrsjxJ0G0kUQ
Vibh5uRo+kWoyY1L/Qchd8QQxZ9jSIjQzs76XT3g7lM1+qD1bDDUkckDnp7WsIMN
vrAQCo1ONEo3/PkQfDHdrnSazshH2z/wnt+sitS3AXeNa6knWfFU5+8OG81O/D5M
5glCHOv0orHpVRdAfPqpkgo69SuOqTrP+AWZ+CVlpo0kmkvXpbxszHZPpAdHGEs+
30g5JskK+z7095LdTvSYnPrUxPU+/xvcbljsJtuLHYTbt1BFoqJVk6LloQdvrh4u
LAqgJJy8e652fC+YPiHR73/Ar5gD9AysgatbpD0+p6Axe0EFH97ghEmQjkaHxQb3
TK6ZM9WWfD3WdclvrxMmOrZsBiMFQFFKpkF9P+rhFudLqEchLbTYZnYlqnYeluGO
N/g+FnqAhMws+MSNQuFI5C5mNexbIH5cQtXpi2+KM0nenf2nLD2JyfCZ/wMLr77/
GpYCucMZQf/oP1lsx1glsoZya9ek5fnHRPH72lRQHKa7p6fQiuNyf1tPAhPr6YM2
xJD/Az5oqVy+NPxWhXzHlkoaF5PeYaRUMkOCP8SIlTvxmHClgXDTgq9Edlkl9h2C
1sqqlif3FOGiZ9XK1KY4mqP4a/DYS2VSkflcJObOfKAH64LJoAYr9G3hRn4stI1g
AApCAXL0qz/Z+JGJO8heB09JeK/d0SFHRT7WytVXeuAJn8C6+ITu3wh3VokRSMKg
8eeV94eQ3Z9iFIDOA9oQb/B9AR7RGqwKVy4QsJba90hk0wAIpcqxyjnEE1ccoAoG
4ExrGUa5GKAYmg5ixJ1oi7+Zt28PgcUVjaLvCEABf0iqRKXltO9gz40FgUhEZk59
0N2iQYC+n8ZgzG1mpZFq6zel7rZLMRP5hhLx76DcV1d9yr538LbMlyMGFcJRc3v+
SZsKrknomNxA0VyT/mO9dtD9iAQOV4bL03AVsNzJlR1TuKP/NcN3S0nrJn9jcO56
+WpwGxMlgftCnVCA+mPONzRZyvJuUh0jAoTXXQlO5DxUZeu79aO6WiJ0Wl5Jenn7
hV7kqwqf7mfNrUcThap4UtIMgWkmiu9moEkodp8kmlUfNdnHnGRe6EGXV3iWF00w
aHumBlgFcRtlYnEH0kO4AiW0I370l55i6joAELuGriLfJTUhY0T2tNxhtzYTDfyK
ZWg3Mhf4vFR7QDUs3JNtAgE+yKiAmfUQv+gsT1f5PQwrUyXbx5pcpUechoVNLf/l
oqPc66JOyf3YGjnCYuQUUwHXfvl8bcHYy1t37kKbO1mOv/97V6se7U1LyX71spsC
NpuvySd10T0QR0TsSx4Pm3pRRxp+dGfkFffhwvkE6j2jLFs50eBTpy23HNZtXCDx
rWkTyaC3ME+YQAYK7xFM9o+ahXN3D7WqBxxRmi1ySWrODGcU6cYSl3bQMpedR6Rw
ueUeDGVjCOWwvqk0oX4ln01gsZWPYst8hOFyOtgIADK8d8445M0Hzp3JOQsnghhB
WZ/NK+xNUqAT15xjcZKcU7dwfkolXSkZGFa877nO8FIWMmE83DS1AOrL+Uboi4v5
kHv0dSI0UmRdpy5AbK/Txx4xogPElCir4niRfCrWeULe3k+VpCi/Mud0q4F3FUO6
k3Jt0Dc1ELkCkm7UFVrAwR5Nq0UfjgxuTKZRrW6rU9mKPmL5NNW4blfTOsbCMxVL
ncfzbjpaJHPIOhDxEsQ/5WSKXi2vVCyexW0opiFVql6i3cqhIcuzoRWhVXJb2+if
WliQwHANtMSrZZO0J3APB05IMDSJ/Ij3TA9bvEsT1pSPVNn/suNllTqAW82Cb7La
38P3Av/1YHc7zfZ4Udo+rIB1r5uveKNeovSe4u6ZzrvbMd98XyBqKkom7wF6wUX8
iKGt+RiFAQhO+srSZ8etTVplOMnDkXjb7UblVj3KjpJgKg6K0NG8SjmvSR8a4f7w
cE1m/i7/R8H3Iw1IoCCU/ZkSGdhOVf13+1t7O8tqEBUf8jByuoUHHC4FQOLlz65W
i/SXOoyDQuKKTr26PhJNlfAriCGMz0YG5c4QjjjNRvxKuiYg1ta9aD/DfvRA1z3F
XNxrm5mge/n3HC1FvWvValE8U+8z/hZv+FM56BFTOZt/Uquk6Kzl4R+g2l3bQuZD
pANrgdXS62MmqR0fytOWeSdSVhPIZNAyZ6C6e9UFqlTrRdQsqMNUXo/UKJoghcxm
vJxc45E1mmZoZG1F7jAUMey6xcZ+d8cWY9Nx2OMUf72Xc8EQWGhO92UQGLj1YUJP
LDFodeRd3dEJWjHbre6XwK0KdugMNc42JTf7+kiGuLuCpEI5u9WrmHDaeJU2yvz6
2zdKPCR5PwdgQp2vZtY+DqyAfAwQtofKcZk4RFuEcUMjHzfw4CjD9YfTWtsK2GzZ
DkLohP+o6gAvCA4+GR/6ex+nzDGCZzxXdyFILtBPgCFQ8kA7NqeqPfO66r/gn3Tk
yTMHxTsKPxBjwkQaZl1kbma+izsMXyFrpLDbM1zIXosOH4HZNCAGBMVJtfNdgPEv
sjIIXMCbzsX67VN2E9XcyXc3fPrhDq4Suxj3yM2T9D9AfLi4Dg8OdWwf3C8zZu3R
dcdlS7RW1FNWmW3KUyB3+PaKf/RIqXEN3mBhHTmMOIvTx6cE65QJx29ZzpnmH9Dx
yzZWr8RYbJHySFaOzEKQNzLMzMbyZZgCLSTdRWdo+yvV3ET1UbXRhtotVbhnm2jX
Se1dxjlT7iORfjEOSVryzNa7dYgr+utoTRZdzV/9K+Ih6w7znSHlGRJ+yIWWse+A
b9lRP1lbtyjg26j9CfpqAWZ/FXcmL26969a1wJZjKgHW5fsxRubt1rqRiBHJeFqK
sZeWlLEEzuxWy+ZRmpx59RNE5+MdmDNcMDoNz/1nu1SrGu1cjyUVZHwQRT1ZjHed
A+mOdN8ZM/mOpLYkFe55KMOgeRNBGy/oPuFPKPqlP3Gnw4cf5JOLeh/hki+aGl+0
e0UhTwhg9GYQS7lUQMJyo4dSGgYc36CZYRQNO8bF0iV7hM6LDuKQVl05aM1LNNc/
JMg6WQIBZDhzlPawkrEFPBt5DEfldRaPM5uuuSApBeyrLVBTLzqdIIioC2im3TQY
9Qpnwkw3NDy4LaJlxGlpewio3sjbaPqKSKSYNZaAkxYmbI/ZWqBsw0mry7v2zOnE
kGPlqzuyft6gTcnSqs7ilW0hwGp83eG9ItlXs220Smykn8ZZQ723LmuQQjB5OOu6
znQmwB0LfZxiVolFGwYXLco5khAHeDmcs+nEVRI8r4G2b7zoiuFzQ9ZvQB2c9N3s
qb7W5ynC1BNZcEaVI2gA3IBLXlPfpk2P0U84CEmNuu9/S+73014trc4e1p/eZ/CP
PL923BWJlIZmkBQQGX8WeDzAOZUzZq6aANhA5NJHqX3YDzZt4vRQht+43twgiXrD
u+7wRga1bGNpPfCbRRiD2SaUpBy2aAeL0b3IK94ep/1w1E6txNKRKk4nlMfgfBMf
2ON6truu6Fj7ywfnrQY/92c3sccFp5MWM89pjWcqCVuaeUAgUUNO/hhODWwmpKgD
9hf6fydVQO9vuxN2rLxCsAE9UItY+ubyi8EWK3P+vzXQtPgqulaysMGf/5NawPp4
l/Nvwz5UDwTyAUAphkSGB++IVdwYsf0DGe/zSfGoWxcD5U/hmo71CT6TDyWTgiYQ
++Z7G7hkMmGrHY9jGImsCFqjj8eIGlyJufmVKYyhU81qW6tEBN+NkxmLfPj/RgYV
9WPjiF+xDNxExftFyicM+5Kc+2IgWJ7k+cvjk55iTFUryZRyOo1TG5bfSn0KRmwc
4TE87xHIgleP8MtvI+QKcwvCUttibPwKBBwSTSEbC53zRBTSdZTTDqxsb7kyQF/W
qnpMO3T3vmgDex5lj5J2fPxItduOyVFqOfcISJsGmhZq0nuXHVHPyVMVusjht+jY
i4quAzzdzzE4JeC3vH9yKlPX100VUog649j4ZhGvFlUIyz9ZMemQ3jGcQCYW4BYY
pQhkxIHZPNumypJ3lqdyFmXG/kibG/dMVF3itoY50BkYorZc+E4uwMPxc5MKXtCZ
gyvNnJOvgMiweJKo0qxHcigiWvGQBr0ct6o3yDLWTYDSaEqYMuijadsfs0+111Oq
MWeq6RxdXT55ityQ5P6WTgk+dgspLvXfBNgeRJATbsc6BRoxBG0Mfm0yldUxWifV
1VZm1YPYBV3MrtXAj/F5A+PgollhKjV+NuyUE8TSZqJJ/RDWvzdK8vfRZqlJMtsg
wWAJ/F74A8RDG4/GnltHYCBWGZAyop3+YKsmr6oXPcwrCJgRDOaq5rWVxIWDvq0y
D61WcYEyG7wPsT0sTjL7qmjYkLp5VoM8DxwZfgdp4SOjLOzLMwb29dY1uHhdfXMg
f0b6lxNlhMB+SXHFxb2uyuE0dv9VoYweQr2ESBP4OyE1+jDYh55/GlpPVk1862qH
tqRUsBchCLKdRqAVNoBiSOHVeyAa0naoKFp42H7lE0U6lnaVkv7NBloFrqxLKate
XeVJjbrddomafRnGMITqaU/cQ7EaqpOLUTKZz+7IkIkSMftDk274vKLfhhUxUfbG
jyjDY8LiW7rok1ClC4OH1d5/c6UypFBajHQHWYuWILeaJhokhk/0LHR89upvb9go
E2k6em4HCW28KQ9qtmHdc9h8pYXiTMHWO20gqCoD5BmqwxrWef/obYK1Pq+5khxl
aKJhPXnmQS83pbZGbrxrgafWjm33kv+yuq+OP3QMMN+9rYUoGVs0W3/Ua/b4Q9QE
e7w3y+se4nkI5LImLPrY6264sG48S441po4MmSprizROBlVV7l+sCOJqzKyWysop
oNyotuugv2Ix8Lcndxrs3aoJZn4++6myuZ/rrdze7IYwIsENg/QI9fEvcpJJxMca
WVWQ+BcK+YNhyoAbsIEZ0d2CJSuEMNfbzPhwqx70oqUFxW2VkQNklBZNM0yzD6XA
X/MJY4sEO8+4GfLKbWy6VHk24EojDlshSyZImP656za7uLcmObVvsAO3bLkn37ew
IdIDuWnCxBqkgDyGeEEYhof+XJ5DBSDMy6oi7PJlF3++u87lj6n1hR+jjR3C5Y9E
yF7dx7cO8GQCmvr/kqf7oFz/V/SIUpZqB0SRTWBH8b54Yc/zdUXYaM72Kg62z4Vt
x9Fw+cxNCsKyZdgANH735RwhsevwSslZNUr05By7G+/ZVFN2jnQHGw8BShHzSZh+
fOd+1B7RuklQ+9LZacCoNk7nZBfSG/T1+MJOA03A70xwLSSco5kgwpiyExtxqVGm
s7id0XkUti252cLyxOy8RVRbUtEdKsss+Tp3sT5zQz5Eat/GCBr18Jyi9oQewS7U
RaEUF2ZjwwgPkT+P4U/5hp1xp9nRYUI1i1pXVGNN+ArHEcm4WXWhRN0e+27K6ROm
tFkGC0a6j0Ne7SpWgKqo6/bup6MGPn7eNrF+VhAl7FTjP9LKrDECSgM3eGvuNsj2
DBRwy8OSQAvsFn+jY74QDP/R0An/XuW3aqtVROZHHe85tAPhDXH+5y2DzE79KBdI
M+Wj2n2nB3p7vu/GYsONAkLeaMI7BG6GvfzVKR889hhZ5DXOjOHyoymrCFvmgyGw
7mTPQxaghj4/CHB0YiRnJ/3nM+uockjqo90BoKXeuELhaEqWTk7dSAW14iYGMUAq
2Blin6z8blvAs+RmkmVtaOImXt2jYNL0S5stcon+jQ3JY/RLbRIAXgGJNoYL8qfR
M67fadGExebBrKNZpbfWfNFd6jpXd0pA1fSDDtTNufuXo9Gb8naOoISsYbZwhHVy
MWs5orBdPh6USDUUfbWkC/8QO1+DVt8oC889lzcmwvmhhOewHAtmJXIZJd83whhy
K3ADu88qgoLLaT1Rjk/r/cofvIWxB1a6X96RccYeaayWpmuPIvL5RrHl5/nz0XFW
ATn/dbnIfBMyjXq8JH1H0M38XU8MFNZ/6GMk4cyCRBfatdoSb1xD3wYLtL2Z/c8b
Ju/NlHVYmt9BKtHWVtVGCeOBg1grzW4gTD/hiYSpkzJZXJWx3FuNe5aTwVnFU+rC
SOwlnwjcPSW7D5sb3NUlVb0Coz0hv5UlWSA4TmElXH5jVRzXETAbgckSSiVdhAcr
zHDO986OiIO7EII7QWmTF+sP3vo+FCfTvm0xfoXg1w0ls+w2+1RgPkJAmJQqbmAL
1+CHaJQJga5QYeofjLLHeZgC5wYhbt0WslnrdiCSKAU/N3Gd0785cSs0y9sdIc0d
Tpck84iPOu25FMhFjhdojAst+FFB3d69t2EbESBQFMpcKcRkK6QGXQgWY6bxROT/
17y17TvozFNNPA6BSrp3RvBKG0A+p5z1Fs4VWpgKH3ahoAM6wJifvkfdLhdMnlGX
WMuT3ViRaROPh88AIQtZewFeNdp6Ym19JGGUGndBKHXgabhf+QpA1AVUAUEHz+Vp
6+MqaG7SJepqocUDQMv72rOb4hl+bc/V88/NLtCjLzD+17WR0+ct8K+eXrAKPlAl
89HVk3v6HsWxDRGsIe3EM5t2i5rAKcdME7OOKyPao30WJyt16kER4kI3H6sgWOrR
xa7ncAFUmj1E87AILl3curX1pAx6gtQsdbWPH5+AVbev663hJdHuOfnKEmhSbxVA
hcoBz8j1vdZtRvP1MOoJz+L39yqoEdjk0hzRB7Zc5bq2DDDaXZtCquK3dRRJMMV6
A/XMVJ4qOx5hCYNzjz6ShV9UWoxVm5aYw4wuOFyeqqWsNv6UHJL8dmLJoM09I0ga
o3ovZ0KaZBnsnhBYeixkUriHkWWXNcTV/qZuRrjpX3xA4zpWeXJVapsKQV040Pq3
JdjR29IiDIkUoHfOWMtMxObx3ILabZh2fvaAWfssqiw9fbtodRACwJCwLv9PBfd7
iTIHVWVqBx1i3Jq42ORTMvAtNyxOsNnSBssgm6I8tNrN5rubhI6N21S4YqE1vOFP
o86qiIkyyHZFlq9fEwtld/27MtN8M9mBumPewkeDVPgiAQ8w85MkjoRWWKQEMjIz
ELi9MShF7xjkkegL7sErBeMHLaBGBjrrhFelxHLsQXI7lBnTYl80NOccIMp9pYJT
XHBtIynJoH8F76M/Nz1rnzVi37t5HHVIHlaIgVFNIX0gagvqY2ITHt00mpb8YyZT
LdLaa1k1ETufklFWPGxOEdrfT406fA15j8g7U8B+/+3z7zNpfPvnGed+bqGl/v/x
q9TFWe0cH8mM8OIElBTn2nyVa2hyA/Xbz6oVLTfWlheZXaPcia4jNh/NrUB/R56o
HFgL9LFNrjeO1AX5zx9g+q/rYlDEba93YIuwukXzw+AO8qPCuPQzEdaFZF1JPyma
Vh2Noj8WW6Fv8vqkdQSuD3TvKcZVG2cTuPbsxPA6f1IYViOshdQrgO+sLcFS04Y/
iowK08pOZyJljwgIjDy0mCH8O4izbAESJhNy6tM++BZcggTr54bCDPEzvdtz//EG
+7CpY1jdU8gpeYnitSuZu6E/BtzTaZtQKsXN58b2hNU8amrHKT4XADj4Ani2dQCI
eKFnfOKa2UhL8IMKdEFodGrY5GSpY2fjQTqoG1UubM6n4EwKdw40euYfGHFg6Ybl
meVk6+RS/f6QCqel6oaLOklXg715IyTv6N2qqfAky6i8tOFdlZJuZJN+J668PqJR
/r2yNzhqwU4m+I+TcXUW594uoN7o18WtQNsbhh5PciwMn6RRYxpfHCdC7y+iB8eY
m54PUuhp/V3g3rPZtjryNEDnxAiFsOK6UhtEjEBSxKJFf69WimpNirneW05aMmGh
KxR0/TEzsoHRHzGC1jK6jYrbwIoLv0F7o7ymVRRnPEF1xQmEU0P7bdif0uVBW6SE
yowSC+8tnqNH2tzAfd1Soq0jr+JKhmHOwfaDzXH73FPw7ETNqsFAHjUwhU+dWvCg
C2JnWh7L3W9wQanowNRfOuxXvGv0kpeWAWmTKRb0zRiz2ikwF2+LUdgHbhIqhRhr
mIXmvgOpMDhYAQ79cweD5Sy58AZ1f2hovL8UGebfKvPa62jPbkFd+FTZttvbjCSj
r4kdfXeZjupTLeStbOcIlRWxbq32DWrwvtGmZt7FsrXr4ThjgamrWsr0Hqgs4Xnv
HIfu0PArPUJkfROJ8Q76fJxKIbY1SxqSXnRaPjTSCftHBJxPFzBmVZd283iDfwq8
ZdW6Bzd+myz8KX7l28UsdveQBibN6O2t28KZSteEA4AQys8gkPpvLdG8sSvmDDth
8++SpH0b4ySnI/QNktAWgQgSKoVDQBEdeYqTpW0fQ3+7iVIdRnR3dFi1d1cXnS6P
gFvM2NXYfWAdwKooeyvbQWdSKgTX704Btjt1V5fKTO4VLk66h46kwLcte6q0ZuoP
W2TiXRw1BhatZ2G4F3yg97MhUmQ0tSHLYbjDWICq7dp+Ysf/tRnrufT1jFcv498p
E2MWBaR9KFGp8sj4Z7gBQzxTEINV3+M55F55vFp8lhTSTHXlRP3AVDyNO8ZHaNEN
tf9syrXNrT2noTMaT5RUjchHamzjSTeSpumXJ0qIcpaUkP1fOpoep0pYX7JEPcor
lKdSecDhtbt3ydR5K3o3EcCNEkSOzEfgZamFePx5noM6Dh+Vz2PRYQPfQnDNw2uW
uTWnHvKzLgqQI0ULlayC0lXDIapelEnFcFMHzfykFZZSGzjqBIUc1B5GZ0WsU7O+
//lQu6zpHYhRf8h7wB8pmkrQZ4meCGfcRiP355/NFLqUnWlOAq8L64bRDcHU/0Pw
dcrPPAcKVm1zlpdnGPBAnhT74sGcjAugNjKZa15lMRXu6v0UwTMPa6HNRP87ESGG
ieA3QpXpqgv9ytf9lMv7an8LrWgYy9Pxh0Z7tdKF8sTAck6K5KAGrmHL0uc1ypIV
kLpmXJQU4crYytk69rRRGVygXizkdPD0deDjm/UAfobAS1XWzpXWrmKsCaFGwk7i
JakW78wjblXOvdcxPFVrPdtZx4XS1T+imSxgb+2gSiRQaU5cNqWBvVAk/PQSaMIf
5U3/udwTywV+7a7rta1idlt4qmrwRqXgZ4ZzZlSvJnoJ7kI/dI38nMV+yJkj11RO
jGejGUl8SU+EM7pQIpk+rK3+/Nm7wz5uu7IPsd5Y8CI5ZR2w2l7VRA4VQOzqO4d+
CAJb7EM/0FPdoas8FlMpUUm2NRrCA8Zti6o4fpNf6NZgA87eCNW7+2dShl3SoUuY
GZaEMUF6HckBEclIFdzGelasuGgJh72OA0um0KK4fyWTAgWnNVLVKGxC4oHgKS7o
lvRaPaSXXarjT7qnbn0vGBYbyCTm5213u9cd02qd/qovq3w1Qs1ejKy0V3o1cabe
8Yp9TQYCdIIZi9P5Ka3pwxKrTjLUuUG7iue+4IFOaCXtj+k5D/f+X/6Pmee5XUBA
kodGjeTlNtP0rLZG1aZlhtT6FDIhC+S7SBstZZV5/FZ7YwU0zYu0SKBs1+Pzbq44
9vCThaRBzyaLP5ToBK/aSAxbpz7BSQdCBvM8SEE90nMFR6Ql0ncSSVJANS+QEk2S
WNt4UybSSuaimzJDicQMg/qWJ9I0rLEUVMEKzuLPfBB0MA/cksTNxhleiBjQBmxF
j0bWDAkGC9OHWtgP2y+t2ghrNC1YP21aV8x2BndQXkm0AykcqpDi/GgFzQwyKQSY
32MJFFjQyjs8Yvpcs5DE+l20TYF8StmAeTknScwco6TbmQb2MJ9Tcp36Qj0PZx0y
R7WXHY8S0lOpnfmS6HzOpJOaovW6hT1gVgK3qmxytxnI85afpksizHhwCiZf4pvD
NwXM1+A5rCGtzdEjvNlLQcr6eP2C8+cy1GFq0wApvjZy8qfAg30Zem9BCyeDqvS7
tJvoB78bOx4jgGpeSXZWnKH15o/7cKpDA2JSy4CUBoJfmVbqPC+i8dr78NKko1h4
TKCADfLlc74iYA0S2Vo2BW7HbL+gOPiyhWmbdNd/mqGHfqqmi38uiMf97OB6yI1s
E5J75eLkT1XIapStr6dHwOxB4EStvzhRpyOKBguO9J0gXsIS/bjrDiqcp+iBCOUN
H9a6FrK2l1U8nlfjttbpbCw7lPvj7yUPBcmjzrbIwZUildVtW8hjTBIh5cd80heT
56iCDMe50VbFANj0d/C7ewwjfKUj+ccVjSXp+/G2744SBFjL+lWgtdpkwTUp8IRi
siRLYgzvTnAcm+6ZZ3cSsRrfyBOag1THUstYHj1LXhzctrffJvStdiPvZFA40YaZ
7jgsk3KDaMjfO3KNUlPQUM71uZ7qzgSJxvKnchpIZiQnkHx980dGfVDcmEHCULDO
nVXwZgFHRAa1au+kEgQUJukmcCk0B8vgAszo6pF7QKh0Bt7J3L9ruebxpcVCD9pn
xpRpCsiJ2hcR8fYZGYIk/f0iJgms6B/CBn4OYQ9fW66DPJASR6r737jWiKYvhuDe
37HjflPHc9FLJFfU2TfpaN9bV4JWzifc16wT+VPxq6CBr7WYAjf1l3r3WxdeaPF0
gJboyEfsQKGfgJEcVIsZRuQ2JurSG4s9YA3qjCkKVH/B2o+Ng/WL9mobdsg5LAR/
I0IoinMcORDU9w9eZtTW29/CX/6F4WxryqFxJsxOkuPz/KEEXD/Th/nQ2Eqh9CBJ
fGluSZwF+uZIxtdfJ5ehUSJK46bUOVI76mDu/9twnJMiNQweSaCgZUneVoJBfJP7
01vmjYFQqMDy/msBtXFc9UmJ1F7CgJ+T33FydpKkuEXWVdLzyMC0n2y4E3bC7U8E
5z2swwoaHcm35TrrOIze2UaXH0Iqt6ffnI8R4PNzvC/MtPw9VDYPDZwfbZi17o3e
gaGikayeftRC1atM+mL5ja2FDNm56XpJgNksQq75xGoFLWfEbS1O/xm3wWzb75gy
q6pxSBiIfs3JWSClhPTUvCoIftTBXFEjvtieODIaZZSz7Gb3FMNi/+KrZrrKbviZ
JRK6ndwq/0/0WG2U1tXP3Kz59UGIyRT5hlLRRazBIFxysR7/eqS4PDF7IFZqwqps
PCYBoZ6rg1OvTEdlK3enHqu09LxT1Wks4P3E1De3nccV5cztRwNt3QPy63s31Ksb
EBBPjT8w/LSqbYEylmR0WHoXw4oTAJQlgL2pAtm06sDz3nqnxkl/w1N90IpKhSp4
rnMtA4fAI5YHjkjSrF3oM/Dnivu+39VWT2sDryVye/5OsNXIIFdJtz1xdrrKS3l4
+8YnB3LGYdYwIP9UNlYJRjQA54lFvXEfgpFVfRdhMGXnKkVY9ZBSC5QpHoawdl7u
eQZW8T9NZxM5s6nptItOx87idSQsUyMSwLP6cfIpx7zzhmxh4dDFmKup7MbYELfD
4fhzYt6HQM7N5TsekQpeUbDEtSaoNgwJeRE1k/TGvF+segHivdvUbLwDnAkXVB6c
L9MVrer0wpKcvOq4SjqhYxKy0YtyWsRLegORqF0kqci/ODKIVGYfIBBnecZ0v62D
H+Na9f1zJPIIqHczQzSvyWuD+96HRUScGnXMxDBhabKAjgOkm9bdtWlnEAEzAu4/
A+d3tT2dhjXyKUHazx9ZfvKmbGAi9XTg2aVRAc0q+WsRRXoErvWIHym7eRmVo1Wc
PB6BbsxzCm0Q0QZ2FoW5/mePzNWq18/EqdOHc/OcIJMvhvFEnFoE3d0z9ItDDArq
5H/1zDuoO7IkLvAcuUvlW30Ocsmm5A+eXsng9RcOFquXj/BWmHH+uSZAivQES3Gt
hM6hC589ym0LJFLn+VF8+Fwq1SRFeSoviOMBPGyk+E/gdHi+0il/+CoXLPgIAdjq
OYwXTr6xqiZg3Zp3xhEN3qv1QyMQIfFsghNnrJM4GgcgfHprSJMGpugxs+di1cEQ
rXfQh5/HXcFd+oSmAsa81mCAYYaccu7GYm/lFeyv5+FE/judj7J5e0Y3fA+DiF6c
t6A5+L4fEfo+4e6Q6/cZh22hVNAK5THh0aCn4sJHM9G8h9W/494mBOylcTnNj//c
a5D4Bw0iPbLL6R4fdzEH9C2r/0JqpnDcOtdFhrlR05ceVlNrZrEfrh4OCZ6NwQg5
3rHXUlqex5N02gmuJUiv6a8JWFVsQDW52pO5Vo3ocvbRz13+OPufvosPxUPQF8M4
lyqzrqwwUEG96mjC5tnU9DZ1FCRyzq07UBMGL7KOYrjZ8QjGVwBBhvk9sVp0RNNf
1jLLT5UCOpVQvOBYgm+1o2DIcTvW5tWtJw8NoJgNJfId1aXJsM3n0gE6XtVk/Vkh
xysLAcdjpYd/vBffwlBA78vyx9tLWmN5pP26pHHj4EmqVUGz4kU+mDGhxYTBYY2J
PjfYvY9IPxdytROJt3SkgQM66zTC3sTXNCLTMQzKNrD0S+pte2E5EBsOLDf1ra+M
zNtnThVfO9V7oBy1Hq5pWvCOmYczarvela1hTprgMP0h0hzzrM/3jMsDyftkW2Ld
wWSx+qnfZ/oLNpuXeFHHd8D6NScL5nIq4qKdLbTHMHZD4xm5LG6BbkurD7girAsm
+NSh5hzDo1hN0aAo8ingTyFa6/uyiE2a2TjQ1Y0gSfZAEvLmVlxK3RYrjYAorUku
vjtjQAMT4RGURHRM2zHiR5Io/1ibPRxEa3NbI8qrNERMceoNY4J+Gjz2TfzgnN2v
89vaBy2VLL/sIjHW2j0nXFqZ4lBdXc+TwndB5NPlQI5ud0xKQ2q9Ga5iOIpU1qKK
oH+VdKzzLXoX5Kkfg44qXZRnEg+NsFe76OvQgwd+VpUj1auV7DWhNZ3UvYEPjk4C
OC6EjkoQGEkmSa4fgXEMRei0DsF93Cj2d1pb9hJKqGDR2wheHUEFHewPfRdhQdFx
edrWVnA9oBWug/G/aZ7h7xMdIkhyBD73b5a0ZraMKEOtn6xyRJsbwr5ux3uOhROt
SfeHs0IBygsgwjGRJ6eiLr7ZCYmP1pgI0Hvx4stjT3KbFPc0QHNHJwNGGJdVJ/rp
9bHeHCpRqkIScU6bBikRHOgtUa7LCoa4rtKGJodjjAThQzO1LM3tctbuQOt1X2ic
XVAsK528j8W5punqfKGbC/eVvnnLMaAdOoUVdXxLMDMGDpCTGJj1gXiCFdS4mG8q
1vYTFdOsXGgcLuyECSrA3Y5+1sLe55eSk9e9EgJ6a6JOQqcqos7kr53l+uu8OPak
1nLuqC4ybGmmyO0Qx7iiilCwhQJU0HZi6PELbALOV8SCoLkAJSw75RxkmYSWbmdo
SMIQcpEomH7g8uT1hXyOHGj+g4D6E/nNqIpA3nifO2AR3rmFKZ37l8RBLUmWhav9
rY2vhc/NmuOwwsVH2VwB/9nAG0+W4rHiKz3rMTCdIwPse/p1v8du6C1/2257GW/K
9JIQ4B6w0JR/jsfVJcC3Ozn+kcOQKcSHwtPkwcK5gq/wuHYe+AWroTuKFXftZ1vh
qkcD2HpGyC4OpkVqU27cz6gRI//I/bb05WEodfN8a1ae45ely8TlYI9doIvvNpKt
a5QcvbnDDHpWT4x+zR4sF83jRb0bGqwOlmOyJgQLwjszCKpk1PNcvQB7DuRrbC8f
z7+ETxnp968Snh/qZk4yG4idxxoTHGA8HJF+mAb2SLebDJ768k6IuAteuYgsyLDg
Kk1vmvwW3txZSOIG4Cdn6WdGLXdqhQzVXCnKlQbshESSvYFozS8GvGmsgmXAkw4p
CT6tL4tCITHMb8f6yj7JUSeN0dLHNthCCSJ4HPicIh9a31S7RHkuhK/atvE6kRHI
pORL6+Jmy2lHIFJKaP8jnHW231salhix/gXu7I1jPw1tAvQZHk/SYYOIZlGZPuqY
qTtzlcjkQJObsZSm0BTxZJMLlUaLwC+kawGTf9N/7qxus0LeyeQqNDRrnOqmwct9
pP7umYtJA8mS6N4y3tAXduK3PskfyCKLTJMWKmpjLm4J+FrmCsYkh+uwOLmHQXnp
O5ByptsHdgED4LMg+EhwcM2fohQPEu4fbxlfxo30YtIxbDkmFRYZhufo0QFXnt5S
PzVrWgi8MgTZ4DAeF+zCu74qSHqI1A0RNq66tzz9gCX7ifzhXud7l+6b8gzPELKY
gn9eGf+kurRm3DaSEExeEXrzCv7CvtsJQg/ca4tWxu4LV+2lyfkjlq1gciq3m+Qi
6S8b5BjmIOzNjnic7noRzUlCpIhFasXUX/rJ0qCnOLszffqHRyOdO4nCWDUWeO/V
3+Yfmi93pry89c3smNxhPoR2Jv4pF2DgJKVFXkdEgZllV+UZgKJiv89+qWrHjjvO
q+thGkT3aczcAhprlkVie/OzqI+Wx4e41YiJMkKGiiNJbEtz+nychLiJKdGyIYJv
IVG1H/2KiJgcvU8I7uLoD/NhUxuuQ0l40tcJ9GjA4Iqxf/0Fb3JYrfyTlzWEjl8r
PS2Erk6SR+vF6PELabNX99YWFjDrYl+mJNaEU5rETHUcTaDaQbwKfA0kJ9aKXQdE
83oni4T6Hp8OQ04Pq7rVi+GEr74dqVdPe3yokaCheLy311fUFKwYjT7YR6DGB/fE
l6lFI+SOOwEH8SOHS0jKtvkpIc+S6kbjL5IusxIq5A/sDtMWIvcbjUb+i79H9aar
0VnAzKskIsUOF0Vx+eeSb8o1PZXpJ4qvksdiohI90/fGKWjyYM6HFUpRpqVoNziZ
YEKv9nZZD/n4p0469BK9GSbsl2LulHaO1LGrGJVQARz5TrLF1CfgKYEO6uL9qfZj
7S48JpzVTLu/zlUco1k4gWNLGE+1ESsJ3XSByp8/NZbqYLiMTS7VG05tncTMJXTx
wFzPdIlInNvW7pZ+wyN6pp/zd/IpmeB9uOoH61Mab8oHJN+zf9QOD4L2DybJ2KQf
LrXXBDd1SST9YcT7VUNOPCGUFeJSaQsjjZqhT6kzFsDD3x/fkJmIUvg7DJZZjU45
Htfbr3AQkroCqG9u+0BBv4gsHqCHGby0QcFEmS9yeX5nZmoJ2A0dHOmL0GweVxup
mmZk3gCqWsdC4rJE7y1B/oOTu3B14eKXFMqwr56eEJKGSpMJcnGxSXnOpY2kaBWU
R3FdItyneCFDZDnl2YanyrrGCPFPQ+eGIx7wYTnXIVVYfvqQrOB6V8PvZZBzGVLt
GolNdGNKgS4L28/l/nQn74OHlotDDi7Jq3ACt0B9oODeAUI9LGhkBodFt+pN8hIb
b6ZaXfBZVVEzigcaKfufo9PVE5HA7XNbHXkhdhjyD3SVM+KM5CNdHza/DKrlu5Sv
xKWz6dRYQai2KgCWCUe3Ed7r9PP6j+slZZ1XdNQhNIXH0H7hMYrznkUhWf/P8u6/
W2MF3Tn+ql/JZBqUE90hslLI+ux9q9ZZZE9NwqL4qPQwBpO4Z+HsNG1iy54DUT+E
j+WzE02XOhIxPwADICka+nvPelVbpvuTp59be1ckczVki/czJeEdpz+3N9LGSCHc
Hd7dOM6QCwRT05Js7G3DyeLjr0mDHZf0fI0zU0pIzAbbEP2OClfkqULHTEnZdWui
VwLFrnBHBYLN74Fmsrxm6+E2+fQwvv/quH/nGMtnMFXTdqZle8OyTWT2yX4Bqk7t
Yr6oyhNdrXJ4cs9at1nBFfodPXvee6jLxr6iFT8+JqlLbDLyhpLmVVsIvu3NtIel
Q1sjjoiibybAwODy2hqiOB0JUHi2qTB8Cq2V15DZtXOqK3JvYWGIqYIH1RkP3l8Q
n6EMfJ+7t3ETNxBFHpoFxUyxw39rhAj8FsHDjWuIqDCTOOEbOq7Y4D6koX7Ravzo
lyJBYqUbvpew95yd6Yi30vT8qthmu2L0Oslz5WKk4nwcdjEL7qecVo9ouuUxc0Js
lRMBEl6SHccfiyjQNvNlec0bBq7HQvzqufjo/4s1j/7yk1XPBrpjbRyVCHYxbnfI
0w4gd+Bt5UeuTtUhGziQeV4N15TGSIMHpoZHjb1i4S/OvylrT8z8W0f4eQcUU5ng
Zgt93opgkkf7r8sStzS6bFKZHdCy6Om7EDFj3+PHcw1rYUe5bdjXF3mIoslO2njO
vHrsc8rA4wjpxshMAA2Dji0w3XLK3UYMu73wUBKmyejaCSjzg02xze43pVuvcEnH
6ZHyutlzaAAI7D0HfyrU16nW9Jmar8YanMiu8SNGJqCK1xIE6/GKcjIz7Xyvuj3N
Z9DrIPSfJuK2ACkEcvXtWiAuM+VVoAqS9eQkc6sQXy7ej8Ni2KFMzOtg6G0ovSIs
4Ptkw06JtCMUj0j85T2YzwkQeVH4R7YEZt8T6/cEP/WcUvoe80Zh71QH2wSBLjot
T0dK8iUOngaPvzMiYHqXZx8rw7vfnQ94qVIPXlcyBm6khUAm1gcfGd8/74hvzOuv
qebJ4DujiHeP/ygcCVrmoEiUVKTSiAny+sZUGddxP+k6l4IYzw1f1+LTgIVsFheu
owqJzNVWcPrnFAH6ZJoOS69j4zohyBfjZiJo86GwNjWWrLcJslFDhMHae4TiaDZ/
OS0k1QS0PmuwbllzfW4Kh3dsJ7lcxOBIu8xsyEf8s84gAZfHXU7WDE4e4/gUCH/h
ebjCSdHNsn0HcYY+cUf4m2WfurEttKsq4oILPi+7oSJ4qg2VGOgKpnfWRuI4AWRy
Z2z8RD1dgjaQ9+f6SjEiYoo99/tESJZOBSFDxtNvsatDEx5lWClEsN4M1XZtrtlY
OYPHdNDVR2HMi2j4r1JTxh2aPiERgsee7A4YY9E1pKDMq23qcwbz0cD95QVSsluc
EUZ0lpGg+3/FgjXAypWuDUJsGvG9LnoT+oOOcKcodDAVkY9VQ9bHNBRNymRW8sA3
fMVcsxEQnfvGEDrw+CP9oXg8rA08kgXxe7IJz5E0rav8BXvaFUu6KesefToEIUY9
Pr5gDU3xwBF4Zw2vqANiW0+SPg+a1IKoptwNqA8NvPQJxQxrYqurfmLjVD8+0Mcv
B5wmRdOPSBEfwlVrldVb2HStwZ0XyfvIpkKBhxN5/Ed9Mol/pptL0/7JZ5TRvugP
L44XlZihcGfhMk1n39xRB9YULsiI6RAXrBmTkMALOtK/JtENpZMy+H9zApaQiVpK
hvGc8pfH0nY0ITDNID5I3rB7cW5lzuPtPZtSx/Gb5zRn4ipkSsVre71/jqIDgdUe
yZ8+DFd66G7wUD3U+dxNWdSH2wYWnzgEjQY83kWi6+YqmVoBpi5DFYGPOkn85JvQ
G6kC0faFUsjkKPTx9eCjvwDndT2OVhOLaacmixfLR1hkiXZVxKH3DBrQInVG5O/P
opf05PUVICeW3bunK6S2wohWVwvf/WHMbUj/QMf/3a5U6dCQNNAZ6zrh07cxCxxt
4P85NlB6vJBuyMovdCzf8i663Kd2DKtJiTeV+jG4uGv7NVwDzLG7hikBCVibYl1V
RQRQHRUhf+a3bBDMsXUnc3pJRtdqO14qGzdSK7SBqJqlplQuNidrlMsAngcjWVoy
9jUh9QaQ1GTwS0OxdxblUkAEelk8na3E+EzRBlxRkOu6WuIDmXukp46E7lIw+ktY
g1cyoa7e0Q+DNKCUPsUdXKWwBdVbYjNZmsX82OH5d8GiPIexs63V8bE3cMU3HV4Z
ppw/XnH/1uD8Kj8RgvE4Vk7tYJKA1R0n7T9Z5CLeZQCa4mAap7dRX+zKdutycPXu
4gcPzWbkGyjOj/JSndtx31RLBPfD0q5IM2frQNTAlFZnRCQl5zlP7gFkkS5GtBSw
wQr70DakuCb+JtwzlZ1j3RH79nLd989ajVJNdFMcb3v7iPWloXTWjxBxqiPmVr1k
/6NlFiThUtCsSo32qTYVSQycuNVvF093MRxb6LBAwiGwqNiy979Gp0flhKUTjiHT
YAXHuYyiFvT+ogszUaP/L+IApGEmZG6Cldh04Iqk1A0dG+S9pWlpcsxeQPLgmGHA
0iPnULiOrTlgMd6oYvHPY4bKbn0KpTbjgNhc6tnpKrewI7Bn905Zx6e2/dz0tQVo
7xPpRdcaEb+vm3B+8z6L4y91ZEEc+SB3rOj5o1nJ6t10NRTXZGghRE8LE+rK+4Lx
FpVxmvTmt4PEZU3DtusWkWyTmxDyVSjWXYorHG+l/C2agAvJAmyEYLuFX8Fw05Ja
09v0/mk2KZXRd8OzcYcZAIQDrnEHKxaumKlpzTXP82dA/r1cM14veU3w5HI5qNw6
NxL+r0Gmcwo6R9SP5pkmeiNq2esxzqHK9dAx/C8SUr9J6Af9U1lhzQgiTLTwVh6h
AfZ2mwMvAo9LyXPg2+L4YMsd2+UjNQDmjo2rw5Bk14B33MWE+GXtig+sTyNQa3aB
t0IIYEydqgNq7CpGsHMdqtuNLlVI/N6GuC9KJ5v0ppTwEix4u8aDW560Ofm5Xd1e
8qiM/bpe3u7Bfgzt0UYz1M9DNiYc0XvKhELRCLW7pclps1KBdpGymWM/RXfFmAQp
mqkyIgiJqvDB8x2rUo1p/0ezBkTdgj+GBAvbsX6qlbXJ03cS1VPJ33wisouPQTeC
PDPW6MsGTk86NTKdxynudYhgmfLRUZEunoYUWLXDjzunRct+DVrZdqDKUyh/HtN4
ThUGRM7wXliDTU4YOjlpIdHYEDSlEoxP3M4/VW0FbLMXvyhRK7ronvuOM34NFQTE
B53zm1xGzL5xWgDsIW2yoXaKZ+n+rK3EDdCFI5TukeYX75+97kA6vaP9qG/RPEz3
vnamJwhb8KGrBsLcdVgoYZKoQcLuVJLKpZk6xWmjOMTZ2xJ0x+tied6/SRgFrFjH
EVPZ3B/SrQbxDSgHswW/8LDA4G2gYcs7VX22rw3gzB+H6DIS0EHAftwfhp8eAW95
rLZAash9UA+aLvXKG3ihJhSn+I6fT2XeJUKVBFmt/d33IhBlQh0jL/J/mIwpoH3N
7zpeuu1JuVrv/mFd2tw5oAlWL18U2tD8uK4n9CJtUStIuEk+2VIf+fUcVXpQ0xNl
xDVXWxk9iWZN+vx25fx3PJ0qTualk42/7v3iVKjlzLYJzWm65GMgf/4yRh1gOjIi
nxSpKLQMbuuIgMivNR3stBulTso4DP6snFSyQpoQ3i2gl6HVUmPikVwXxu//ZBdo
liK8UqLYfNz5GXqrIhoIC6S6h9bG42tslZBrqhp2wbMD7EQBuGAi06lB3/v0oFJE
D5SWNDFkUFEWqOq/LAML999rBRp1iDz0vaNOI/PnlAcEPF2yMIuWIWcuHcsaDqVN
J4nSXUr7N/qly2BmAsDM2APVnG4okqjNhLNHhKOwVrlMFLWCK7BJ5nokHg8ZA3DK
K8MeYjyKgzFPlWHz0Y0FG9HVQz65hxcIOrFu0HKsBTUVdvigx2YEgTaWn+pmdXyG
/es7kKrbo7JFH8Cd7wNKKsTW2tv8hFkFGvTdVFRLAHiy82b1u/MRb7aokHrV4zqE
66SIO3/GfF4flTtvbPHDZDHpkj1fxWcnNa40l3o6XTMFdpXdvB7UD9ZX0ZknPYC2
+WAWi6uGaKjngMoMi+2zxyu2PCXAmdgFbvjlDN6o7la/aHGbHgC+bX59lD2c+x+N
FV85UA6NZNU4UE2bKNIeBiZDuxW0Q72ryW8r6rYm3xqeZBMMlAdBskO16FhlqHJi
bp3QJcpq33P71DZ3n9/8LpofBBn8Tr26kUlWhNHrt2sZaKtwDYZOMcaOnDgnj9aN
4sV4FfWVw+THMuAH7iPJvgQwCnyT6ZzyLL+YKthZhMYO8D6VhVhiI4SlCGFY18Yx
38hE/1r5go62k6jnvNdjZuJSFmFxP3ynP43EeQ+uPak+HABztURez0fE7aYCLOMQ
k8UUjmzc0oKXuhnMf8dKy7+EX6wEHf3ov4Tc9uCPX8vaXwgFjIi2eHdRC/OXl5w0
bLIVH1X5iEvOJDTkQdrDwmmkgqRFGgJuFdFr3ffSunGb8VfM8z8bb6ztSCfbKXKU
4OtlXW8Zkn+CQtFAbbWe7iKyMjVHEH3Xv0njFU5JX99tJQBv4BRLHGMGLH1Hq33/
3J7iVT/sV6fNNkIDSyJiwOeq2GLfwJ2MV6HTMBuR+6BNiwFmaZ4yCILodtR1OTqZ
dNY1R9vuvg77k99Lk9a8Akj3CE49WKCB+uS++3HhX1pyOnfTa5sbrEcGmvIaRyps
i7nNSagGdTem57VHz2U/W6Na0SlKKOyG1PE2MqvifejZrk6bkjxbzo/YP8OJCLgJ
c+xca6Wx9ApJUIcU/Cwzwvy5fGVDrwlptYTrPtNXKoBCY+6W13Ee1mVcgYXIxYME
B8EAQMiYaQEDhLleiR8QtZMLPtsze9Ykt687r9IhW+Wtmik2VQsoLa05+8XiuPFl
ESdm8Hngo2ZwfOQB9hoyIAxRqjD22RxvgGcROntXAYYg+GW3uV16iYnbAkOFV1WM
K6L3Td/gr43j19X/lp0fUAzlyZfySDfWCy6U2dXxvgM2sVseyTUQlR90n2YekDDH
yusG6Dl9AIbyLjgTVaElAbLbYjmsI1H6fWPS57XpyWi+HGR8eL3tb1v3Om+e1K9r
dMeqEn7m7709Gf3OF5GBapBFKyMXiCkET7vEdYAaaD5Txv/uNh5quSfQWHgLRoFa
xLSAnTXxX55ZplFcjLWf0yWU/Jm4XLMmTSANjue3N3M9qamsOlfj07Oe6I4lgsMY
eEp/Em7YBlz0rgIh0HI5o6ECFcl0fapCc4IP8Qauy9HWwoJbaJo6WTD0AwcO7X0U
0P/apFbpIkhD2TBE15tHsrCqiSuK/XtutSRL5A4QryrS6FDXClqbFqlP2wpHx983
d1k6qZqZo8efaNcOFrBECxfyGDvV5q+mt9hfWMRgrWoNyGmcLkjYsvVFAr8WLiA+
KfnppY/30AyAEGoXv+Kg93r+GBADXMLxyiuZBeXCci6XCrKl8cewyaL/DcFN6kyx
911sI6n46nlbAJg3wVx3mnViWMrpMrLlip+Bd0IVphJ+l9txKVP9j4bgJbB6A846
gsxbadb93iu7fbRFw1f4GxWphXfeRyFF26BZ02q0rexQMPIVyXK9v49Rap9/wgmf
QsvejRv0EuFahH909aNP5EfwYitRXcyPxXZDM8RW7nC1hjWDJ2j6B+wmIeqZ614h
XI+6YiG8BD526E7UQSquD99kbJC9tSEljfaP9CgPa8BO0CUcbS5f0gwtrnO+mnzG
jAzNZPlXc6aing1T8JpD6OuIi4VBCoHftQv+m9hKxh1ez2RFca2V4nqjBtshCX5r
vstn9Av70MuYfoL+JdoSlZ2NQGEhF5WAwRsPg/vjUd7svQVMtTqXUVa6Ab/rvBNj
XyaBrwKGO2lQ+Fl31sGoKiqFx1GIj5I2sLo2EIygWqEQDqRupJS1pEZE/CU8DHY7
3SkHyoydpCEa/aF0IKB3yPXIYsLwrTL2etvaIDhNJKwUE11BvjeBLnzfcGeHXWR7
aFSqf5fE1K/61xiVpjJ/wIy2FXn4crB94KZ+ZAtaSADJdEnuky5msVG2KP5DDJ8U
rwI1mSQP+jLDp1G8jkleMMsmsuDatY5CwvwOVQYr3wditu0U6TOOqjIuNT10Iqf4
z+na9DXHRq9IeVWQCOhR2It4sFrqWtF0fu/sgcilxwmsVaIa6CstrNe1SBaMsapu
PZ5//TaK8oMXjTf100N1oedqaB8e2JLMFTD1kdRUtncvgMDsFD0+/du9ASAy2FKx
O3NaSlyizniFnYr5iWGma1VaGFPsPhxpG7BIsY3u9WUjaYcD078phDzWT9WIZldR
1d6G1PuxPLWdamiUVzCKQeeqcHkUwblPT6SI5jxLR6TNeTsxJ3nldo2mwntllicU
vIqLq94E4qSonILILoLxYLa2WGiYFHFrDF8gyTV88kIKGmyI8STtZ5U3Fa+RfxRK
XLBecifJVKetZvtDHbJ+nE4jVnudhJmSJwjJuYmu0cOonsmZY6wfi5FR4hkeql7/
KhdoQ67PqTwp8xntdQN0YXXmbIdzHyMqloEij0qTTMSK+8bwQ7jY3EowikTNplXr
210T+DgN5RU6zZer5JQGrFhJPmeuMLKiFCvu2Rn8MfaV6+Ok9spTW6enHktgLFZJ
Jk4NVfwNCjY404PdjDrGnq4GQLAQv0ovQ6zQ9nlioq8L08MnjF8BtkoRBYuBoG01
YpVCQOoJfqotx6IoqFFlT1GQKcmKP64kR/72CkIK7CHd5HMdLb9U2hB8lU70KhCR
7Cs8gx/tQFgCrk9rrGmAliz1mEuyy7dI5Z69fj5KuzgSNv25llu0T/wePpJEMeWW
LXef4NvO2xC8MX1K8xfJbZ/hxOFpB47KtF4wJ/6cpX7o6TKSjQT+TsBxQeQfp/ZT
E7tqbT5xPJzBxHIQZYQZ6jZBIv8FpjuvUFgPk7LQ2rJsWgZHibhEdknotuir2mTw
9vlBBJFxqx147X01Q6lPL0W8X8U3C8gVgZqoyDKzVTJ4hXlbfDRfMcE0v+iw72Fw
2yOM8gIhygst8Y1LaQlUTiyWoP7fcy2DOwtpvaEFqN2OtapqiLFt+dNUKlpuYRTK
iC1m4Hw99ZCkjYkHj7bt2vOQrYnsQjGZQvc8+1tIOvdP5XjXaBPMA3kVzAfjgvc/
PPbIxqU/zArepzMYaNPUWkwN++zKbm2gtVJGmlMyFQ1Iorn12g6CE1uSgXKNiiyJ
6Q3rg4IRW1DplrNNRdWrvg+N2z4QJBatAcuDxhL68KbeuiWG0jBDT2jLLkICgLuX
gTImPTUDy5GKr4nIDrlwj1vZnRjj6evhsefBMdcian9ILr6zrA49+SnNnfuAtMNa
azLzUvRfD1CeJw5mTielkRMgghDLGc/MYkXk3HReJIk8t7w7WowCff7JT0YWmyea
Ont9m/TtZdftRrwiI0Pc0+jT8rC94Fp4i2+xloRIBXZ+BPwGzJP1YPSHviaM7BUs
ZYz43YxZL4LQNyTh6YxBhfaIUhD7sxtRUr/b5HiZCtF6t25rnlyyaZZkHOECbRFu
FNTZjDhYmBJpAqSnp625r1JW0NEp1O67LoVjpUEsOVhzv1OHfDIZ6FLdocKztjha
sh/xaecz915SEytuLEijqSRvMOjqg6tOnr0pl4RRtKsYGQcv7OKBK2JQmHqXSip+
Vcccf2yq4HkAymUX5Eiv9qD9+ZF5What/STnGLPDAo+nCRPzde6jSoy3yKIlAnW6
Gvr+VLMVPv4CpfcwDFQInW5Iixb5DYJemCMpZHVHPRdFvmO0I3aNtxSgxK+KWy6b
ZlVSyuQg5vxobmnfi0wJwTa1OM/BGRuZhsAq0O2IPF9o2z1xq7z+BzJEHeOhqD01
BNZa10oZGjEwoxqsyTU8JBcN7nzONtMpUiasNW39YpUBOfEbAf+zb1eg8GueFgfl
2Y32GjwfuZ+8Ehg3CLSIc7yrp6VkwFaYPhcFI/Ts2URj9WgVgqCuW2B8OsGg7Rro
8PNUuu2s+DbV1TWUPDU4q05R9QaO3BtJAozAs4wxqlvuzwKbYdVpLnBt47EUUPO6
dd47VbWZq3oiwm1sYhv9eXg0PK9iTvqIHVRNusdGheQrRBJ8DGsVFO/z299EFsEH
MFGSgdAIRsOwUQPGu3ljEFwL5/ZSvQEQF40ZnDjjZtCotNS5iF/qHNSlRuyv/HJB
8/WWum1bLJ+ZSB/UiVCYjvU+tat4TQKBYKGDtMBzXQBMiGYGXFf8Br8mihKGoS77
wNUbId1jJYfEX+K4U2RJINunXF234GWp3nsYVAAwALJsiUKNz/f1pSwacBginIjm
gdJZDC0zcJklVVNPW2dM2YBdxhlox4oHHX0wQ/3DqOfnggsoNWyyzHZwK8yUT+V4
3blckDMpcZ0X9RbmmgwBI4gTd2rOoI7OY7+a2AYB1n+2bWlfKTkS/P1SV0M1xFiE
cx5sKWSNhLAnGs3zZobNgDfyUCccDScRNWN3QCIlUqyq1yF9Q+ahx0DsnI4gQZgD
TyAKf8UCt8tDXzolbbPyKPqEqaFT0x9FFuXw3UMhHsoh++BZ6au1vUDzPsRNStBy
0jjC4IfzpOoVE1gBOxEFc424uHJAXJOPCrl0ixiJtHIIT2xE58aQv1/07NWMvTq9
6mefx/AdQZpovssyr1RFqdVOoG/1wARD3Lb5siAf7cmby8vaW8z/1kFwDtjiPRDs
BimAIwRckeV7+5/PP4LBvuHRN2oyk4tShMmL4tzzyLvjxuX+i9uQw9WRoTtomsY2
UFHuGDygN+/DRWi9KBfxY3ihQr66Pw3Rpb4BYQ67Tk2IFqVBDC+IfdU5N6K0P1pi
zgj9bNyF0Q2qxGYaq1ClYnzRfNl7DTHI7MkvTMBg7nC4uRBESYLOM+NBcJQ51EEh
hsyuR01Qr27iuQgUsmAM8k4A9wIYfdSGQ/L5bRTvucdjVZAf8onH0t9ohF/T3Je0
a1XCwASkdKDAVEAelRjkWw0gecoRP4EgpJndeP3WxXwmknxenGUauC7k8/60/x3Z
rl3STIid2AXMNnIR6tRTMfXVMu86+Fa67O0weQN4omBS66An+700EzW5AQZoYjEX
HcnVGGq56CCgy6z8LkzifkuuFEDMKE2TIcpl5AvTDbLANajFVShsob8JFam3MQCg
yUQDZI7+emdxtyer6pxQOuHOuoRDjvx2y7sp7bsF/inXgJvqlAINioIHqVW98vNi
UEWtU1TbsKIF4q6U66MjoJVKE2+vIgH4Qt1DBTYRO/R+iLxD397JWpYlzRC9Qedr
RGLVkDu1t0YjWW/H6JgE0tisaHJrBf4JKFkXtA94azoWcJxWmvBYPBpBCv9ITLEl
+gpi9AuqFL9R2FaOIMjxAIf5c3BVPy9oaKDtyIShXTMqZrhAHOF1g82pm2/bzLWQ
WSzhTb1XKJhFuaduzb4jx80mhIYYI5rpQvgTlGE4He/T1I7YS+LYDPQ2h9tSZ6RE
UzjmhlBV4/qUK7qKQ5yY/y0Q+udxReJp4MbXHnutxBkWN1C++h3Ki7SMLoJVEdpu
DuPoADZZGG8MC7b/tc2yYyLWgAGsw6+PNg/TXA7z7t7pfN5CiyzeVsa/ua3krr8O
u521o3U3p/dNINKHKZnmVT/25r6EasWWLoYzQvdG8Be9mnH2jugyQm2/LE6CytbZ
CLzuYXLbrtZo8Dy8+e0p+CVc5qqoXOpFNYAUuapmBlQLhElv+JPb7XBC8X96myHV
J4LTPBwiRQS6KNw5BTo9U+sxbwgBJr18Q1S1VgaQ7RDDOHveFB5sfKUN2Pmcvfnk
036HXJ2nse3WP7tncF97SI3QFkq43qOlXG9S7WRsgob8XTQnwgbOpimZUNYQ1eKX
wcd+Yo+umHh+Ai5Bz5j+onA/sRSW7FPCBagYyaQl2Pe4Ukbyqn/47/8kKXI2KhJd
RXcEhD7KGI8Xi2SmU55i8qBEZdwZ5+jkarg0o9gKpI9naEuM3dPiSBL2cXdlaq/y
4STH85AAHiZ1tDiHDEnMI741YMdGfI9G1bejh6kdROADjKS0UQORSov6HUTzHC1i
b+xcK238IBe5x45J2VpZIT6sZDCVcpj+dqcejZMgJpT7LBgnx8KBzBCOiCe5p5yX
zwLy6c3yJelol0lW8VD4mNHJLgmxVRjrCutdbj2kbKfI+WK+2/ZsAxywoym7R6Uj
DB6tpCb5vXKYDJXF8EVX5YYhPN8nVtJTmvk69hvV5cOXzHM+oWqd/1p3OyHi903w
EyLHrACNVazaJ3dNztX67Wfv76YGTqbaElmyPSaYTDT9U8E/QTAHsXxkxP9u/FsQ
VkKgD0I56qe1vZadEG3W94RNKcrqbjmFnEidQLy5QHlyXFrLIizt4U7L8z0EEcXh
WRX8OyhdeO9FCEMgR9wVqP3Sq854H7DCVasMc157B2MuqVvDUudU3Yo/lnMETkui
yYHnuMKL5rwT/JKmBha5Gjvk2l8il2g0t/FHpydfzPFATF1q7z3/broCZ4tdv1rq
4gH1PdqNnoWUBhghZVTDiAq9/LZ2g7KiE+dBrl5h3gfwIE2bgR3IfAwnImcpR9aA
MfmEGJBZ8cSNyNx5HXRTj2Y2QyHNv4Coj9ZqwwYSCL2vWuCfAYyfuC2UEXHR2gFf
wQyI39PRslswwQpGpzQngSNIXNuuBpKjtsJBQv2NAViqJ++lSFE2OGxX8goKsRYN
ziBZMr45bmYgulEFO/EpE8WHC3nQrKfpQR01jFHjoKYvfSjcOwVcdEGL2J8jqqny
rLjiMTYtLG0cT+Z9AnDlgZNPFweV5j1lRUuxFn4nM8UQlCaKYZZ6NYixQP6SrH/K
x/ibsRHWyCenLdS5iP27FalnqF9T3ZzaLfZoClG2ULPy6k0ZMv5UuELFTez7R62K
hHWMtzdOFaRNrRbv85eZQgA+zCo4wngIpdi+x9DomC/JIGZE92GclH7Rpg+MO77P
IIjU+uCwdqsm5fDly7jxTKrUWNCFtOQ35ioC+AxMNtIHsR/9/mIDUdoOp7gvVj7J
d5uicDaZSKXY1WcWd7GC+OL6sgPoVIJLbFY3nJKrugMbDo/TUJ3ZRFtzaYkn4KYM
+N9B/1xZKfNaTsVhAwA9IQUaoTGb3d1Sl1blgQ9uYjIA8B8MSAJaSEoRE8ibs2NU
ENnWS9O+3oagziCudOwGseDh2tbuCedL8ucMF/kxzhwpF46iY0P42O+tJXK810BV
dkfwATHoPWwRwgeAqJXIjYR02wxDmH/lFNAO7Zzo//fB5Hsz+5I+Fl0wVHARZYIe
n4X25+GR3D1i7eRCk3+Ob5bu21RBAYP+KZG+6R2y+TIhUd3UWwuRTcCSEr70Mn7E
evvsK70t4ywCJWBda7qNFY27p7wD7kSmLa5e2TEG1sTUps34HVdsU/QXixKIPSOQ
UNZL2zRCynl8VC8lmd9T3lj298Vl6LKv9Jcz8Kw/9uV+kqviJ08rwnXSxUOSFLY1
itbnfx6iTqCDQUDGBomZvcEOb+GHE/Y0aNvF2C7190kpCPxqBAug5P79kIYcvn5o
P/FnUZkhz1Mm3rNHGxnILbvOdLEy30Cgi7vGWuRad6gnS5YaWKYtLIi1YEhysxNX
HLU5hebpipxyPQkp/R6zkEHL+dCTFRW29zMccF7+N5Q7gwmH8gOhSgxlkADylULN
GxqgEJVHgJXS0nr84TNfGZdAeswhGA5e6Egyhb2r0TDkJcvmcUMi862BUp6bMl/E
lzPrG6yAziKOQlyk0ilhXvD+Lfaq9whgiHeTqBCLjOpAY6TGQIUlc6KdfI0WsApu
rpx3biitrZ/IW0js0MSlAJDWTQZ+nrjGr03GTL26bxwuvklS3ZPMJcEW+QcuwXuB
DOJCtS0e4jbxplVQ0cNR/gqMwjo5ux39lxfD/VBqS/C6dD60jjMRj0rfpFz/kjzD
RyqdhNHwSSnSxfMauYHkbhRdx1ibH2ZlP2giSwVbIHKBv9jOPA8urT6KLXG4NCbu
PcQmY+Nf27dHoh3oNPcleET9ukYxl8ymCc6kQXpkg/IWYAXj0CNcymxZpp5HCDFD
+COcXGedCZo0AroTwJRIzgqUhU2gtS7Za4j2rhiqX7YQu/SjCAIGnBgG7jdoklvL
jCjIrf89V4kWXey6MoxqpaATU0dPbKi5mkKfkHjl3FDvUJ4mKQ5SOny/FK/i9J4s
S8Qr/yNyaHBJeZJFBQZUxRi7M7ro+EwZjaEbiTXItVvztTQSRtlxvQd6g0vYlHuv
S6P+aJAgyufpUjONQrDXYG28Xh9R7xcK41FRAHDUrOu9XG7zZfE73dCEML4VPvrA
tJxmJJK9HQwI3XEeDj0gV/5E4f1nY2W05TaR82SeqSywFolsAQM70+YCt4aSUUW/
Rd0Cf/Z6i+t2OcIonttJU1RrZnDsfDYjg4nXDv1jaYK42MLIc1x3HcBrSZ6d4n9A
km+pQ9yp3UfzJC8nx9weuo1otl7E39m4Ow4kYHNe565PScmU0rHTIMz9WMCYmvH9
rNDi9Fgn6xkIFeKHdWN2xjFTP/TNfSr1bsF2K9yu9rQF/fzR8SGFutQ3AAp4Nabw
58nuDVw+Inb2fiNL1mpBxpRgTIzKavLzF5tawtJkXTh349de/qjBDAD+PqcTK+Bj
gmclv4A/cBfl6v0EyVFVd8RygU2nK9R1SsC7sRcA/OVeR9uZJ8J3E30jci9EesCL
UDZUY8Xl4X3KzTKhxQ7gvNKl0+mMi3K2Ug453XSeK9fqRCw9Namp5OXIQvPNxbrA
5963NoyP4ykZvsI4VP5sJWP0CPceUcIyE9MJ1CbqTZUJPjDSEQL8oxOy0we9CGpN
6elIM/gktw2XYd6ITlFrF031eLs7e/6n9tLmcg5/AqE3vdVu/DU2rVUfnjghkEJC
wKan68anvYRc13N7Czx9y0GaS2HkYU+yky7l8R79tMrIsB7M8xax651/oEFzJiJ+
4l9v8+ZI9SDarhzeGzo4iPxh8XdPDSVSfbqk8Ndle7ftIqfzemtM4pbO7F0X85r0
RR90YG+CVI8b19ASLudSmmZN8vGip9z+hQELz0+gIdtfCEQ2pR9zkcmNvrcfLYKH
MSyY/hbbRgeGBJGDnR96MrDAG9k5QBiW6xsPmTlJjnKkY4rHYoPcRe/sYu1uSOlu
3ZwZd8Ak9lfLrjYd2sefdwiNL+bhcH6JX+emMCGhwyQ6ewxCd5gJIY3sq/RWKFam
oeKUfBnkTy8bRqXnuhqwXDOczxHLx1NRc3G+JkTJajLHoKqjfjJe/DT7gHedJVvX
TrdDGXR3DXNnGzBDbNUUF9VDsxnB2BJIC4S7Qr7wii6LiuNHrxg8FbML+ixgvSI5
JCaJxKn299kSKsDqReSyTK8RyokEWD3rd2HTxKF3UG+W1g1ib76D+EKVMMS6aoGc
BCDSJ8/m76v9aIdWiFa8uFfwyf5cdS4qsG78k3YuwHKLdJPRnANnfHQaPG98egtp
Tc/Qe0YakiYtj163QSh1KrPJk/tibg9zQ5kywOtqToeT1aFuh0Wke2bt+5ANhzKM
5X+hnRSsfszvuE5cfCmwjxjGUoVrATclS8JJPwA9YJeMehMhXlVXM8n/nRhZ7ZGf
h+tEBDTDXjtxHVc9uDvCJrHJQgV38Ioi4s49MkBqEq7i3L8qV0+PZxf2ri0xShwZ
gRiROt5qLfaGZ3lROpCsU/NpMOc7XnkbdxZq/jgUOmNaoCZJJKrgt2cXshVZwn/g
OLBiqbRsU0jBfU9LGJ4PMy/h2o7WS2OnZR1B+CAGICvxhZkPBAYhqW6Bh7W4iZit
5jD67uBPAwf/YtGhqcuOr7oxR622yo84XQwJSIgzbnOMrMGqwQjohB/uWx2sf9WU
Fp6uM3/KSxIzJQgT6nh5e6cXnSPUqw0Mg74sJ0GazN5Uaedcp7w4oDRucYh/OjSw
kzXSTbURo3VlrA6wsIdkRWWwhaWH/M1x5Zv7eR1uFpRxoAzd/mRHjXV9nyTQ/BCD
WW8YYvXNi4iiCsJHDGXlkztp9oRnCRNoVw5rzhkXsysmvuAOoJ+kslhpq577uN62
QjkLfl7nh15syx+jNfAT3XJwbDlezeTTwAeaFIOW+kn0Rbep7JUaApYuu2TM/OL7
0YQblc/iHLF4s14ZePRhgwiEEIxI+0tdXHQNAFqisG9QsIB0/YRKNxphlArnxZye
aZ8wxsfw787INI11ieB6u0dPNQQxWv8y1i3+IhCpJ2uJoMMw8BTWVemWTEFwvNUT
kczBTFi9PEft3Xhaziif1vV46IKbR9gnSS32T4fV+HCP3JOn/LmNM8HOc+LB2G4K
nKKNC1DXYrmN0pWzTbTDq21yPQgPfMonkQwIGl3drfzhl6TbHSTlVGdWdB5Ljekm
lK3B0Ur/P39aH364xKS4U0hxWg+az5pEm4hfpIRBu8obtUtmJYdwXB+8MsBxsFud
IRv39ksUNFRORXyf+NGrS/TouPSKA5CM5r7mRZC45HyOBzk5NzDODOGrCD/rZ8VX
VqOgUdtqi1rk6qwE6MSxbigznUT6lt6zEBjDdNgbr26ZmhHGCwnhdWSi8+c0u5wS
GQQuPHye6JgPBWx3stt0Q/q7uzoIBqpw5ugsWpIeDOvqCO/ELICNtxjn206saqmb
TXcCpMKpFaqgk8/LU7YU3YQkaFXHufjuzT0+i4lhFMQFkY5MdUNruRqSjx8McLBH
cj/AfOxA8u6VchSubTmoLvyM8J7vpPOpYJSx3RnQWrlVH5UI379B85sW8MlJBnD0
XI3f+e/sJNp2NCXNMrTsIoEEj2XCfn9r5ceK4AyHMk1PVNLNZQcWFeYYzcwrorIZ
tVs249unW0xJDbENdoUKmWgTJMb3HHNEUQP83DkzYShP7YM8ote3Xq7CMgh/DACf
NPMsDlzmTfblsZYvUTW7L79v0hlPxDLCJsxiKzY8lVB1AHq8JCgeZsqOsFR+Q9gi
Gs9uKYwT0sWKCPzFJ5ma6Mp6ECFpOKM+zWMxSxYuSlsEE1Zb6tnXvZrhZmr/kevb
8L6RRtLBjODzNG6/VpGurGq0JiBcm3ZiEqYk0X9NPbp7gmJofUJB7c+FMA+SbJmO
q/WMcJARmNsVCOLHFBEItHUx+nuIGdssJsPTG36iIDtwcCPb1wn4d7mr2t5fhMDS
9/DUFpqts/qmVSWaYh54C2sTfBHT3FkJxdLhDeH40hZKxLpR1IMK8Ah6CUz9xArD
U+EtTu/ES8gI+VlmR5ZuoESod9PkiwTrid2pd+V/W3Q+JRuyEDe6Ivf6f7Hm1mPk
ZAmHXGE1GNSqp/lrdfqIYhHuJtq0V91Fh64fP2RIMd2mDl5wVZb+V2phDGANyA/i
qrge3j4wpVVy9k1neEe81PQp3nS0XI/oyhFQa3eR8KS/WBGYuWUqIMwl0JqdGgQA
jSH3YDzoLWU+3mJjjWRccshJrawdk9cAOqEfMsGchdLkJgAR7PWaFIueJOvPsXao
JP8gKhqrNMDOxHlh6zBRtg9Zg7PhmwaaUuzohH7myCPXGo1za4OkkTif6hZPxFuy
Imup2c3X+1B2pQMUY17dareRQ6hKbIkJ9/9K8XftLUzUH42AfArAkqRosYl/ntwc
g3ZCvm0mEhy6Bty12RpYsYCufSM4tWpiHQ4ey9z5ONsFW3QeP7P1IQ8UJidNo+1y
zgoYSTrCKmx3FRgAb2tGE10Z5qkcQ60OtouSSgOySyb4pbmF/VhjFHG+0vRGEMua
woG/FxReGScUuxjtqKrq8rjmCSObemxeHCVED69KbGYk2MYlTOnwl2X6dPhk0JQ+
NxjyO/XUTqlSxjWG8f2TQRKixawzXL44uvRZjd7OXIcqFxEdvcx89CEyWlXRgWRL
729J7piF/kQ8USAqZ8SkaWcJ6RzV1MIseB/l+b8HaDGo5qINnM1XlGRb7nl3EZI5
tykwecDEMP/zf/wonEyqO7STbtD/BES4hZ1RiYhmdXE0vx7peFXdLiEqdiir+6nZ
Sz47TpM0XC4Gf60x4wB0oViJ/2ZrPcxs8fC85nytGRhx4+vm2mEFo+fizCF8Dr1Q
8yNEj38VFVZOygvSnq37o+dIRPF4t2mpebLSx18aTGIfYFW2vLB0rUXVDEcMogk8
jYqeGKoA9JIHaCp1OB0h+h4nY4ynbKk+cZAf87huegLPjGyoEkJQcAJ+UJICC7mv
gJ22jxETs9Umit/eFvvvd6BbJc+94NYu0CP6hEkdwAt8NTTR2Ar2VPj1xdCH+gy+
v8wd+jKtfTtR+nsIjefjT7B3Vy8nwNZJCD/BUd7+JZNJmgeZ5tco8hkM0/9cvmyi
trGBpmUnJ92lnMBaNuDesXzSkbp8XmPKZlS5/u7DRzOiHFiML6SMHs7qIiwWewL2
XxkVlnyJaATCOR9iJS/GDDRcwbJ3POnWW7EzIMSIV1G2CpxwbRUpKp/t/+BTQr2H
bzzXT4eYtnIzLN2I3n/XD0+mkNqbh2SvQVwgOZESG0iWtD7D2BW6OANQ4GO7A18O
zZq7hvoUbVWjTHBTOlwqKNGEx+lgOe6kZMNVI0PyydM7Rhw8DQeA7H8tbu7uAmfL
h4CWFzBvSjmsd5VXXSgz0S9UnGn9Qr2WRFF20loZVShs6ethc2ZgHQYgeTWvIcsk
WDhe/m7rQjHe9uFOFUJoTTFi8njbWO7Y0GRJxwbLIxre+x77/tuNRabEWLEcIYRw
Kczu+9E7Uqow168BJzU3Jj4vaVWRS18YQ9n6i6x6C32o80h2tCGxRq0KHbaQZJyM
wJzLLrQsWXkIvGOS93I4qcKxCpN7d0jMnlx6AVM3HpbX1i+CPRSlgNvHr/Kwiw0S
ogGdr0R0i09LM5MBMsnFDPBXwWgxGSHdtD9he4PLD+d/9tzIafNQY7YHB49eh/fL
5eYK8tmSbym8BVqN7GObznPKwMnCB3gvgPFjpFLyBNmhIItophJ8p0zlt0fRqaFA
CtAiwBDvS3wS8t+8H0RIFiKfMIo3jbI9HFAYQ98Tj9kMIPD3fPA5y7Rg59NDLp8q
rQyT5JEyXIszjJRGuaUh1MGX6tVd+hKfbGNmzroYiUR4d203H+fwlcCq7uue/+fU
73zaB1R52FUT8E6VO5iX0e7UL4SzY2bycpB1k175a4QjN/zGzmHFlAaJWHCodDyi
eJZBBz/MKGKoPH6TDk7kohLhOP8tn7w4fbMHkj8gsitOWmJqdA1ttmlsluqE2bs5
Ohu0MVCYCRRsxkwWyRrAqet08uWmk41HzEg/sUFrN73SmCa2NQZiK958Ghyy2koK
hPVNEWVYA8iNaAynbsm+s2gXIs5Rg7Yyq1D6WR7YJ0ZKimuLSpby7NC3mMyUV2TV
0U0YXRwnERdLlf9rx1vVP7XBob1BvPGpat1ejDUOlfAJVSmg2dWFjdkLnOCy/8KE
qrNAyCZ0qFd4Lb5OCxCwuAdirMbmFQLbQFVbwKPBQlbAmDsqcNU0RxmzmDPpsLO4
KxEsWkyx6huEBDxoRprI/6fldNW96iwHPGXqrFobOsEU1M70ysGqSsqN0ujDBYES
aIJWfMitW8djDVEYWqvXCyNg2MBmo6ot+irLHjl/Bd6CHPjYrXr725S/xK4Wf90v
odU4X/YBxrCjxKzNjli8mdLY7Y/lQx/9XIS0PugPFOBLAnUqZbeTzsPVHxVPBrkK
3onX8TdVfzEaoRZvF97/F125zZIiA5ulAznKAO8VpizKp5w/NiV1CNCKhsC+Z/kx
9l4PlPF/cKwM4VfKIKpMvp4UapOx98a8ARsbRcC36YHKM0hdCcFqCzJI+enRL95N
QTrX/8I71wsfSFUrrO06xfITlucOia/Bzvu8WVJi4TWWyiqtDHM+gFbIgNJlOrts
wXpSv/7esl7RR8NPhiXg/tCkQauureUkoXyNbOfSaeLt6Z6fSSAq1PRO7qhNU4/r
3PBVXGw7iP7uvBiKbRZH3FwDBe7ML3XhmC36wI+hcoAoMcKXzQ6d3KQOoT3W8lLm
7tJQI8IXGT48QymtNqOw8r+69u84u6JDhsz4qzszCp+T7TFqy1YOK2yzWd4K46XC
QckSrJu6j7FxFF1OMOhd5Q08jbhhCye7T99hmb97rinX/aTy6ae0xbpyZwjRHD/7
Sw0nKLWf8OtLkvmnnlzyxck16w75AJc/GY85nU4bvBPMpaT2cIoHwM614E384vai
4X56XgJ0MxlWTH0i+reQR8/l7gualKfyOJqG3Cz7tIGYLG/hMlbwDrQLS95Gyo5Y
NM8twAijGujj7UmMQKXt6yG0Wgi0sN21fPel5VX/duLcBdnbZDF9uujaaUs28o2w
qgwbqcNpyam9L62YaQJCW0HYtgcI6YcAmFDJ+1CNrNETmDUjR9ZxCqHCao/sY6pf
yjnLSHimznRMV/bWrHI5dRITAgadtvqQCj8hau6k3agg/X6W+GXByCRhqcG4rUI+
XTBcVOSD3CEIM8i2dgJ07GAMKyC4lrOS1+RMjiSKh1AFSrWh/V/ciTzdPTnT/+QN
SY51sVWiz122EcRtTfh+fBH54uge0qk8LnzItMBEyvnSsrldOmYWwgS4RpKQKL8v
grPky8CIuRUBcC0++zm8ebPCxUb1mhxQ9eYyBMKaWg3vRz6UDupbv3aXp6QIt1dR
QmbzLykEwL54fgZGdBejmh/sJrT93MAjadjpYTke976MQlUqVjUtuYM5HetMrIlF
E6EzkxhtxKeocGM8I9fnnBH81eB+jOcmtR7jfe5W5HyecocUt+hb6tcIjr3xWt7i
gr/39OjlKRQfKh81bMWx+uAW3cGSskZppw9OzCJJxDeZfmRnxmVSnAhkYfXxX6fi
fZkztKTSScRSc35AooKa3JMOFpib47Rd8Fz8mnc/kLQMJgA7yUIqv4vHbMVM3g0M
Jjl4VKKyIE6Lp6hLZdqG66a7xn8GI4qlZaLbpqzHYDx0H2t76HoX0z9+vQ0uQCcs
3QiQz06xcSAo0qXcFa+9GsWDJkBKT6w5Kqs0hjnJXFTjGa+EalfVFpAGsVoFo5cU
APH2If+F2oV6ECZlIKEeKkwMvlhYuwxqgwWZ+f8CwQLz4bbK9HDRv1DM3utJE66p
Cpz0eKD9x3Iy9nXfCFqOrv7CvGy/EreVYopd0fdyHmuvCJKZ+TOhX4auT0FI9hAo
BuWi+1CVMXf2wjnWwA0UxYfzHcy44JvzmGU5+o9/y3Do77S3jmt+9mjBWjuL1e+c
PwNLDMPP+IcmWRJHaiRzPyEMKQvWwdqtoLLejFv/xzxtacLduOYlq7W1exrYwMIQ
luVHprjJCVrpw84TufSR2xSLN6VEALtT2+XCt/53QzZtvjdONcL4mizhQHQCMAko
6EEvfAOcCPmXn1LJ+crDwygnWWuPhM2nTwDY39+OynPTFn9Tb0saers7yXYvGfN0
afj9fuZWgUiWAp5AyXhixljLjHzWLcxH78KkwPb5oMvYcN4wZ3DiI/mSpi6iAT+n
RwqtnKt2BILAQINotyem3/+QJ/fmykg5toa3S5kfLGZ2q9U+/IwE6y7foZg7/6U9
4GRhV0tRqihQ4Dr0dD90+HLLvqDKM8ZsyC4mVepSEUjVKjrU8NEqcJgFJBqlqWMV
0DDgOCFCRPPOFMKl7Z2feeXCBd0WBjXvvApAfaSoS13Xp3E6tuqDdzfaCYhC8kkE
vIN5NXV42YJau1+kMIjesJdrF7uKYxaZl/n+eW2pesXGg/cakKb+ZTa6mmEMmRNW
CF4rTIAhsCiOfWv1lNTIdZMmFFH+CcOjQmuR83QMs/0PjG8ZUV/XYGBBL6AGDRAT
TfkVodmhuPbee2uWynzPzLwMIV4/QitZXPiACv4bfTQC/Q8wPxxJIWlpUxxQ0lLO
7fpkL9VwofEiIr3nzVHx2WScMiPUZL4oPRRPKExREWJwUR8T7hL0XdLxz7V304cL
byzdEyDdXp6kaPGbu2LU2ptFQxLlz7qw+BkkEK+X47dSrQaufWoFXhyZkr5rlRyU
4cINNb8wGZyR7fcUeIHbPD1DnWSR5QcczQt/1knBnmN0tUTizW5eo5LPkgxFYUib
Hwgy3U/YLqcGhcDZHnxDL96cqzbB7qvNpJxypf38EotEEvRzvaxwlqFR7cf4cJYS
n0fmad7EhEp3nSKqleaMjhQmc9zjygSfjLPrD8Mi2yHmccs8VXsN5oDqnhCK7Jch
OczdcRKsiP1Djkcag/SUz0Ev7d6FeJa/GvJl/Z+CP0XfPobu4zSEIBgDLDaYppba
kKqY3RJPJ6dlHQTDWRMgI+y7Bkic1nr9HojAl8IzTQ1wNL04tOkDVZHjR5dPZbe9
RFGU/BmzQmh2fIpJeKR7JpO8RqMg4xiIo8Tt5T7mnq1AobM02RE43+pJsJxyHBGx
CO7LW83QlbL6YMv6OpJDkgA+3N5OSa+xoGtzCewqAELdUTVbbxNhveqaYnWHvYS8
oYzUJKTpaz1EaJJhS/nKl6W3N7O2Gt7lQqAuSiV9zhiT9OVOJUuSo+6kR58b//Fb
R2qXv4TcMjerx3OcgeZ4slmkQR7wPjkq+OD/gwQfzUSFrHYk0JFwDdON/1p0L6V5
KGY45JT19MWVGHEx6/1C/THZLlI57JM0h8jPGEViue5T6uATeVSzq+6qaMcUjAqA
oWW8YaLr6VuJG+vjBgRMXe9qdM8dUNLumniOFRQi2Vnr5V2OHLgK8Q+AvucG7LO2
MHAE4qlt1GXcdndrz1DvGvXojCHF6NxKoQ88N3jrFn61qqH7jVnCVZOyNPl7rUyQ
ZayCz7zWveHX4FV0oYPbH/Pf5nbdM/1PAHQnMfns+fWXuCgc863DBM8w4fD4+59k
LVkhZafRHdGPSs9bRV8Yk9kpPMxrrnFNtQxeB34X3DsqpaNhLoHYxeYUP4iLQbJm
GY27OLIZX/aVATa0kun4qmTO9puD2i2loLj07fhyo4NbJiKuO+L+dOEDlyFlBDdk
CL80KxhDEWQkmk7JZO9vdX2uVpnLst4KVFpj8ZW1PD5XSKnjYmTaM7JzX/NAXkGp
v6jvJnN0LyFEDIHgcHwzrfyuS1WTlfQUYR9wTDjX7nOH9YeoOUSaA7DhPNw0BETY
`pragma protect end_protected
