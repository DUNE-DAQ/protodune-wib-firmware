// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dC1SsobDu/dWIoKgoj7ap32thH2glhPkazWfTjilXeIjUMbSxDAsbrj2/mG7Swt3
8vF73HxrQSATsXtEx2YJEac2QizAJU4u3Z+X4JuS3/tyGA9mXVlUjhBvESS6Dlxh
oYtBOYGjgHn0OVCvruAON/CMZbPQTRzSHpIHvVk9KrY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12176)
nyx2EEoZ3lxyGYtH02LrMvqLyBBNLBGldXVIOLsQfZvHgGbpgI751swFilM5i/DJ
DhKeRsBn9JnHw1PI6na5rDteqnluID4P17szHKwUV/97qRQZsfH+t/uDa0Duwjy3
EHodfYAm11nn5r/PEbwv4nn7QhNKH8AxUq94F3kgh/tsvekNsdpc5HgTXQB2AWW+
hwkVrUi/ARaweHP+xl+UPMqV+01yTc6Rp29VXAdVyYK9sAXYpiEB8RW4REiM4uO6
I+RvDEYH7+JFY+nwDd/RBLv0HKSvvX2bvXBam4S3IMsMCj9fMpL8Vcb6OlIzu0f6
OIVWXI/6TIGZPjxd3Rh4ZwB1DFG00pfIrCUoiaRtAGkdOVeWldiM4ZmFNtOA8NKS
HmWZtTRocbeuVkMtdZfXFL1Bun7wLgP34UqXpb9+XXjHvg4K2NavbaedFDQz3jkC
f7OdhThyWhKakMz2ZiJLgTCqGZGchnahV5w6SCKctWwyw1rt+TT/yFxNsaiIsFdx
IzhaeZQooE5rhDQvZyqior5efwV+o4oz58/DZeuONTcUHfy84XZ5iz3qS+l2gwYc
DT1GJz8JBkHnDyJXP4+v8sUzr8fNdXyVPUmMl3ojwEjJjDELbCGencIwS3oXg9T1
JbzEMqCrwtYUyl0o2oA8wOdeDX9WTgo0sGQSvPQSqE1GC5O9PwV6XqhzMXmpabPl
M3CQVz/ReNfmAN+U+OgyyQAm93fDr2NkfeWl4roSFxdQVLhI6f4POV7HNBPlOyt+
FtBkDlxUDRI8tvxYZkKq3IzuEqkgLYiJQnBocrpC+1lnZIuZsGPD07a5LISS55ru
gJcfGSPpa/oweYOdwIiVV+c+I88/pBDuE310fU6pSe96fy1ROLP7WaTR2WIlQ+f2
iotF5wuPEpo1mMmMhJJIaShb+/HOpdVWwiXInkQbDytrO7G9Cmx3VWV77DH6DWoq
PyJhB20NERAYszuc7eIFTZt4fdbsRwG5Fvkqx0TeHQ9hSNsgM4imv/5feJpDk2Ti
Mk9YrHqs5ft3srMestXZCo99XULX4+oBX2eCbpKzdu+o964/Q3ytx370qhMMSeRh
mkRmGV4lGE4d0B5cwfzqxbi5T/ATyDksWwwDeYK/Pwb34rhFmxrtUML4N9DYAgsA
+PTv9Pba+QYNJ1CWep3vfioTn8Ju3U5XngFJrS0DF8aEuj5AmhFc2FSMSrpKNUan
MZEODfJXppBLDL8yQmMXcfFa6cB9Sg24iTbUWPVl2nZkytHdmxB09S9JcKUigdto
9RkFwBkLUzHLF+TSzUBtf+FaXTiZa1Nery8tp+j8WibSBXv2MbeqFUbU316crI3v
kMGte5XRdwsb7Wc2RcccJ1W2M1CaCgc/VMgnqFaGR2Znkxq0aPSPoVQN36y8abrj
PUQvAN+JRIK7MzXmRTqzwfSw0S95ZgUOwk0c8ed0oeQc8RtWD26J/wFA9nsnLpZz
tFDxqhzHvtzoZy1+EZ+liENRun2n1c+oy6dS9r9OSb4dcXoAKNCD++XPPaLc4Hop
BaaSqK7sR7jMOcvS390M1rwneABgq0eDJrSAAicEcNnYuhGWA6qh9Bz9S/X0gMEN
UgwzLb0M81nTW1QLNfeOCUQ0XhwNdLerfySuu6KdKRspu9b0MwbE1FfzRBFV9nPg
4+/kcxf06fm01zQi01n6vC5lLsD7FI4ypJBdH8g/r1YJGCSbHWj09UbUW61F80X9
e6liruBWi+BM3MjOW3h70VlLWYhIs7Vsb0B3rUfV89lkFJevcw85W49U682KomHF
Eb9iKR5rhM4WT0/RIQ7aN/NcegWToTQz6Jgmq5joexOXtIFiEDxA0MM89dYsB/4J
ZJiikhXTPCQntfS3I3CbGTzo1GT2ImncFTgs/pAZrnYi1TZfJYFqwn6GnL7+eoCy
eGiMeCz3kaLiUk0q75q+OMlHtCvvyIdH5IfQ36UOJdGQGpxmBAXWbpVeqmdqkg6/
UfPb59uDwCMC/dgWRh/Tdu+xKNmcrVanMynsQJcwmON4zaHhoVzlVtSRaKMpyji/
UOJKOT8gF7VG3ysw1y6IBQMCp7F38yMIAuJX7kqNVs+K9NeCkJyTZfuu1MQLDmKn
0eci2PAxEAptC6vc64japiQh8wBygHOvAnVJu6UxCrhQf9Lwpn2UdQfxlooxQIqh
SJD2G+djwR6vKLPD/nlaqB9RK08pmgUl0ZPAIYj9+DaJl6wYmHQagcw+Qk62TdBw
4nrmxWvyVt/F/RjMeZM3dfYfHcAvanTEr6o47Hl4F0w+onR79LPQGvhyDPeygf6C
cwjbFoSYjHMP0URRJYg8tIN4nl0LM+jpwqt8C68CngCNscH7x3F4QBC+i26ZEYAX
3zgNmK9FnwsLM7/qntzKm1hr0kJpmgLkbms/ErR0M4aGtr7OiKg0NJS1JgJjj6ow
TghfWH7LmuCRj7kCkAAHNM0jRgiIadRtEmsfDZZAXrFqlBcGf6bkkhAvx7O94G4c
nSMCX7benRcZgFD2cZ+LOgBzeUNOxbBoiDa7xgq8DMk82XdS6+6o8fHMu4praGFn
Xil9Zxf1ojtkK8Ow9Zb/fiP3b+X06B8mXKK15OIi3rBzGAmbKwTQbbYsu6a1bZZY
tEaqwU5jaU/cKKAG7FmVKukrmaIgftN4aJqMz67oqB3kG5QdjX/Y84pO6yK51eDC
ypTqSFLJmsGcuo0tCGRrMX9pUDMxLKhYf+KCB04byzdyvtzraF8IGJpiWSiRwDdp
sAqlhSNec25gGQogzRWipPKZjHnZm5HCjB5fkvsXJwgmck7eHl4ErSduedweFvcs
Ges5/Vng97Ii5mzshpHWWV9wLzTzM4EM8NkJsB0Qp7o1VDO5jqNdvm91Xv+ipKP9
ST05UvMvHjtgo3scc8haDMJMMW7ZryP5++frefBTBKBLwJBvJ3UNsY9v9n0tzpGu
crSpe1ryc09aj+Sx0ASBiX1tuKoQbotee1dhI8VclFAC2r0qtn656IT8ugpwhVk6
3vpipOSBglLFEL4yeXVgdYvOp0oVlrAne1VQXxa9WV2OI7Lacm5EcLarirHsz/jO
KtZdXtp+2CdiU50eT9g8xcTGcraK7PJGC6asyJQIzMwWPP3UNEjU1v1NTH0JN5M+
OtFHwOY3iwvuifPxlJLRNtUhL1r8W0MMtPkh1eqMS7xAGeNVel9aoRq2zvChTupe
PLShJuNIpfSDlzPo5bjQXCBPwa9WvK8vX0JCSuSl9O5GYjEk7dDlyO4FKQRJ85JN
2OlZ7SxHR2UKmH8v2wsNtTBtKPAcXgK4FhrWJtZVKorYVRfKp4V/s2RaCiJwRlqe
elYLKRH9IUKs0tc46PgcH+jTs2Z7e7ayXSv//C+mjcmFK/egiFBKMDXTlmb3qBz+
LlD+M9WyKU0PvMySu0j86UtBDW6TNLij/Tew5TWnkbjHIVV23t7c4yOk1sTMtqah
XBT9tfJkJvFvBm+OxEsghZ/QwgxmwSiRwMN5BtQ/dO6W/TfMCvMcnc3NkrmBwU+z
VeDUAQ9tku6GnpqqKAjlHgANDMx6XzzvlP1Yl1S4q0uQhkF+TqubsS3HSkEVUn2w
6LRgD32pyvFNZg0eu5LwBpKXYjrQ2S7cdtr98kVZLI6c+orJAihZzZ+UX23ODxvi
C5IUXFbaHla62m0ybhn9WhVgedtLZ8ndICF9AAB04jBm5LtViBZ4TiflThl+xIMG
NWKc37jaMFsepPT+UHkX9Ss+fin4w7jTE0lflM2hWku6c9teXRP6J1KkZ+mwa4n+
1v7ZSAHhiZR4+thGblvs9yxaSO6y6v1pZTCGyOxgDrxez8Y/ElPW/9oaJ5zgETU8
8Jh1U59c04B1OJ4ZUSgQzAAo/soYK0rDaySff56mYu5pYMWy/ZXe6CQMQD3JhIqn
6VBn9Hzs+4RYl+/sZrn1VlhKfe2Th4ev1B3uomTS5C8gGkhSrYWBvJ5fPmtih8Ma
1m4whMXHPt4c0XRVabEkOzvYIH6fORe5bev7j1a2ruRqyf3H82Y3NB1vDNdPj40i
bhbwTOfC7Ev7ipqTOoml1oMrIiCAo2Oobn+ZoGb7/c25GUTwnaCOaRCE/tYZVkDg
TxY/70I3NZjHdzpgOnongWtRry2ZE6SXUNMi4VcUZ0RkfHw3oTa2ZIUdVyA+GMe8
U0IOU+2yf3DuGrMZ+1onncfXtRhcYZ2Rb696o9Y/7JKDDHtf8HVFMcvEla4e+DX7
AEq9/NQpDC4pOq/+EHriTdiupAo2vI6p7rwFibcKah6bbHFYeHamBecGLhWqN46P
MCrEeuC2kjnlNboqeDApnS3m2AEhol/q9ydQCVobZgiQP7Jl5AwxJkBejtzzjsU+
vwrpdNvRRJq5KVUgcDBPNDehQTnfzUFspAqU6teMTl8lft1aSytxfqD51EU+jcfK
TGu5R83xkdlAsZbiJVrzbrP90QuxA1ZZbBlEeq0nBy1H5TgZfS8SoO7+1bm9xos3
UH/NnB6RZDYQg0twm41Y5yQg/NIgrg8NSqto7ym5pHLYAWHau0/w2qrtx2E2PxXZ
MwCQe5/08WUNllinlKRTH1YupoWy3anIZTBUG9RpAzgKBCylOa+uVONa673pt92r
LI86dKC6X/lujeCUM5F7sDeux6kOGpQw2xbRsrP+j9zjhxlfPo0YS4gCtBnDmrJL
LQMP1U/dXY9DJG1FoCmCVFLa7IdtkfBbcPAnOiY6SVHlN+gk1rOPfJM34/nkXU07
BsohDoArncQMhy1yFg2PPHKUi+pJ122ifjuBYu8mHV6BkxE774vxOgzE30PzpkVn
Ex/Q3JbBQtzcaHaDBvGlAo/QowVdRK/YZtCj/inM/axsXI9Je/vXrekrqsdXQcsO
Qp1wyVj+OGNV7MhZVWC2rp0pRFWiP+nYBVtBhAB24TYmKlGWRC6pj+r68UAm2TUC
wTmSyCVJ5klrKoOg6hGQoKiSEvCbf4sj42bBp2zYY09OETmwQJxhNOWQVrUvkvNg
dY8x/KhPecoxTgS1ArPvuOgAedIy8iqwUU5f0g/2o93DVjPPjxFjevlfX8IwFKlq
C9XzSMB8RsG0Imd6O+ap87gU6AVxAxQZFTZrVlAajv0o8Ielv1V0xa1L3Ya5tdK6
TIQy6H9fnb30R2oaW6bILLy2T4siG6nYNhsxhQY0V25c97RxEPdA8jlDUM/BiNOV
2CYLIVRtHUtfhEPg83hZQz5+gBwWJw07vWZu1pqd8WY8kVLR/G3NxP1Sj/yo5Mdo
OYtwbSi+DZiCP/yrJh2FWsabu2KFSJSlsIg6hEesa6eWlKeWObxJ4Xri/rSdU3kw
dgL3Ae2QPq2GZklJsfcReCl90lEs5H8IUAIPBhhTvMJ/C4v0e9/rYgQf6C3KHLgp
YqchMEBlj6uEDIytF1ZYVtAjWLgMFtEizye9r93Mg1mY+V3cv8d3m6OYnbIek5Qp
1xU3QPBzgjRlS1/JcmuJwg9vB5ufLNhse/upELhSG540RU2CEI3vrTOCwdfeDCYL
SJtt2DReOzwfXYLRo7gzQowhM07MeBe5QHOSo1L0j43ZQBDECyGWlaG51Am+zFt9
Q3ydlWJZCM0Try0eswXS3eiNjJ3DRfJjeB1QFGXDbOLVvbVk8MceFEbXXVlNJbbA
JbXakJtCH6Jk6CGH/bENTFlTugz3HqROtEm9DKfXML20mC9lgOeKaOFozUzY225i
jT3D2OXPwbbkSrhTiTKrNnatD92nqvqnJD02M/aqZnMZqq9wRGR/8LqnPfK5HjrK
o3lMylD5xVXtAOb/ylcsylbMDu3e2UGEyKgBDk9FKWtpYIwQlOUAi6LA+lU7PoxE
bVInTZuQa5VVy6T+Drr/MVEOesAZXUyms/vFHCFhMLgp2njQIneKeu27et9y8BmL
aPL2TjnWgoKXf7beQ0Evg6n4Kx08A1l0uunpKVV/toKaBUyvLWfTDNX+CwVPieUA
rOXR3WTTzat9vTkoP9s8de9v1c8BSCMCo5RukC7zlTelwJNgh7Gn/biwFjih4Zgo
1wQcGh9WC92XdozJLn13L8AhhcavYzERL6iEc/ukrfn9F/Wl9NaZVL/8MnD93dbA
ubkb6duldOPNMAHkorxS8DJytfTFHZ8dFJ+bhpvq7NUZkh0uvVZAQP2Enek28DOT
uSj8EgY5uKlh5vhhThLM/twWR3vqyylLzIgHa1Lw+aJdxzUSu50fJvZrPK53XXAZ
xSQT89TVyBm5eWv2vnV1F6I8yQpQ08cjH4NC1cqbzfj2WjOFRuKNc7FAfZ+T30Mm
CiEYZ4Q8y7oJRSxqbEKklZ8Z6ZjGRw8gXOW2iT0ff/xG9OjByXgry/H7U3OGUYhg
DG523TCu+55GmHbGrn4y3H9qIBUmpMHgHg3VIPkwl49g6WCQomYUzb9VouExKO5W
dxQWBVP2A6aKOPF4pAZtebIf0zI/m5My2GB/3idACEAfCyRcbx4edXarL582urh8
HlqpyCBDKFuMRL48OrfK9tU7Hl/iHrpNl35PsgAh47FU62Qru4aLksDEX5F5ZfH5
quW+Gf8XpqtFWYYskXIBDc10p1aP9ssiwp89/xeYQDaNXbZJmgM0Lhd6vRvyVR/R
RMUtK0hEX5ej2rKwcy/GLqyX2D4xcjWRZ5Z+7Dcm382PVe0CDABXKM10duWgQ5P0
33g+VoNwX2NLPAXv3o1pGSF1MoKj8KzrohCz0jXgb13YTgjqj7YDQOR1fvfd6jLH
OKPa44/C4uAl0zSbRK7WurcATVN56hPCo0ix8Ru4pCuLdIBj/elJH9zcMiCSP7S/
E4u2wy25YFXOFSiyZ3OwDG4Ym+GRBsUxUVPgsglQ2W2yfQ1cdMBsK7P67fLzArZj
kZPnKVuRUFB6C1oANrjiVuZIpKHyedHCOmdshCvULcLfkqS9thVstDy0VbZn8l3m
KQCt9QSEh8cimHvN65H7LMr9JcZKao6YtJe8unAa351lkxhBBhEe00ePMc840tno
DSy23kekpfiAzlc5nAsd6qwVwOyNFrhYQXI5Ez1IJZvr3bLQ22CE9D/IH+J/ZK0+
v2UmvrqzvR6qGgEvShEIZmi6pZwg/NdLPnkIvCCR+z+F8CVO6jQi5lZRt87lV+4i
FuFGmh9R6pvZ8E8R2C09+lxrRTrvWs6TA4Wb5FUJZaEnfxMzeWK2SLHC/V1bk3eN
NYhI9tJLEeLgxmoQzmj8uZPgFp5kihTkOAHsZuOF3qWY289YvECCE9I3SEnKVokY
6xR8MI7wZZMHBpz/4lchHjHkcvFXt1oaxaa9Ebj+tpNJurnpJGzMoFfT5mAh0/D8
4s3TVx7mHGJofCedt9IFL75rkl+QquR53tmM2utoyOdA4emY/AyJ9agdIAUoGpDw
NNSeWHbVTvDMlLfBOLiDUqVOp2CLS09QBvY18s70ymTiONMuuaxYBhFUxmilIRxa
9daXy7z+bdauStq+Ex09OHdfErdEVOCdSCTixT5tS8H1BDtwY3WnnAT8D8czq4ja
LS1WL2UigJEYzWLVf6fGy1BKSnJOSQPx1ioP/e6qzNep3T5bbD8HvO3HEpOtzZ7A
fMpA1aTxCoY3o9gcln1UVQ3/M725cYxSYdl8cjT+qZNyhjulmJYx3rIvTjpgSo5m
o4oq+l5Vlh7AT5ehYK7rLmR8UDJL0ohcRmQpUxTMCARcAiNJpbs8xH4HeTbD2R3n
10E2PPC0W/j6gp0WyXO6Xg4G1DrT9nW+m9wqR+Gyk6DUQfnwrvIFjdq7B2RhC0y+
XnWaRZhVYPd6IU6vs8zhj9uvBUD/vyqYqGioFar6p20s/9+Ltt9N1zw5HfDBL47j
gFbOK/rWLyRseSubo8Yu4clHD6n17Mnkg9vTIRVPyqmOga/2JhhwDta56DFX8L5X
jIDmSCcQSOMsVutHjaorPgAk+quhQGWbMYEpX/f3nql2Rqn4g2vrJzHSmPaydF2a
0jdKYKic4PS5aV9jAMyeO51YWWRSYKm83OTEtda/mXvAUF/l5f59ONvLQ8qEd90v
PiUOOB2XkhQQ6y/c+9F0QeYHz+JRr1kltnOj1sWrQ49rgP6Ar32RDhkqhchzUncT
BI4h89Z2YgLdX0fqYpnWS1Y4ftXPa0ewv/NxWqHjLhnf64gUaEUyXOBSGTp7Jqo9
9lBK91SZFVnqxeFX8EYB+YCBr4gVbyH6k9I7T+mDAauCj1/tvXP8kK9t2muhhiAL
0QmgeNOdoJdTAPqOm24IosB4v3mCpuW4snohrj/VZYUJgthzSFnkqfqI4TwDrjfM
VLMOXf1fdxzEf6ewdIT+6nyibkZv2CoXoGEH96+CDmxNefn8bNDIIVoUHYjdLa73
7C+AAt4kZhBJ6SVno8frN+xUhoojoyjcZbghAzmRJ42hc/HtNsaBSRYOgzwykxJI
asw6h9Kk0arD9tE58YAd5kdGCA/TfHjV0UtJuQmhmzzOsZOFArSnmL7YkQrwgIer
vZS8juP+TV7182CyLeUofJckiF4QeDZri/zD74VGdEpEM4LYaMuci+bPyy3Z3Sb6
Fm0ZEiaaWgj+1h6UzLY5WnYOtrlCKs1bX6j2gB/oMoFcEi722sgZIRTn6eI8QsuZ
kaHi8n/AP+WC1QdguZaVdFPvohSUoXlofWwIsPOBGSZ4ZAA84XsvqQluTpcwWAqi
GArbsYnkjBG5vVsjL3ewr7FZ1rHrod+SeXcnqJjQIeAdW9x848xAHS60451S7n9x
4wc1oAdkCUCNvz9BjB8gZX84+pJMnD3pdwqvMmIaW76UgiZ57GAbmvP0GpZfNisH
tFcnblIdQkwe2RKmFxqwUz9L/KYJ+e6mPSehAI73FXK1v13S7Lx2ybh4XSaBczfw
ZP1wZmtNihwv4Bp003qlnuk0MpQni6oWxCFGC5QuHG274WpqoFn8O0vm1SlYan7y
pGSG7NXDCkIM+Rd9hLsiTaZw8uQYq02TEzLI2HmN8zcBKTyb9NYotIDk2t2EScoN
Isd3gw4mMQqba0GGB9mGs4pgc/903DOV5jtPJC0mN2omyEMC4WzOqRgBIkkmviar
wgGWFe/+5mAd7UMNFd4zz3/0zTADK7mf6MN8yW6jr0J3SiofoCAx0J3dXDD7IHXb
1+e4uc35uvard7GxeLjob7y9V4ykioh6vErIsV0lXUm503nKU2+JQMQ+bVwhX/9f
7HZuCUp4N8QpBYXH3x4Nd3DVJ/deaDUfwee5Oww043zEDCeixz74iKeCwvLPUD3H
xD7UMIVgdslUXIlrwEpPgSRXiszj5VW1aKyHuAZNnzATanzDIiH5HsbUqmAetz1w
RVJamiYQnExmT4LKqTNo081NCYHYXQDNOy1YQAzOKbV9n2TcbIHqDej+iqBruq3R
11CIREsZgDAcBo/trB/rjViKiuO8lThGJLW4fUl3DsJ47QJTjXkjloiLJM92czEd
zV2E+igDv41xGi6VtOJPRZx6SE6UH0kKxihVCn9HGAyByCtjOmFMk1gMPno9/t8W
zE7uwanQkhJ4qELRaPIJiamKHJeAxJ78HwHBsFg7QPwz/jXulyU3ry/UfzNJX0Y2
ERb/H4b8Xseo7vKFJe55OuJ+10xvID52K+5jFunFp4jNlhQ8VQG2TkO5rma+KOMP
b5M78WwujO19DjdKxpsIc5RxnaYG3TIgkOujX8tEkg+w7jbBuyISTLi7HI/3VZD2
pqw4kmsElNidxJgEd0g7LsAAh5RPQBrfqvUffAETvtkl0+ILZL8ETKRxRD+6lElC
BvPw6R3B7yM7W2wmdNrUF2Wyc/mrhtPj8hJSF+zrt5kBTTzNsTo6qFeTIthbVIDQ
LQ1sBPG5q+hflSTlPyt4JHCtesSPpu90Mv7rzfNe62kW269Em+CrrcWx4j3RhiAU
FsbD6kFpi/vykLKnaY4QPY6Tax0TeKox4V9tGukVAMV/o3Vcjxwz016w0LkGqOet
+rWkgnsyUbbA/C6g5rdFofVv0rMslg5aNLMu5dpdc+4W6/a+u90GQdVz+ceoqIRH
8aIOgolbDONwOKADwgVDlWAGKDa+t+orM9/Qz8UbHoiyMtOWX2i/ClhYHvrwsxPx
RuCFOJAc8e1O9nGlF1OqcLEEp0DDmdGeUt/kD/qFOHPoIWQ5+Yxez0Cl5gFYpUZQ
S+Uh7O62lSjLiuBGM0hcGm9kqD9bZUugh+jFF0JHCT0mIE2Y6+bWVz2JQWo3q/f6
N0ETZvK8/egSx2yze7sNpDL8AbyBK51T6Z6M/WeOAspm2xmZmJBg6Od838OUM35w
aM5Vg7bfbm9x4lUWNmFvkpPX1OCrFdGyMmyIvrqO/ClHrMxRVXwnLByUNRShV7aC
b39wrDHATI6+AY/EvSWuScOi/GeBuW2Msj9+/XR7FSFVbegdYt37FxCgASM0gndY
WcOTjV92xW5UHOCiCTjSRGBFKRy3S6NI8AHH7JaaUVpIkiOfUSO4UWsrTh+zvcPI
YV3Qsjc6nCpKZ9V0G5jwZo5psao1N/Wose88wEpE6osygYq5/ZR5sTaqSDugPyA2
ENivkRHQSn/ea0UkCCaKxk7YvD9fSHSzK3QOqHKLtm2zy3yihJohqQbfL48NDpjA
OxXdCv2iU4DmTaBbKE82zUKA87MtsdDesnvy8M2Q48EAlbvjgyEIlRnXMMxCqxNI
Q0PRncuqozrEGoNcNmzv0M5LN9JCtVXe94RYPWfsinPMoJ0uTHB/fmrl70Ze8FON
LakL/uOlh/NST7QIVOnezwssXbgqw/5AWEisNt/gPTJ9sPduOHOfHEs20QHfcTOV
rAm5EMg2hZ3CKoXXwlnGKFolpNX07gKPW30RuHEUtc/yXkJUh6O+JFCklqf7SK/0
BEMQmuw//IHr/Ecn0EBfYx/IUZ7bCNrix8Z2WrW/iNPskep+uiRE7gvK/iWfa0OS
aah0kIgm5l5Hyi7fu/Pjhilq2eWIUMdl71FFnG3hAWNtwSVv3SjgjhjwtDVk09ZX
k2GSD4QAXjMAI2rXoAPU82t80zb/gT4U/UXYuLX3ERBUgw1C2aNPabTx/I2RJrXZ
S0FOVmGzh62r56lhnPfUldeIgYcwVIHR2xGgcJ2zG1T6YopCFzp9I+B4Q9/c4xb5
WXvDcJwRQTj6SQ5UfJ0isTAhyORqT4exfUMK6Rlf5ARxtEs06ItWAGjy5Vcx/st/
YByq4CcSF/JNq6zyJSVD4eVi+8WslL+CChO0HLHeyNDtqtfwS8dIopoYFVvlEVag
xwCxW65cMgb5jmdLSo35YRHj1wPIHjMhG6gwL5CyaNtASPukgLkT9+cEJveK5h5K
Jypv8lhNqoW3ADmLXVvwR0hKVZJPqyGjKrJ6nFD6E3KxKYn8MWJE6YoKgqjHtmh9
cbPGzxA6HVmWkjJf89jLqsuQVFaDsj3QKaZ2p7vt7da6nSXXnNtJ79R9JhbhNJc/
GijllHF/k2fQ912P62BN5w4fR2HR1WK/cjnSSsXdsCOxRQX8Vq/MCtM6TdfuTvg0
pVzbg4bsb0GgLPeR8rUammDz9oO6U3lr5/piTGbceYNu/h3Va8k/kaojvcmiqTHP
2fvkmCbQN/BlteFBPCgh72Tqo/IGAxbmk+h2hX6hQvWJWy/tna0CX2x+yJpikh/R
FmSdsd+xGro/1ojnRCfZQe5zAFmlXTKR+aS4TU+IBOg2anX6xRGPr8sIAqWeeMmK
60PPS6PFNR/tsHVqJujULYkIdbCTM0HUshxXPiXfT+6E3JcXbwcE7MhAMlW66iso
MKSf2hxrpNvuWdclBIvnesjfxZSN3+vloV5J3z1297P3z1GpOPf0BhxAf5W5q9HE
MekBWRNmED9THdBygMu47BXhXEIU4jbvIFfo6L5GorfTKrcvYiLP9mvdp6uKSmL6
rZ8XpWta5dailbPiv93TUDKF6UXcD7dKJHLdQrCIdmny4sXU2U7h8E4DZ0qzloDT
+HsjU3fDMhW0UOztlMfHhzlkQMbeLWjcDIuY2Io6aueQZHWegtvnJgXETz8Y5BVq
kXUm9/4pOoVGD6m94sJGoW8AbGOdx+gXfOIBpPiIsTwgzqLMJeJ0BQmPKuuyzV8k
fZRdjOZJqbY6JZAaOGQFMm6zRL5MJMEXQ9FBPGZDDVNUvWU3WauS4RJ0Xxd3NB0Q
LCNyvAAfz2U3zrJ6XNL7YGRspwryCkG4KYRJS0fAnVoZdGDh8Ze2T39A17u6KUAS
ag8GpWh/8EZriTCpJLwINOOun63CAJINzrPdbcjl2F5iB86mdAVYLapm6J93DTSU
WO6D8km3P1sFrWruOefDrAeBu7DINQMEPWtgoZShjnciuYqwYWW52XPPbjJ+ha3P
kh6fvBXLjwXtdXwwzP+KbvP+jE1ejykUmwKo92gW83kyPKKW8a7cIM+inpe9r9wZ
zZPOJuH7v2QrepRvJyadRtp4BmGKa9AcNLtxN/jqoyhp9b6519z55h7oaf0iqsBl
wsozE8wKu+6XiFmqW5swjWCRZgSx19B+GZb/j7A6Ppx1nlKU1WmxM4jytNUcHRv3
3RuoXsWuP2YvOBC8oRaHa8jZWuMoztSOXXj+4QPwKHmO+lxSu94xMvTI4lXuNsQH
epVfG6KGwzY03ws/LMhE5P4bq8ySklVV8gFKwH2wVS0EbeH1icXYSGXqzFQTR9ri
GsrZJxTVhjwf2aLJALOw76MSE1QVsXpv7KaDvexk+P81/sTyAbkzvLREHqBWV71g
dxjLlX8pGOxfVuyLVtuk3gqo73Hl2tl+F9rYnlIkoTS5w6igljGWXZWZF+ZeOp/6
jNc6w8VwCM9U8wc4VazKSYcy3lKtfuji+EQ21SpbRYeQUBh52ewbOJonVPLFX2pq
tudCjVzWZ70Yd+YWKvaKtuac4WhEEilKwyJMzSBgQshjanulFCcgP4cbOZ+haYtu
vqR51AM9f2DU7A3do8KQjX3/W6y+3LhWNyBtxajdV9frXzRdEFegbktVqoEqf+Gv
6DF8+snrmtBAzcJhFfbKfBofK60YfvEw0nLh7SKdjtTZaTIG6FCa4M1Xnm9tLo4n
3cytw7fratEO9abxRBoNP1kk/oWSgpAMtkufslsVNu1aaYcYLBGS7vX+bQjUNgrp
SCNNYy2RlgvDcqR8Fh9HxSWk1LXQe3ChIWDuJILvyKeDOkhxvL9/B/6zWha8jVth
KKx3YIRN7CWaHG33fiqXm5GqglN3dNUZlzh4T5e0IWmDNWcBVzNU6cV2oqYCsP9P
WvDA33YLfTLzzzvvzvYqfCHs9AUYhpmPdsecnGLuY4rbA8U4fni+GGHJ2UFmWoFH
U+jZHyH/n3ho4edFAPkfQLukEvxaqSi5zEl1AXeHjS+5kBhsaKnwvc0QyzVnu3cm
nO+aLbJ68Mqe+7ctEegfseUjnc2EMrzFnyusjhttf01GFuWkcrH2DO3/tLsFmjoF
QZ2Rci04YE8dZaZwRrXa/nrHRXFA184dIU5IASp8uHgtd8qOLa5X4gIkS1mnCqEf
ppVqVYlchsoeFzo5a1cE/rrL+etiIP+AHxh2AVEfmNV/xUansKo6Csb+ZHW3Bvzh
ZmGWb3mUdB1MhPcJXTUUjuMfOYd/hGPveHuAhetiKiVXPZcbPrYRu1eP2u374nzY
+ZYoaiFkebI5AmE6N17YMENQLNe/rhtwujnBOioDluSEv1loYOgjNLMuzMClU+Tn
Gdg4ljQpfKXDKTISN2KZFbfKnZvFwHLlQROFq4FO3Iyety8ZtMEPAgCJMDFQSSkR
ySHsC16+neUSmJZGbv92rn8yf3m8JZzAGCMYJ4N769fioq4Au7HORJ2SeJWe93Lo
LxWhfiRosfJTetzMlHfTJenOzrzs5wCoiWXNXINov8GA35b268es9H4j0HsCn60q
2YvXjj06OmUe8ZjO2Vt+84tv/YGSkljfsNYRi6bGGoUFnPrPgbV4D6lxjP1LaofI
ZKScMhSBR4GWv+zEPcKJ5JNpxPiTNnTVNkPq45Ns/LU7YssxX2ji+mypRL6bpr+H
uCC/BKfg1e/fe4gujg/XWxQmSkhH579pglfjlTXQ3GSo9bXJJJnHffdf6ZqViLGL
KVMqxQT05Yzf22H9K1ag1zRgoca66i57revqrUE/rh9D0Ik97SrVZMuB3OiMXt1+
BP/b1TKl/MIDa+gq52rusnS7zQzhgKXR+8xnWWo+6tRl8vUfPdqa4jIDlGbYCsA/
2Y+8v2FR4zCAL4DRyWv2u/nYFbjlAfm67XmqOYQVxZFT3tydPguxhR2Pz9m00M6s
60Hl2Jek+SvfD4c2MLuIz07KoEFzj5R+GFf/jzpxLFE2vCXtG4aGalBuBmjtuFrV
P4HFoHChIhJNG+zdpEHr8GsUCDYU99kBhi4KmDdmCoQ+CbOfzcElehJHjTRHjZWW
fLflBWPnP4mJ+hHg0uTdwFkprwfU1DI5S1MMqx9XiWea85Bkbaalb/D4UOOLJATl
aTQJWZ3WTD6+jXtebCWArmKpd6OecUVpx9wjSmsw8RqnbtCeQ0/tLag9dlGwidE8
75JJPeCfB/KM5LzDkLbGNX3F42lKklrdTRPPjUpDzTGC431NtuqTts7dMcS85k88
EO87rUTE7pk2MRHGzBjygKY4TzWGKeDMq1Cr/YQeEsvYZKMjFF8xyzQh54ClZqFk
I9Q4xiRPLvIDiUT9/3/HoLVQ/P5uroJBvBHoedH8GYQr2ZIKFB6F3pAVCULkMWng
ZgY/epF8KcTAQRsBNdcW8wUntBi1Zv3Zan+OCFTgWs98OIKW7NHNel59RTefSiri
TPqXRy7fpwXhlojbBX/mMRVg9Poq0j05cVO6E82C+bfoGiMv5GmL15hZERvGmMWs
hMwsi5vK5/8xYY9r5TY7PB3x3qSVzRjvE91VALvzGPQOA6NCcLR7eLqlXcJIPsb9
jFhs5Gk70dfg72KTHKtQ6lYfyzfbHc2MFfGSzLEQ5QJ8CHEuWJHwxUHTHxJHZ4Fj
Vtl7+Jxzl/U3DkMKJZu0riXxZ49s/R9nJzgfmK8qfZCqXWgi02ZdZE+2Dmy4I93k
fh9QuCms5Pkc3Gw58GJIO3LdCF+rOi/O9/aEMIppyXPQBc9NQtUyUTeBPc1OdRXh
OhzI9ZH7UyVFkEO2xW8aZh1FewEZxMPFvJ/IVG2E8+Pz5s/be4O9iZdejq/f+re8
zx2PRDMSLvINHe5SXhulPWlzoeeCTeucv4Urwx7C/zonliU9oEl7dEYl3fZI7sNp
tLkvy4hlPHOOu76f9YhK9rzQNjnPXZahw4jN/h2TZDHRi0vA+WmKFJBkb0NY4/BV
QeQQOEwoz+QbWIcsrug/ZIzeDWtfd9aHuV1u6/xkvhl3DTXrj8Dm2fnrzucm3YHq
dQkzGVpiHwxe94SPYVIA2c6Oq6tGrQDRX2Q8V6IQSCwj+cXyBD8G4SYXuYKnNWOq
6Z3icmRCJk6VxmxiiANxANpvDtX+W3QFOr8MgjxH7g2WGPCpMz8En4cUqezLZb24
moyJ7i1ncUk4Sp3zGY8G5e+f/+hpxreQ+5hl8uW9yQIoZ9aNAgALHKy71XWCNx5L
RWLOIdcv0vBXezHCbs1G2SNk/vIdlaP5ZFIsoVokOBJdDLAGz/A4UhAqtONSKUBy
qZUqEpwsMZiqXLWor8dOmUroaXjyy2V3zWne2sM7Hl/ZAb/Llbh8r+9hp2k9xFK5
2VnL2PMepzW2TYkWFSkCaWrlaronrixXIx4EGTWmBd8lkF34KqNX4BHh4ySXJAq0
8u8k/BecvCeTYRki6uEiYPt/L/Sp2fL86HRakcmoEmwYJFdbpKYKdYNsFBEX0H1O
6wl+SysUzmxma1n0IY/xaTZVozaux9qlfizoxdORHM6hKIJhXYe1NKIWedc6+91Z
kxEzZuALM9dJpPbEng7Bh3FGLyOLqmQ92KlVG/IcTF369G7jPusZw6xu1M9fqyEM
H90RJWtuSKLp9Mz18fybeJJTVMu7U48QGZWwZKej2pfY1tnufWLHDWrEIRiLsnOU
Gl3o+t0ml/pN+Vz3SwXGlWac3J6B6VzoKFCH7rOMrSK7K5i3OUk7MI3VwGytiOV1
FLeeaHZasvHFebcDckH5iHnsBzkZubHaAyP8PTPSj+kpQjZ21XxQp4ckrK0IILu0
Gfc+V9fbGif8Rya2mlWK8glFVecZfsQFC4F81Mz5Ts9qgOk9a6/zsb65Kq4dovBy
3BMi7BF0k50A+RcUGgIWAkGcyr6L0Z/dSmfBhRn56EMbrlYbd0DOOgxtxfbhduDi
qGU3XoMRcPh0JMyTneEwjFzmJ3sMfcZ6a7pBEWCILjA=
`pragma protect end_protected
