// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:55 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e26nCJ00jPG7/hpYZfTYw/A3S6jUgU+aGZ/DbPFUA1V/jS5DGZtAthzFu9m7fZxJ
s2xiqqZMOyzxzNMshZjj2XETlPDKPCztpzlK9txUiJVrrxj687IXAxCWajO3HODp
mAXDUmDZ06otUm4RFhmW3qqquta35r5dbG28NqIvVXU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21472)
NAskNf5vsJ0RECZkWb3kGm9F/eEXkN+HbyMYupjvtsCOoH1SPw8fPZ9zpKbr3tRd
1hzzVlRQhGLodN0jIDGU8zSfoYrz1wxXytmQpy245czedKoyUhN2vr2VkwE3+4yu
D2nZDJB/AajibF37PGBjOskrnI1T18JIUjsMtJv3vRlrMmQWwa56XjnqT59RDwo5
B5gJGDDkrxMBeosAMj/LzUybspEQ6nJ+0NP3k6u2kcad8MfzqlKqdc4YCLNBsvGl
NLbaETwGrVfPME0dxAiTujkiD00aqLGC+zhIdPPTNbBIADqUHM8Bffna3A/4ZV+x
f0dxPBlA5o/jIQtRHl5/NwT83CnNfwh1SdBBUsKSD/4KnwVzc0A5JfN7Z4X8N+Bs
c+WjuJpNcT2deDQpMMuMeuJho0pHtYX/NkyMsCny4nKEFid21aZWQxTE5sr6G7LT
NQhDlfYrBssJBcfC+Kmu6m7lxsvNFHOBFWtpKTCe1eK1gLwX4kiZOGwjwtSt7Z0A
EJks0YB5HP/Bc+Ar2NK3wX+wVjd7T7iuJTSM5Z5AO2XatU5zSUGf91u5zt/g+11B
8DUK1Z3hInMwuqNuS9p+HlEMhhq0L4WCRkvDZdi021MM5ii2bTGy2Vh0DPGOHp1y
M3ht/wzVqOkeNLIhxSbB7tSwFaReTKXU70tqTVr8CqXgTxcWqkYfXI2Gja5Ub4ZL
vQV9Py/2nNPhP7z/r5O+D0iebUY78NMH9LMaSIbIL/sd+R5fiBEJoQBaIEYDn87N
EEZkADLmf5Gz14W1FgRBndeuRUP4mLMzYBhmFcSKxfnPEWgx5nfYCcKPnxpECA/k
PtiqjMdsXt7UMmEMEeVWytgqbTFFFeIbfUixER6zVLNlQNSkMphLrf030yE5IUPG
678LqwWCYviTcjpIZNwlCliGM4aAPE1IeDBHTho+R76MBbRf37R3cIQbQA2hOJJ7
pa6Tv+INx9nWJePvicvpUoiWlixuyfoASrXfXxqnDCUjHoITlHQBOWO+qJobIkaw
1seqsG+PMKSudznUiSVtuLcw8YzmvqQJA3WvfvGujdkNy2Q9DUFwFgiGBH4WdSgJ
2YpyAQAkp9Fnw/tpCVaCJ5mdXuhr5QIKXqhhjAylyTWCk49qQWmwbZrJjFfT7VwH
iuCp6H56GnIxYUyF4bU+uH7S+yl+W50usUCMr6yhl0qXtBgtjhEGCyrI9DVPS7yc
8qewXNGdJaYwhl/6tSdLhx8EDHkrTRP99B7e90XpYAoMWSWw5152qDAxnAY7uz/8
w241gakYVcAtyFkAouTVbPphjD+EIXwhO31L1WlKftwWWf8mj+02JBT+s52p/OXS
oY15jx9upRlcUWsoU4ifTd+ZSFxuU1G4rGdL+e3+AIVxPXO/YLxb5qF639FhhFdT
54ZGS4KJZvoouY97Y6+2AlAPZXruk4udN3QVR8sfTYgXAIG9WCaYoWecYfSTYvUt
vnCIEhTB2EtVwgkL6Uo6p6iBzhsaLAHq25ML+fcyywXiNaWDeEvTcHT64RHgw9tH
pwWRbUYHSRUdt/M3Jl/B0Aq2pGZLGwwLEMRDrO9d8bpeo9lAcUBHkZHo5BY/45O2
RetOrTEp0Ujhmo+6lGmjbFpf+m7zDXcanrx0wEmiRiGTmdsJ0hVPACH/VT+phaiY
u4kkUu5hPfwTMP9ZO/sufRKfhns6mXbd4grT8/FnLtAVF6b4z+BL+TpJoaeQBiEN
Q3FDKQfa0EeC4sSc2F5+hO9RDYtO+SQHK4qOYrjb2cAzVEZWFY+ucQceowwD7ejx
gvNBm7OR0nIfqWwba2myxJ+XpS1I/0qWo4qxfoWpClIRldacpukn1P/gHbCi1Gda
In1r7SxZIac+nQtiQU1vUfZF/rJbJT4GkDpioAM4p1VPkkn8UdohRbRdbR+DFbhB
higycSHKR3G6J6vpcYxLeKoiAjzT1Ess92zH4iWw5vW4MU1YWkW5GAn6ugdK8+vB
DLxolBtA9ghxd3Bi4XKL6l/5s8EfDtcmPusuAefGZmLOw4KMzorDSi0gKHjDhXSQ
Ei+DOCdgJgU4VrdhgwWNyEvaj2wR2yi9tRjkFCUcod2cEUsuxLcIkqV8iQp9BVrq
zlFMsLvKttIS2DaJDpT6E5ETETOcZM3zeXPS9fRSPEXpfeOdPVmyUB01FxQx7Pix
BYhoMaB4zmgx3YcHi1mKX9lcC/F9OzHorxl63sdp1Zni8VkQwLQ7dXPWZaYuznyq
dvhsHWDmE9BP0zDBMSyul04wN0eCwH56gz8qrFIhY3mAhI9f/WHpS23f8+tLtITk
O45bZbkvMmX5k8n1CvWmwW0jtUQShQ1k13ngRMbSvZHXfIu1iBIg7gUI6dxJ6O+/
cxZbNMV+wMAV74W6biCigO96DP3rEPFw5aYtcPnMVsGWR/2k+pgJ6Dd3Oubkg1Zn
Gql4WJwjxFFg1uT9tY/Lzf9qbVnnSYAifbLOWRnDtj9ndRrQNKBJgh75gmLDYuvW
itn2Varvz0cbLoEqa5ZDyUCGBfeubjtKmkNLhOpYMPIye7SUjYcK/gzbcDE9yhTp
/m/PKEZWY8Rtaq+ZD6qwmk8kaMLV1jIzQ1ww9+21LNPvs9xXdOEWaU9/WtCJ85+S
pJ2RIm1V9J5+jAnXPeIkE5H19I/2tNJaWAOAHRbQszVeGbBKNIzy/ZUtyoObBcZ7
NLMr+VgSx73Mm5gr/N5qpFa0+QVEds1WFoNC5oVsUJiztAHDB0J1NjAFqct/dMUv
hCGajAp98JRSQPlH0w1FLIvEQyMzMSpsUAWdjjiPHhVGhW0B7ShWzrscJhhM+74o
qj7DyCVa+vloVLZB+cBcDRvoY5I6xpijsCWDUHlS60wuY3yPj3BVOAJ6gLnVwRUA
cnfVRnuUEV84nDAdVWhvAK73RZIcbGfNCy58AhExDNc3HfMFVF2iFD8qWBh01w0f
AH9VS03vSRCjNL3FxPXasm/4PeWpK2fF5nwW1//fhFbpciK2dFO3Dj+OI6IbfV5h
ShNvlrhAmaqgI6Lk2lERlZDH7+1LtJ0U97hAylyZrlLNrEiqHUoz3l8jIRnQsD8x
eWlhPwJ5ByLS4IYNI4/yFbVFXr/9qaBcTz+is8XrE/ieqy9IdnM6yEzGN5Magjbl
6tI6UnJE0s/bnlIr2zsVGh8CfKDEFhLlugnwU5M04wEt61plo1/Zu8LzOGItTa/D
nNAzPL/Z5VoKOLxV8EUZ06jJOzxSguIMAFl4pCk0GfbQfIV13LKdyFq97VBdRvqa
Vott+cSBMyrc5G+lzttWzwWsh/wZ3sBqG5sAJl3AaY04lMC7XBraLHNp+a0dSxu9
KJR8pbpsDE4jshDB4E+OH4CGJIDFOvBgd14k0rziFZ6gfpbH5EI9trlQ88rabEN8
GWci4TRsXtskH8M9RNufphWZtrw2MD1BVK9VBhcGLPp5B/aCC+CLdAaX2qjiA4Wn
9PMw1HPOClEb+2MvM+gxdRvh3tzEscET6WmWkjLlHS44iZ94Ih+BSUYp9mKnn9tb
SNv3m5H2djdYXeolesmYNmbHC/9y67qmhLnarLzwY19lQA9iDnJRcs9GJlSIkJKa
x5aoJLbIJv6gi/Bhapb5VnclJCh6fPGABzt8T5t90U1jxtvtlbrbqSY+1CG/b0/a
MDX0W167OM0dkvq5sMFzFeV7g3MFFmZnctWxSsDHTvkCKvrNtoaSDsTK655wYR3Q
rd1VyBn9G3ivCE572bcVhbALXeJg+ffjuy6c+DOqu8/3V9QRNNOISfCAKTZNYHVQ
vzUkxA7+cPCBR/ONCWlbhtAHL8VnCnmdKjMSifAiFO2u98xjs2HhfgbC5Eg1Jcet
KyFFKzCAgtiJn6nnTI3tzsmm7yi21KvJZlMPNWu5Hb6eG4sD8tl+2vm6QkD89XAo
+OcgW7AGg0o3gVs/eDjXvnl78Vx8dxpJAGx5AB1eGtmymEWJyo/Z5ulRGAPjSDGg
fMciPnDs6dlAs5wbe4OBc61pGFyu5oRstm2CE5syf2RJDCS9Scax/JaVM1rtLDlC
QM8NUcQBSoqWN4q+XjVhWQvTzJFkFH4i2PvCDoBXedAGBt1A8XJf/Ir3GR8ncxUy
E/sGfP9mGViZV+qRGJa7Nx3kUMkc5JqmMxeKFs440uFbuOk4DZ+EB4gsUMNSYIqT
8lFktC1rvWyMUesOcEbmA1Vd6DuZuDh/tc3hWF+tkzfkWlofouc3TmQXb9+VqAKT
6IWSsE9OXGxtet+OpmAj+OlotqFq0GK7OoUxlNbeYTdkMjaujX0KpTuvFxqlC85v
V2iu/g2zUvaX65SbOqEQ9xz0Kh4e+NbNSzGlp728rP3U1rmrBh6s7EyTFnILlsmf
LyWb8vCbmgAokOUEBsdCV4lvFVfx1mv0xoMTu+TQx2D0q79DbcXh01fg6otQKGMy
hYjiITg82D5b1Ht3JjfimJBFK6p3lNsa8Uc2FbXhnBzV8iGrrmjY2jpDVTxoXN3V
pKRaYAEKXg6p9zGHQEt0xWDplkmnKee3Yn31ddBAaFwvOEGmnZ2GcvQVCmI4iuhw
Hy6hcS2Lt54b2ckJTbDJYzkVuWMXC4oRkXZk0ANihw0dFDQ7EYUbxZE1LgWUdjVV
Dz6X7Lw+s8EdAVc4bAcgggtiVypCiwrX/+rJprYfuVi8MYuHF+xVjB5t0oJ9zNoo
fYp9Zi0ERHRsHLWuQhoGUzzjj1kQ0wgxCTxcq84QiQPIke+prxozH5IfLzQDgex4
s2/j0rBo9FP+/SscrCwCCsHypRSZEvXO3hh9PGEqq0ubLq2EaGJbTzbDNfytv/Rk
4QOrlpsxhpBwfoEZGzq3NWmu3K32B2yO4LtJ1ZCSYmBo7UEFFkssvXe44/HOXFYz
4Efz4wqXtHRFHAWRtoldIjwgcVZLNhzNLHRRHV61IfPRmfd32TeJ42BuSEaVN16g
yL2sIpufb/FcLSwJUaSMnoJMeXMpoKTKRv0DKzgEXDRdaIF4dZZm8oZ7GUe8HCsT
QkSzq5uose+Dq4gccPKVZNEfsU0HrhRcip/yn4KTfdK2SAk3VXPrVjucwe5fNgMO
jngT2GYwKkNBQ5bZSv+/JPfp4tJpU4BZeRhH8Je3t399TgRqFinXKG3XeyJSDCvA
poyOrNxcPh9A8eqEzZbE05hnhm3L4SzkswlCrhr19s1pHXWqFcJRbXUdUSCVXfwE
ex70dT6zu4eN+mSpJiSA73I5/k/KJKyc5gSqJMR0xIKtwCR8etGm0ToWyPUwd0PF
KGAQsjjMUDYsfry8gJkCh6yzGfaBg3cVnR5mlgwLOBE7iEz8Y4L5LyG8olm6NDIQ
CciZXmkyutof+VBjWulK1l/uYTC0Rn/qMNEV7QgUoKgrqWZ0dpnVo2/Hqjdyk5AI
2A4eRo7hAji4ntK97sT7S9NiRMZ1WaT7OHCh4QTCpot4DjIBVjWNe+fFknbvflUb
BbSCjIamnLbeRI2jPKd0dLI0Ne7W0A+GU3ccFgzEO1OiLT2pL0eR5K7W8u7kTmP1
sExVHm0wY4qb6cGJsv2RPghTbIsurgqfKqdPmS5wk9qxS1eJUKAM9NFN0lqAG74O
Bsbhc6i6fN/8bowynwqGsawMa2OhxJAVwdQWh1TFIx62m950c97eQkpyMCKS5PSX
AYy1vxBSc7W3CriTthJqF78rM7oLRD0n1gmu8XY0sj5L4NkcLNaVqghwRO8Uxnxf
S+Q/iXj7y9reyX5FVhO6QiS+3onYVsnqcBxMIpN9V4N8kekKDz/PQjYJhDDbvZ1K
OZNX+PMlPvPSLznyFd5tBwUDIT3JSGoiT4FTCbsUgcm+H+W0N8C7w4cDLyKIjnpL
8/WNYQ50oYzE1m3e4u/K/XLVgsNexJpsbLHNN4mcH4eQc/0U/7UOO88mRt+bmmuM
4HFt3ru3iCJEo0tXMooYydR3lXEVewF59Y0bXp0ikkmjQhSyaoweAO166ZsRQPe+
mX0NiUqnD8/G3t3jSzGa/LO3pERv309nZQfc9fiudlhlznkWLsC9v5KZRGIagget
PumFf9I+DRtXKXTnRbopHt9li8Q6LT1ZZKJ209bs37V/GE810Km5k0SwT4h/IUSO
8dJQaOkfDM33pQsyfUwlU80CnyYzo+iopBkYWcm+jkrcQtbzwvIEGVU5Mc4I9O9i
OT8MFmxulcKXW8ZwwSmol86i3Rev0wDtWaIFMinslhiaZ/JXIER+B1/JCBwLn7GL
F387DM2vaTS5rcb7E0e7TdZGaqNOHqr2OScplvQ6ycufTiDJc97/PKAMS4N0uGnB
kXvH4Vji8Z/E3NRuwOMmV5jFlQQjehCtMltVMyz7rnK0WBX0L+dO6EEsPU8H7bBx
YO4AHtZOZL8Mxne2whJkbA+0VhynK+/lvHb6E/Fjd8uovK0aAsaHU3UIn35jCFel
PazHGB6bAi5D8c4oN70l6xn2Sm5vjk9vYC6BYlRjDA2hDfmN077+hs7WPNB5pgrT
6+KxfSIdirwGnnhgvtfPiAQezYGI1STpdcMMpY9AZfypRdNiYAHHSq/qd+kl3QwU
KP7fgX/EUwWpK7xQTLiGdSfbioM7AWo2ggqe8zLioath471v1IfGolgsNTum7Hcp
ASMic4DtPWqmJX0EjtESApOdsrURGhD50EJ1GZbQUDTJQZGFKgOHlO4QKPeHvE4G
fJEZZlQrtVPUZ8KqK/qxy6ueX0Bai5geT0xObT2SQcdyaag5YChDNJI7bydnyMSU
PISMT8dlXrTbwejB/FSlXru38pqGabkeJ+A0+69kWZNtjDutyzsmj1b2/Qt5yOsa
sDVVRfoQLlULG7wH/8KpisygDbX6LRKQJTjI/YJoVLSPBdKAJjWCgNDeyMU3Io5q
2bmORqy1x476B89koX+BLmx85H6E33s1SFXN9+WJZ2l9oJ+XYtPRBlLxyCc14anr
U8Cr9MjC7UHWhAoaxgvBJdlKYgQe7AndvwNu66pwpTK0gSU9u3pLdumpf6uKKW+W
GrCA5zHBajChAcGPwfhyEZEGjvrbRAWdT85ZEpLUoCX+EkRHrxMbZbQ6vQa+FwcP
YqA0n63/iL9X43Vb8LW/hzps03ygnWVpmT+JS+f8i3Cw2O7+zMhdRQMnCiBOzU3q
zQzW4xDfGpN9aP96Z+8JJi1v4Fqr/ojnUL7N/nlEeCyBc9HX+EVIo+Q27IDczPHt
jE0BQubku0GnPZBwZqn4IZPH4By1Fu3WfQoMxk4BOqC6R6dwH6EG7uSvAZUVFInJ
rZ5bwLwuBF3FW2dGlp9lanb7JeedFBtOXKTtOVPXbk43u0mIDiGy1ZkyqRxbErN9
WsO5ACGlJrjvctaj9khKep+ATMdTypWadBjNoYbmJFpsh4Vek46/dLODZNMFo00o
ZsM7M4y+/A32DGskOvMzBOCubnhraPtiGHx2c3VewjAvi1aoAkxjbjQOo1Fm7uau
+L+WCafoMbnFi+MvvHPHB2RcfszZq5GWMNNCP5VVMs5JfsNCr0M2+rgBOpIKx4Bk
BzqDufiXQ1pBPexHkD10lJckA9GeBynVe540Qs36Wru1IkSzviVRanNEcn1CTij+
1Bvj4sFTngxtNxWFOYDaWOXcCmKXNz0ahkF7z4AgD0lGI3XHdBBQKA0tloOWphKv
kpdzTs42MY+pMn8GK1v2eX9oAubtjU24Iwww9QiwGt4f9c6TfrRVSHW8gyGhwVY5
VJH2oqTwg6fAZd8SjBGS7+N1KVjyohC3a1/YbnCnz2M/4bD4XSQokOFRaaSvwO2U
IjjXm5M/pKK3VElDPp90XSZKsXhQmq5eA9hKrKrXIxChJPm59PCJzsFmrzo7W03m
DTGgXtR62q+PteFKHoEj57g0rE83n/8bwcRtBu5mrs2eA60gbkrXpat6ZSswRZAc
6c0VolPbS8hrSSsxwrZpUOrT8P91EMAI+KpFbegefpQy1KLiDUqhMdsZV45WryHN
y1xsGsjkpsKySXjBxwO4XXZ4EOadUXTHqWujzg6HQpf0UEi1nsn5wwsmkvu2Nbr4
s0BagwAH2fkEbhNf8LA/b5IhxmWx7MP2J516hUpnOoBBGo+XIbm14fRNrcQmNOh7
Q4akRSE3Gndmbi2LftcV4llcuPa1WiApkZBoD8GaLtjy0OHrfsamGE8FEa5o+nq9
c4Ai83RyZ8y9hOMIcmS6qQMTQyo35rXiLLTcozIzg8zPIOjImMafJeVdzf5wvvj/
rBVrlAi2aJhvQEAaPnQ5x/7Il+PZKPUjaEF8YUuRiENPPfeoefYgLBQmfSfQWa8N
ZqFclyD7RYgIDd/ZR85bxOx3isrLzMA8k+l2JRL/OQRUglmA/AqcEe4l74m4y46z
8DnhwU4Zhlu/kT3S91w3mZI9XUkqRtG9Zr7kkm7I/MW/6KdU7ZSfa1gnfMvuy2P3
72UDJGEVjR0YUa3684gt7sNoT5vTI84qe1/UBb9IDUO5c0jpkwIHP0/urCjIHNZj
heLGwysaZVjdn95tz4kbX1aMBKSL5xPujZD1fxFi4H61iy5wuATGLJc04OZSzm5R
5gYmLlNp7FGyc1SO4W1NtRv3vDlsBjsBo8WsxwGJ2O0/WWS3izKmZfTWcmHNfnS2
+6+0MkfWmUWlkMuaQpz1TaGENp3ynwhpPHY6afYGFl0rJIdjw2rjJxXpBCyYuMbN
VJSD3A8jZ83ifSOQQ2pct0iKN59/wtxJlVPNvLMR9eIPq1lfeY+Opz5utiXYlFyO
pULUG5YkkAoyz4QaAVPIrwW6RRWUazqfQADMN+QM8MtaYdoxBrnii4gM/3vXjAdw
jhsWWaQfFpKKWcOAE5ODLVmnhY/iMDdkoiCRL0w+7U9CWPgOWtMJYTPNT0XpraFr
eS3zLSVKqQ+9OOuiFm2U0cOrA8ktjpEC+TKuxHaezCNkSPA7An4/+W2KigGbGGkG
RyLTuW/YZXDwc6akUJ5+QgyZLMuUMm4ifyPSYIeG3rH6H2TUoLBC4DunYwbeUwBf
zeRPTpDFaWcah4k1l1D4NYIBHFiqhVk4bdQS4IAYW22yU+Wa8KQrBwL5NoUzwqJz
NOHsu7SR9A44ZR8ecSNS7R3GdWArHI6+PePjlMWqfQoW4Kro1oqEqiGjxfCa9dkJ
hq7nWBY3jla8B2SSeWi7m0JWE50n4IJ0ZuWLZTebifii6JExNQ7UbPiJjRXyfZcA
z5koP8RLtC9VjdrGwCMVaBvjpyA5m5F0hx8HgvrEVelScLPIFJAW0DgT6pG3oPyQ
LBH1nd0S520t4uj+M97l7+tDEsqboOqcX6oE0jp+ulenGFuRfRUdlVVpBUcpIVNd
uTsw3ld0vITuDYA4Rsw9v0eWMYmvpioq75lNbGF3gNCJUUmwD5CUHqoYjWk8zfet
Dyixd4X8uLPc8tu5vlTzTs5aZyIqAJkIOSkuJIWbtsIXVV5W1GGBaPwkQaaC3DQw
GYXw7pADRO6CtvJ3kG0n2YdgZN93RXIjD5/cM+M0EEOSAz5vxr6nNpkKUNEHUFd7
IUHQID6LvKE0EECX/O8LG640FXFIAZyo9eteoderAyeuD1+pB5tUjRJw3FyfFf+0
nKRmpBFcQr5OsV9BfRqd3dbwzMxZ0lc4H+huxl4i1O9mHVTU4Fj5y75YzBd4R9eL
oqpXfb98XRHCN3iuHgZjXbRxS2WLZP3Ud/FfJEIAIz1LjwRVHpPvGuZ/vSIlKQH1
sE2RYrYP+hNiE90YGxaEbmhRPqhTJVQJUwUPUU4xfMpb+ZyXfSVTHMAGTXEcehrU
zJ8w2owrpj8muzXK8RiUT5sz4UHhO8/Op7pxivz5KEgOUGPQGgvji+YX8prb9Ha6
qD3RrgqLyAbHj8oFezhHszSfNXt6ghtlwXU9+czVd6/89fvmoG8wNpGBazMTxJmA
cgczDfZNXiFutSnpjaI28ZcNtfE/VkKvlSLCZrLMJ3qSV+BiZI5Kn5YKiIffmxRu
fA/BBWThrI5w/SX2tGfKiY45qJnsSKPlDVqswMUGDjPBXqTp4tbFw9w4O+D3WKVC
hdbyDXrIT5nSWTfdWLJpsCnARMOIn1Mex0ccEcAr5VP5gxe4c+2vBfx+gwGOHDdI
Px3sBmE5rOwDVDBQRhiajbpfdsppW4esFRp3Nj4Bupnp5P9jRD1Czr4tizAS3NY4
Y2i11NhFuBytuUNvqc59gNsKbmQqsSCWp9WrDOxLC7SK+YWfTwVWUf9vTpZYG05d
VEdqiIZBk4NHdK5EhjaBBPhnPTZdNZjOC2vWxzNV0enp/80h3qKBMmIZF07P+0Sa
rTTrir272BIKUH4Hb0QVCWRcwZVbIGt0Agvs0w1c+baV8WfVfJtFCyy8zcEj0yA7
ZL4WK5/5QPzDgrT3CQZFHJ/ZaWXrLkruHAEcRyFM5xlASIYau00/VRfaoiCKslX6
RFuAJnF1DSHtTYxkO5o42P/EXQzpsP+kNszKbAWTMPQ3udEZ+8VLmfe85XRl6AcU
Rse+q3LIrCTEN9he0plPuf9KydRdcUq5O0ui8IVvtAa5k0qGql/FUyT4uPooDWzu
cytFiblG/7Bn2tYcC4UOVKIgEeS+eB/+VHSev1NU0NofVL8XV76J9lxOv9H848a6
QYQRv7TfDca8j7KaFd2hMt4tcwiMztQE+eEqa5Cw4BvC5lYaot2o6OD+rTs4Ksrv
JusQKPkBrJwNh5h6bWbE//QHH+eujMOedtFIFPhjPaW6A6odiDriBWRP13KowqzD
9/AXntg/SqVqnkp/jKP5x1fa/d/T8qr6UolxRX33b44JXuBqWn/pfEVbirCFmlog
/rsqVP1Z0Xxt3riqSLA2gfg7Theaq3vPW8WHvKsGmDFoHFVCEdLlWFDGioNzBQMD
4afPNpfoC5weZP/TICm310IOyphU0y2ZetquT/X+r3fPnGEWf1TdsTZEZdyDp2sq
xlWpBgZcx1YVeo2O6275ouA2h8MLta3oNofTzp0uZsWImzayxdiEdTFhAF773M4p
1LgUAiUn1HQLJwDZtW+Dgrd7q3pQeXyLG6O8e2ujQgtWOzddBfI9Yu5Kt5Mjbmop
fUhtMJftBa14wvsqPPF1YnwgR9SugjxXdq3eH07of+3lnwiLXzR9iDy3dAi7uzyu
FxRtCBZ8F7wtE58pEvilbn2+Hz+zVX63osNNDMT86WZnzkzwB9P389DgeEkK2xXt
ljZv0Z4KuqLzLK5yaFWxWl0ZpC97jNR4Ys7QEIHFoZe5gP/5HoDIIw4zlNtq9AdJ
+YBe1mtYWVk+5ZJNgdJBZdKBNFprWOdqVEqIXe7olrylaRPAbA7hoNlwrLZHQcTn
bPUsLzRaZpuLLqXjatVJLWmljRJTTZjkjij2aeVMvB4lPdG2UyzzzS2cJ2EfvsKu
35B7ZzOtG5Ae+j948sWhnV+6crqR6eBwvnKlbfFmNz+L47Ll1fVwkoXaMZtQdLph
fj4BvfAp5lCGr3YNgDE4aieCHdmW6Gg3wflyOEYpF1F64o7nIFcGqWo+m7N9066u
4sV85ApF9uDpAaQ0CjTM0UnPX9yA2wP5u/9Z7B83zsvVKstkry9h+iAUq5qawk3c
kgtvbgkZC+8zbVETtSsOi0j74623XHLVTvv90SqoKhHp6ERV6IBBQRp59996zzwA
JCyXpm62A33OC17bQu50TrvmIUn4qSbqM/qsicYCk4gSGl9F/H+5TN/UKhn1ECl9
VDTbOK11ZlnPRB/ZMyshI5qWw04bonPBjaHeNV5Q0ztXgVmmsfjZXr0bYrGr29Xc
nJX05BxSEeImCF7p2MzBSQegG4mw3SNRfiaqCbu06OvCmBF4c9KEbP58hWjcPsO3
mX6S1gdBZPrVh+RM4Wa28lITnbSbqS4EqWpeTuJG3XT3k+v9Pya7gu16b7j45Ah/
cTkCH4EppBuw8K3+xIxDDaivTOPtDi7iZgeHMMQw0VSiQ5fUjLNtE3Cs+K8AoDq3
s9YPv2fG4W3u0GxsApV2b5byCHksV+g7y3AwEiOLnqIZs+qsYmK4E3fLcH4Od9Q4
Uh+1ZvbACrDakwHOJIoixz8qjp//oZ09DKcbdnxYYNLm9KyNevduYmEfMoXtr6gf
ZOoy+Zc5WqE2YNdcv8NrPpw5yxXzO+eTXOsXbOmlKtlXeMhq9Bzq3x60z/7v8Eag
lrDXGmF/I3ViU5PiA8wqN7JudfgoOf9EbgDICiY6eqhA38yWNkQvvOV9a60iiBFs
Y4sY0+aVu0qD85VE9UIakfx0nYYIiOgmX0bX5CAgagRcitbYiKnAnXD36h7ullCo
KGIAGE2oJpWNuNKa8SUjTQ6k7EG9sOoYXFURvmLqq2yiFwWG2vgkC57pTTs/vbEM
8yTIFxer+L8rlIZdrhQHBGJFEQATJQRSe9vKv/b/cG6Ae065UCz2/dzpFO8ok+Oc
Fc9bc+WNQGDg38FMXU9nNiwtS16p/CXaceK7qyUXKLauZhrZ8hwT7Wt8ase9l/R2
ECUx1dlpEMBg4R/cmbeueMfIzOv/6Yb+0a34g/65fG8MBQFpx2H9g8viz8+vbmdE
X9PVxyyHmpgTIqvshjzmi4AIGlGnawlBrWgyZPtgMgY2HoowiFquyiWWFOnFzDhm
Ga0n5nCK3YkcFhJKPq9IIV6rv9phZnCBO1O5ZCN1TxcObZ4LR+r9Hwl/nbJ9rDqk
9mw829337ehsx5AKzqRXsxKRycvMSv6a4lYRwYtkmoDybmk6CF/R6P6+kLso8pm+
udRfEGBAVD4a59B0uaL0fBkyQV1pYza1hWS4oltIu0wEYjuvH1WdekeVXIwveqNX
WT3vUCYYD3mNbDa7mxoxW9L9C8SBCecmk8znwRsw5fYNdTj41xKfVPer/TXY1NlK
SmtYD1ReBzri70x0al0pGGVZOUflQoaYVZozXEdw8uo7G6OagSnozm9d7QSgKYop
+1bHRVYTFjCbRUEZNxcEJRKTujp0atNm+QATBWRibmW6ZbjjqSJWSTGO/ghlJ7vr
d2ZiDrTSjuuA+3ugw4RBplP2QhbnaydfjJ7MWlPiOH6K59x/dpB7zFJbR9ruLpf8
aD0gi4UaKugN/vM6MQdgf3tK5qiNKDgai+QxfxTzsg9KVhreSiYhCOBOrvw8klrJ
4+FmuQCBld/zQiXukkhzYMUhii78VLhceEgH6uIyMMM6BBQgWAEg/l2U1tKbmV96
i1tZx3Vk+dX64q57Orcin6QwNTm7N5qJiGeCvLsNRQ7YXhAEJuZkj6iFiLxGNuCP
PqN6DTsb6QyGJEJYElJH7bNEPz5wSXwo4F7PRSx1JZcY1SHQRIz5YLq9mvdPcxHf
WcSFmXyww1hF4LM8h7hCyGJdixGtupJs296hxXybZ4tYR8zt38eLPwCwSqVNoJ1v
QtAmL8akjio1n0XM5MH28UMWBczbfA/3PccdnSR3mRc6C0lVInptfBZkuibrXunH
Lz+OA1+nrfLPKsOKiS6nYInLudIHUFvCTH6H4unjuv0WGFsG/eRxWy3FGa8FdSji
BeCKP6w34pNr12+euAnOKQhjiozXFiBHZlbEVFuOT4nfmLpkmzi9dUyDM3Yb/Mgw
IeYS0kTM9ceW3w9nk0Yh58Lc/FSPisYkyUK272MKKO0tEBBCcRifVuGTFPZeHzjt
jbaf6InB1mtRHn/fV8wxDXhkjvRqIsUrMh8NYW+g+Jr4AzJIqEf1TLFwgfp94RdO
oMRmCtwRtBZBq7ynIcPbTWyI0nM8ApGmLorefFZJ8bloRoFOVfArgu2euY3HISaJ
hGrUK5JwfqZDBBpn7n6UZVePWUtZUUGolxJ5X2KAQe1BFHkM0dXKnU5vkmEFuuEk
DsXPt0e79bAolfZVvc3qbALLU3SrDp8eSmT6Zqmpf2gXsGztTHMOE9xQf2Z5DiE5
CELFEvWCitwaBt6W1UlyS8sIUyuPzOeORpJf+mAWOM1qxF9m/YtnL+4h4ZRUIr/R
O+kZrwkDoAczYyQ7BoN7AtZ2aeGn/VB0HN2oM151Ft9RiGOmo7zJhYe6XX9cGhB1
9yo30KcWI1ZTCoD2UtR71IZJJ6q5B+divPF1KIFdYlRNQ8Gnw7N3AHXZRTMBoqcW
tVQRW1eT4gSYTcA5Us9kYu1WbCBY797oY8x9hTDU2na8sqBspvm4k3A7ZQwS+J6T
E3IhzZvHg0UYBDq/Mbd2Wv/EES/N0wC+f13hufEmvHFibsHiaqTneJPeXgMMOXPn
EK5Sxyh1+4fbAEDDcjw7L9sHCXJxOiWEdbhKnDrmanMUbTCpDLljpoSFn8eXqkqW
cMXQLyWf7tCRYDNZCcCEcgGSv8Oj3kK+0vf36yqMH2t6Tyc2JI+XrQ4MNP13oYfI
9ZzPkn8ot+RNeK6twPqWjlPP/MwxbktofWn/lEoyGeAtYa7bAmnaCK37vyyj/8dr
44ZMV/PzC9mb7rT4wny8AeH/qyFp+QOMumeUG/aVnQVPHHxPiHoDcqHHr3CCcQs1
IBFuCsJTklEca5bvda6JBUGqpfzlMac1qWRnYff4NnCaMt38fJU307HSLC6Vt+yv
OMiTqxB8vUWPqVXZkUw+1mT3qX3kdsPViQwlAbvACOf+y9YRDKZMC1NDI+haopSW
3tgLoto0Ye1/qkwFFtJaX/N+jkIgOeUQhSrxgtnv30PSNvglOTR9YY43L1xrCT6o
OK4pQf1rlPuKK3N4muhD4+e+fTNePeiIwM1LZqMdtS0PRPhi+Bw2vdR9Q2Y+dOoC
F4syoeB+3VjdKI4HWl+6FCmnheU5iqA4NfwEdzS5eWmAC5Lo5mD7cIx6B1z7iwYq
kGNcIEnPMmyTSVNvAYSyHbWPQgSmWBRuf5BU4NWwwG77Pm7l3e5PJI+d6tobQ2Ff
bw9F8x6g054D0GTFGS94sYp8c62l6It+Hc+Kqt1izFEfDgxqsEEEskGzb+H33oms
M1p76hutc3bu07NrjWABtprToUL7ldxAPpOszM5tT7yELbt82BbDQC+pvQb7TQsh
1jq/G3qzvAHiAD6qQLRb8fescWv5bZTSjWQbqZxHgOC4iLqGQk2ojaByq7Dj8ICI
PfYiZcEEGFQyF1HEhcfnapbv+cP9lQoo2lqIgqfO0ZtraDvT/8j3fNsgHLY+z+KH
Qp1JZq4VRtwKmiLLMEACruoEphtSu73dwGywJRZD1R006LBGsjxCBFHtJbI1U11K
N0qBCtB5/lZ/hbIUYyHyu83mRjdVq9XWnPpqxlMKUjbBj+EC+oBHy65WFa6c1al4
YjiRkrAfV3i86WCxWg6MIDU/pDryn2jxqwM2ZOTbVzC1crWkCwIDlm7ma7bZJyFM
UF4ZOXw6HRzTJL5FOahBlrteZsJdk8SE0klQ2r5H6Hsa4VUzb8IggfrPqF2Z5wkH
qHqrOU65ZhnZQYw5vdan96SKwzP/2A6qZGafvCg1WSa6Tu+rUs+6Y7wQt10JyGDP
EcL7OBmiUdRWEznEMYzoSuEpX3SE36BWk88b8bUGnc/B1FZdsfdKul8vfpkx2v02
8QJrhnuZrMbQh7m3jNSgTveLtIngK6oAPd+J3Z67zayuPbsXNWGxya9rqG+hTCcn
nwG5V7wMj/aaB0MjkC1eDT3tE2KVoTZ0Cm+6UGvmESjPG/sbgc0jIByl2adG4MBg
3fIG3qyfxen37VdcjkQ8Z6IehlHQxDGp1IcLEOD70mdUaHF21eIyaap+pJoqwE1w
Esa9cHIBDbrVbXkgb4bazn7ccquyWRnUtE1jbXofWkWklXr/kj30IoAKRQfrgqt8
z/XWSKauRLEP13b4B9Jp0gG4F/2dDwDfDLlCIN6XcGgMXVH1W5PnQYubGQuu8NAe
4cccp5b8MpQde1Evk4tq1SjG7xwNouqQ7bbSb5MxVssjnFiVF5SxeSVyNqP7AdZM
IYiIq6BBZ8wQ5s0l4Yd/A4oC9iHRGfKaIzBrqU44Y0hOkL5ofzeVJVo15kuXK1Or
8GWCleYVLVWnuigS9N52BWnKbxXIrHDI0QAsC7pjXLrAt4uvphRPpAdxWk/boYaA
c3L2iwxDHWrpPB3uZtQ2iWFZyxsLQdROgpPNzv13Ks/Wq1EyqD6cAMjvOF8+ZqgA
LYG0QBRF9NyhX1xz1TOiVNgZGqZboSs7gA7m3PzmgBwH6bIHP8/cOll8wrpk/7aB
sKk7zCP1rGhA4vb8YTVLHArpZGRK8cr+ax9kPvk66dCKpMU+ia+VPRu/r93QFnNB
AcYKy3uEgDkALjxRN3Cmgg5Y2/WGC33/iF+Tc6oFeSWRbToLX8nzOpLmPXEmUuWZ
rBumCnelcUMTaE2+Ttbw8KzHzvWb+6XnCBBsE36unxq4p7cPg1sf21+0Q/MYV/q9
YCHUfZN4Uh3noclQNSM30qhpiEKA2wa8TBcRSi8ReWGWTnxAxd6wGr7MzQ0e1rJV
suzOEgto6ZVR2mHfP1nBBq9L4s1s53NgnTcqy+Y7K6ohsjZyuYLJGUDUb9Ijt8Wa
gx/G6xdaOeRBb/aOTW2lU+zs124TzXUBoLwWHceonoG41DlrmL5AMBEu0HjITLnM
eX4eiRhqGhtXBjeOY4pSvZnKyvo7ATvilZ/VAlAMzWwablJ7keTODx++XMoy67P8
3nhXyFQ9a8eG80kkpsFtMWecO/IxGeQVySQ5TA/yFQh0FS6qKojC56WhZfeg6A18
DrxJD1PuW15Qv4T/U5Cwd5a7pHLsJbarLmLNo7wSPf/A6AP7cSJnuqawPr8PkQt2
ZRiV78fa32NgvebVNl0JHU5RlMntcMli7og7AnzWS3vDQi8inRUVrWyjTif/8WQA
haCBq2mExBUlERehOUjegWvAazkdgIC+ZW1x70FPS1Kh1//c6C6MK+5oJfqdQs8J
R61fWp9VDfdRI+jk7INFLiNFsBBr/bCwJx+c8kRewSmOm3bOtr4fWakVaWDJhnIm
96w8VDC0T9VCRJyMptFrGVXh3t923GfIpSNheHGIONU609x9x//znIiugqoMbGtL
ZH0ZhA0E1AnZh/0Yv2laGo1p3s7//+pplmWBcXIKU5SXnWGd5qwyloiLWsqnmqp/
Rkvc+xwWaGHthBBy5pTX+GgzwKK00F7ne88kyseLd7RrYCtYMR6yX2fPYNkWgN16
We0FRSYhMA+UxblzQNC5IaOdYaE7+p6MdwVWS7SniZNpUMYKuxx/c6rwcsTw8lYX
sr1yQzg1PM06BaVewrDebqagIzyGYWx8MeaviaCLYJRF3ITGidzx/4obrufr0mry
PqNRxsqVHYxL8am9P0xDEoYU+Qn4OCkIsrR4US6F75c6ttfjyaxkvcmuY1ArC/S+
z3eQUBR9qLRs+R7oqIL1IzQIpZrFAUjt676AQyAFbAUdhldKXBbR9LLajjyWh8Pm
IKmO7Cj2W/V8m4vxP3gurIvpyslIUObRPMH3Az4ojr7orQbOnhXWY84wQeRO9GiM
yBDhRd9nmR3goS2mqQlZrx+z8ispYzT6kn4NQ3hVuT56btfRzV1Nc8KDHa3gz9Y3
As+rvKIhxXDr//1bgLsW15T3rD3l7f/fC5stXwBpjoBTSspKPD2xPLhTStxHiz/o
q1YjEjASabFBuhqjCNV35P7G4GTqRxrJ2tBKwsbNTYoWgkMUCrYZgGTyTRsrM/CB
oQWccNUXm5Z+K4m5mjbBz33ShBolFg2Hmq+xhp/dB8zAHQvTUmGQs3fogqIvE+gA
4Ue2iEXmGKu15tSAlIwwAbtCn6ZN5lhL+cawyNmlG3jbewt3rTXMF9HTkGNZTCx0
p71IgVGECJXe4kgQEX7JIfBcWiBleukudlvL0ldlCnzkzZts1ygagtUqqL13FYkb
uxAfmHg64SsVi6xEtWNWSKfYpC7q5HZwhSHtMYY66ewuqQo3FFV6b2X9GbQCSQdd
z1RaaIk1AGafczkMPbYCVorYQwq/u3sxwV7baLlIHs10W3qlWt7BKGBRzTWdrZlb
3sSJdkuDEePbyKFH3+2+TsZtTArwKXKiM42pkrPxPMqbQzma1ssxEOnHhq64tB/S
5oHkk/cM5HJ88MRyi3C58eMHGg1L1NkStMHwd3azIjnK/LzrXJE7cZFSj+MpS6Nm
c1sK1nSGjx1HU3dnZ/7r/gpUzn3RGpnflQNfPyPD/0KKdgWFRjlF5pZSZif/MtFk
VcnHfU9EoVNd5QRPH7KMtuynoltbLYYnsQTJV5xBZz6ADDjEFDDwDva6AC4i7z9m
xWt+JSlBrEAJl1CZ+FxP+CqNCrDQema6JK96LyDxwtzIXYfgQkDo8ql0xdFTW3B8
YDJS4Fz+zbZq6vYzCRpVfT0wBJa6GRnAVXTFhyCJFD4G0U16MGN3vLTv5sz47owh
ybyHGqXpqp/FkAPeu3BkVeTVYIkJpuvEZiZwIHeyPvkrNKQZwZ+SFmsHdK86lL0e
14Cll5VXlJ+LHf+/7Aafdihnd2zgenBH8q8Ms1gEQew5CwG9WZ2E4vQ2dl4GN1UI
fiv6XfBDmTaCprw+C5EXUUKPn6e4dZ5/QiqWtq7Y2TFbfLJSILruZDj837NCgF2K
sz3qJancHsYZpfWlbWepalKi4q6UfDOr0X3veY+CUJblmGq3KY6IMZC+u4/EeBq+
CkQ5vS7ductWZhIlk1SceLuTEVcSyCOQDgd9trRphbOIQLGwqb07WS5lXa0IHFVp
f1dbc7HjoQNlxZz55lLXwChlDVbSWmTKFs5jBXVXGOkp90oyt39lYnaT1/+aAjJw
qW4LgkyJDmwqccK9VhL5sobsV3jmwQ0loRKWnYgvXpebP1CCkCDUdEUdUQEhg2Cm
49umxDhL2IOxsrJ3dhOpu7HhD7gjTlBqhJO4YDQc/ENJSNe6OKVfvgKlLE8UW+2w
KzgcEs1M5a+vsd+Zvp1Ng/gYrispOC830aCK0U2vZVVZtaxMEZxdZvdkXc3yq4jT
3CpIcB5vK5vUnl3+tLNxuXPEqEdHw1LvZxPyz5v3q4POLYb94p5oUq4xrBsuQezg
Vq8qiSSAYyHaDRn87UaGCX4hq8Rhq9syRZJKwVCCRXprOHp6MdOb8BAwDZL1LIgX
nW3rwUwnLNanRFuPssEjkUqZfDUo85D0qxBTHq/hgjtR9qL0EDq4EjlnMIjtcWT4
TF1lTiEf2hPxI63bQY70cD4xWwFQ3Hq87KK3Cx3V63ykLIuHKlJBlerVtMHU41hB
F8MPJ+fBSplErcdRzYmiEostg5L5gWdk0xUwAWP5Shy4INI0ogu52RR/N/v1m49f
dsrN91gvT3m+Ugbw7Cma4D7GsCJQlJVI3xMuGfNgZhifdtwwabIJiihYwAVF/eeR
42apiaYmMzfDTlGvXrwGBqfVQL3ZFuefCsbTivDnHCs/WDxdwxdHN2EPMzmYUYd/
6K2xz7sxhQMVk0e4gORrx7rn4fKxRxFRoSZIXvjKKgyC6knwuzswrV99uynBCm2q
HGAEPuNZEzCy1Q6qbov9PgSd3aqE1i3D0Cwm/QwmpDnQyzdYsFH8qLUk/B+bUJrE
WXp/D0E47fhOmF1FnZguPOPhOg6m1axgGFzvD5tptvQqIhpaUzyOmCgCIOiVqwUQ
7poRC1HLcI0wg1nHen3XdqTircSPd1eU0eYOg2G0lAG+RwzlFtTRLBcHL95mzAmS
MjRwTg/J4lzqZ0ZCgMkOVvIkpQXgpg5+WBC1DXzwdep1S5gAi1wjF5b1aKItbwWc
/lxy0XJDw2bW3pTMkB6LMooPEn2eDMUac5eSDe7AQ/8tPrSIxKQUUkr/93h35I24
q2v08RN5Qlkpf6EkOKzQThMT6niY/c+W57f2EY35UAyMMS1+E2ZU5a8+b34vms3Q
SG9lHs2pB1YN9uanYra5M8B883lW9NMWrX2GxXTsqL1VpS5pBUAL5USZAB8reo06
ijnXQ7+3NbXfKKMR9ultWFTVHpg/PiLv9V7vxN9V6wooBo4DnbN0Wxmlo/DMzOPd
wVDpJuxFuRMLmEeVFtZ7ejZShgb/W/h0rt4yCv675VYddkeUAxGcqIqWuJm/J7Zl
xxwkKv0nhxeN7Z+vYvCU6phvJzd/HA1crLWcBDp8AsgBcebWaFE1flxZrVWO83pH
hcZKHPn6l68Q1bcio+UsLlHlOABoMw6/BIC5AdiCxuC3mw1J+ovwgMdnQODy7Bi2
JXT3GvtZI4n0Jd0MaSn5Gbvoq4rI4XT1jBWvv5k6E4jiu3ncroY3wBMbeeaKkLAY
JoIqWCcYHtIgu1v2XImMv1bPZdyTb8PmvlWVLTXOm/42RS1/vxIfM3RlZyUxpAbQ
9I3WDhd1OmBBwRTTeVKk1jTdEnSxdjiPYo2WSm4HtZOlqUJ6cON7LujwoSu5Hc0z
AeI6OP64+AfXWS9ysyScvFYolmHmWQYaYS+3Uw55jyel3Mk5Wlh+eH/yaOmx+GmF
MNbRQl+HSALlaKBf5ASlAVEsq4J/v4+hgOHkmSb1k7JxtflXxxv4IZtRFOQW1xfz
DuMnN1xwsb4D2eIZpr+NcPFghRafCdJht7FR/dZtpjiognnd0bLFRSm5zaoMu/cE
d+GZwB1oO6YuRRWlVPXU74yT2VOqOYM5BzOlYtsD6PgEBNqHqQQCzZV8Sb1PKbRa
q6pZG5jpft8uNurW7UsOswHww8wqmdictdU5Y1LHvMrd8YA8KGxjmb0C9djkE6Rx
1dR3qgzUfxUyQGD0FI42ZMlXtWdeBCETq0OVNam66ruLWyoYp6Q6425IqkIjy9c/
272wh45PswHm+41sB6/8GwFA7l0g5h8VXKwIhk52WBrTmwLrvPdkTcFPqqo1Dw3p
1dt6mUwz0kDxzHmw2e31w9IDfXxXhfbOQx7RhJ57KYszCbyyGRXMw37pTzaLFA/t
+dRHWllAvlNsdsG/Mv8CColQ2RpJjP6UJfVNCYMh7TmNGi89nHqf/opIXvmXZksx
J3NkKQEOFbUbXkhyyZtWt3WtXV2xq2NVb1Bry9ngh9pRSjMTynh55E45owVmf2So
anLwRH66HbqiEX/8+g6Jbl2w/XlfRDGpqZCB3CIImhkaHO2Ib2efHWAdk+W3odsD
0COFVz268H2ENezs2cz6bw463LeNXCJaM/uZ2aDBxIUBM7S6KX7Odi64qwQwz775
x1ekdeTOPAT+YEI7BvixxGXANrWqtZs8eEbflbq9a8navcAKGR7FGmUhU+lCLwCH
k5zSSMz6gvxy+k6SOB98g5C5IndX9n6mpEsrHTCK3jU9spcE6a4jWT95K3ZV5pm5
YfTqUDWxb92ZlaDn8KlmCt8NJwBZugRq4RZlUqyn5C/Lm1Zof6sgbk4PNcSPz29b
dtE+mZD2BnrZWPHMGE6cJHPzXdT5UTQFNItRAY4+MPGOyIHUg+MYGDpzQC1Vu/Pb
g6ckNdCy6pMycKrMQRbXSPLDe5SKEq1StitE7SxgKz+CopqCD+fGtRw2Le8TmCao
dc0iqvj6vnJqqZX8Wkx5uD/+0aJojeRHbbS9/E5G6qT0T0uNV0T2z58E9v5kAYHA
U99x222iQtaETMbdZg9hUABzI6EBJKKgEj8NMMA8SPWHIG6Kv4AdqVr4ymH8vyFO
u8ShoGioD12Phe+j/1Zz1qR7RR7lo9m4fb6ZkFTR7oC0GucmW2rZh6a09rhHOpmk
jcv/P1i3xh+vWB/kBWsfGY6q1HUBwJFjLCqBGBLIBwQgVpsmtg39sF43P8144Atu
i4AxZwUqUCkJzqKbo1rPsZET9SUckbfQRaFLUJv1f5QLE8CNl07kXQ9C57EScmz2
Umt7ro/TjVAK9sPI7fDfRcPSSTvzrQGrm+vOyAim9/0XG/Be/KVLKXzIsbeSmULu
rK1y3GNLjh+ElzdnDVgxSm/igiJlK2uHJloNnGREKzQapIBHNb4roxg+o82LCTHj
37Ks346FSn1HBWu04glinJpNUL9g4HlicJ5nGqB5zV0dNxp3ygLmxwnY7b6SK1P2
ZtIc/xN6XvPxj4TiBwfo9dKBQqBH9sYKyw1SN40Ij1eUMLq8GhzRJVDyHfM2I6Vf
9b+IHEkhlR/QfDXgT0+2Xr1gXY02Ypw19t5cu1879rhLIB52KKmduWb1UFahY+zj
wlFgc9SXowTTYk5Gtv47Q4Rn3Kl2ZSTk7eOSB8mFxlL1OfxgwY82HLV5nYwaU/k2
Ffc5KhH28PrhORnBb8FmB91v9vRIjtWrRVaNi2Naerp50hOfRKjrYVz80SmEgaVV
B7vuMfb2tmhhLzLDkAU0lB/VOPMjrxOuAemiONF5pfrDmPc4b3Pk4yE4xZxfq0/u
bxAd9wFEyVOLNgoFPtUPTmmTe+ig+T5kFaHeYhS61apFlCAZeuabWvAr+mS6qwUw
UNR2fogxWOvydJiRN1RnsY/zWjT5ae2BlfI9gWkPRTj5SlY+QANKLeVJ9wIlhc7t
AXEDauaE1m4oXBnfStzokWMSiZvMl+ullN2CvwnvMC0Q5xm/Km2891ftctzcH0Lu
4wJ+ZRN6QpLre6RXam0O2nXld3BAovBqjXSnkuWm8edotfsQ6Pm4yITwB2rq4xwS
8rDevGdhcCKZv2XNZjxis3rWSQyYOuzUNG2QzndypzuoPN6Op/AwezT3Nizh9GeC
V7b9cUqy7OF0iG32Xden4KXjOv9E5EdrOjXGS4oJ8UThGrKTfF931JNVQwmgROUL
zGilBL4YbuuKC9w3dli+CYF4GMz2dsahlpzb7xMdRwkXC3dPnQhYkOFfFZwDsBCg
Kcqod2dd8MRXXNJ/vId/Q0Yp8B8VSWA7K+bNlYc/wGYfqdr+69/ufslukJhjESG9
no236+gD/9U0GraujaMOK9yE4A0oH5jIxeNYAi6NG3irZzorQK4YVsUPYq4QMp7P
xBMRwDjgENVwaGMk3DIV3nQAWgSWJZHYbVCqkv3q7uVvCU5JfGG8+Ci0yODO404x
puNoOvbeY0CQZRYjHUbAfLjwgIGrx77vunj0sqdNToB63UTi/BX3Rp+4XMHFjL0J
i+Za22ra8hJkL+eNtXT68yDeWqJpEkv0BYUuMpSA81QE70oY6icH1aDWUcFUXIS8
ML84Qn7x4MA4Vv7qxRChtieNOemLvjM1jz15euL/AInZu/AOxY+4/9fjmqmzFyYn
dRXOsW8/VQ61XpVrlH6PvQgSiIDQIa15JG/VBgeA+L+Qdf/PlltzuOjKQHJCcN7/
BcWd50HgsttPLpSfIkyz+lPBiTm0Hw4mRWFgl19WHdiKK7EBfaCRJt1we92c5sMg
5QIBpJ1m9deO9uSjh+YKzQjJ7gfmQTtvgbkyLFf5bHIsf5vlRlt2txRvITkYT4Is
nw5sATfdfuNA8jdhyI1n7fKZjbS3Y9n4+tn7o2+NAnungCyIKzv0cBV3PvWWRVZc
csQXjhl/lXYqQFhmxctTQos/0gqEPM2+K7M+yaDwsHmwn/KhaE+szsWYqwvLBqP2
1KjwNgm8wEVR1L7WkLMgfOgveCgEO2KFcT71g4VRxisLATsKhwoVnjXAn2Zy71vg
mDhSEl6jWYwXlbs6PD9ju5HHYHfs8RLrVP/Mc1CWeLpkMwNkcBCsW2i23JCwZXT+
y8SrHZOKf3O1ipNvqG8zl995344S8nygY6xTtxCUc4Msdj+s04ytKHCAE/O9nvMc
fuHySx5mTxU69jacFmAZ+eDUBor0ALWrXn42N8hUs6YNu5WEwrpZux89NLfnzBmX
QfMCf9QPmzisPMENPfDnrIKcAg6Mx6DIRTaJwqqjyidGsxuT4poD8gIDGdsaL3yI
9p7TblQ8uSn4vxZkJRQ1Cv0HMkuxaoPA7aoOVCZ8p9WPmB4vhUA7etkalqljwird
cG0YmPYJLCSHtnKF/19TOuAN5N2fPEzzZ4d0ebrkQuDHK5nl8GIRjIMVypQTx+qn
1S1rMYiCf0dlMWTbUXAfYr7rQsCXkrklHGWoYnXGjSpgi87SV59nHTO3Zggx4AHN
SnluZdoiC2b+Of+bBZNFFccd82SUP10lb/IzMqPRt4sgca5gDcfSuWNoEZuYOPtk
HU+uMb66acb4Utftj/AQEMhF++yKOMD31PW+40eMiAiuOFp62UH3cel+/sa8ogBI
5jhox5mPshhinWvgMDJKDchiM3P2JiCNpeKFJ2zengMQipDBK6VB8v9B/2k2PZM7
n0KZ5OoUrTOtLih4bZgLLXmRzibQgoUeYuWZGpBP0soKE7JYAVA5s57j5gCMRQlw
OvYWn0/BokoVQxLifL4CpIRSHzvcpNJvyFML6u5EuOJ+XAc6zv5sz8zMXXqvFoYQ
zvVC2+Tcl7RInTuu1URnFnxBoPBOnlaTkdP2BDLP9jMV/OcbfzTkIkH5piuphe8m
Ii8FAk5mSSwTMeF9foX9cru5zBDPM2gSxnSR0xLqNv9Sx0/uIVa8XgiP6iHi/60a
LVKpxhY2Ng6tCmOnCIQLrsJrWYTYY2D8Z1MxtjYZWQwLG5EvRnxE6O9YrpcOgMOs
aD9URNDMxHClRq3xsN3Ix+QSJ+mh37Edmc65uqBFEqO66HreyfdBDNoRls7vR4or
lx/LDDVztBZfBQGCYOv6y8IlGOOk90vvp3gsLN7EkTKlgCYISKQ6Ju1uCRC/knOD
3099SPr9uH2jGkH0/4aTrQ7V9mYKMNKcEG7/vHJIqFRkVDPHZ11U7yZFFZGO5JVV
cJgD+HtSJues81ruZi+MsyFf+1ziLzjPZB/oKTHV0a/T9M6axSm4mu8YMMBGhW4V
5QJBhJpqURyStHgQvEsAHTZhGHnTGZz1CiOwtN2x7fZUFKKyq6FsBu+6R/ltaI9s
/CNVgoEgTHGL1Dsc7jy73julaRuDfVFpaXj7mvN5iB2njtpEOK9oUts3KwZVvMlD
CmZvtX8QGdCD/xsDDvPGhysF6YhKI/wd+UuupDuJgo/Eb6ANw5bw3EB7NHDOPG40
nlnzQWUtJuIqAgjD27LnVK/O4ag0lmInkWcrrXyETa70JrjeT2M053F9XeMvc5gF
RJ2ewSQIRQ2kA/TbRYxV8Bibz6cepIbHdxbjd9BKWjIEOQk9gdNNsXxgHZgnWVl8
nxWLrspFZ7HX/KSrpk2hne/ph9qyUe+ENBqA32sIDSEqQwFw36PIU77jB4npQ1PQ
JQG8wUfgBHR0hADKQ8KalOH3EOC/Ok0nApyi0yeH8Jjvy6+zt+vF6ZpVyLDj0jbP
do2fUNzPHah3DoD+/SsGKTAai+OxmJuhJPikAoyxiTg9MdVsTSgoi+lYZxxdC0DV
l7ummqs2wfF0manh8qsQLz+p/jP7t3VoS5kFS7rk08LOYqFsnmFFtAhnyTr5Bx1d
kOeP2bDHf6Yo4c2UtcnzBEbJIo9INaRPEQTUx2pXvxoxAZ3j5ZcN0GySegn/cJLm
BDb7dDwUaTGjExGXcQ6tDXo+qqDXtMC40O3vXsoN7UFRDZWY/Kn5PGllFQHQwzhu
jlrBBv9KvqTjjFhAroANS+sZWUHfMMX0w98zxUzwRy9JXDktpst0uGgnqcacPkuF
QhZf9eYBLLUyXaeioEo8KtlDwaf3wsTXW337ef79EdUhbgmiVieypSDsMj6SKlcY
MFrXyUjdc5ac9x0I/2+Y+0JnA8qA+QZYbK0zJK9BN0qPHj+wMB1vK++GgZ0AjRTp
efaUjBjHWcB4PqS14y0Xv2ETudR2/9iEaJc6REYCuNf5QdzdPxHhiGQyjRo9xoBr
jcNAbK2u2tBycGkMbsSUu4U8zcNjzvCysa5hP3cHGx/qAKdVgLD4CzAmN3s96vZt
cBiXwHVP4sYPwAf0oPqlhjCorOc+BaC43esIsqekIFHjnMt5Rncc+Uv+lIgY2tv1
UurZCanybifUFHrZAwLND2rKgaEf1ZyU825kpq8bQCETMWi8ZUFH7AwLOLqdjOpT
9I1uQ9AFkwmoIYr0vtK8ZIcpNZl52ABDbZVMm1UGPl94us4AtFEhnRHFgwgMR0Xp
H5CPo+Zyx67LTNcaoEVIBWxAQzbWj6EiMMANrEJ+Nm0MaD7Jugt2frlupG6f/5/X
FYH4rev8NJKj7LYlSeYlk6+3wDrna7xBToXaXyqtWxw4bWxWzAj7WTcfJdvXXeRk
DWp4KZ8xjywf0fFVPTw0V22eDRDwJ6vzc9FCLx+ghe3S5nF0O2DvV8nO1/nR5kDF
HlaW/uPXAMcXInqXmVdyxAg0I06Xs/X7hwUMFpMCKpaBYVrHxTZDt5JcJcy4c5I+
2s9evjvht7SQh4eYL51R51E6/TwY0z8eiA7Go86Jl4boORl86GnOTKI2glNeDohB
niuRlGVzt+Gk7VGrWe8nPE+o+IF3vqi6DQOMf5rNStZoCjRrIfZjk6NnAFz1Ijac
bE/8p9I9wnAltiNMrIWgDjtpSLg7y0Ni1kDmhyb91jwUgDHj2QFB82amwErgTaCD
wNJPiJOJ5cCJgiMELOQwCuCGXDbaL1BU9EjvrwL144EpfiZ4EVHAQy9yvLDhe39s
B+tv6hX/PCM/rIUvmYd7IkQnd2Mx6wbHWCihAiFnNKFZbhk7KTR4YWQ6x+w8nGwk
I6Zr6KqORsr3IWZEKO7YUhJVzHcxWg3h3F6wDQHFKfvw0ojHY+0xeLSymSx4VL36
Z9e6Z8LmdEBJboLm45ahyMSEIljsbs2PzOQhnmHzFKa1A3UXLSa1nRqNCE/91PSC
2yQA+Hlby6b1NWg8sOsx6JG12MAYyklgMTxTmIKHLnwliiEos9YF7QCemUtW3AOH
tkG7FBl9FFPt1aU+xy3VzMlnL4gR6PASmQlXkIjziUR7GWRkntfp4zMv8QXw5CaP
MKD3dieGuMl1vU7tWZzP1Ckby2ubOrEaYw7dVJ3rQbPULhTkiMsTfS99stz8hlJS
IRcz3yYKRQywyILp1fX1JhAjqPc5d9Q9ht81YO0zHE3nA2RCDcFBShm2CUiFoLj8
9JV4XhAVG7hWZfb6Qf9VlnXCW4gJZFPzwDU97MonW6pptt65orn+hxDsE37wciMG
/eROCYGRd9BFYWWMK/jbD2OZZREM1Y8MewxjQXXxZSyMFbVSoJF3jw18jkucgSyK
e7EC88vjPCzr8GGl6a5GIHyVIolgqLogm/UoCMmSIjY648yWD82TWB8NXeG5JMMu
4OktLxz0vHWVXpNt97VxX56hqtXzLT3df9P10DWc3J4mKom+w9YHTG2k0xYmPBrj
W+YoiTDLgG4gV9a2qInc32BVi6aPxGnNXUzaQAeZYvheABgLZjeYx0Q9DHYWZwvM
hqu1FsjbSz7Rz6kcnBiAq/38cXlLVVNxP1Z5/0Qo3McbzJQ0PdvMAXlMV9iunF/H
2rIAj3d8fuv2ytaQemc0y4g4qsdV+lAsZXddUmGElBSKqAShNKgPuQdteDVi+Rcm
qPKEAwysSawJQv8JQSS3Qhhf27TCU1StAW2QQda25VGA9OFUI5+u4OKyLxHyikwc
l9DTqc4p4OEJ4Dv1b2NtudsZ68BVv1NQRTNsEc83xye9ur4KcH77JitZl3YYqKEn
0TSLBrkg56M9eCBvonwsaKHdIOhIrnzPkxy4AjeQQ4uPSM59asc51M5ta2DZsWJ/
40pPteTvuhLY9yqLJMWK/0BW9wR0Z6o+Z363PU5e7GFd0l8b6GxsVaSqKbFK1aRh
M44bGXqR73L9sOL6/6IRJriHuFJnNGSCDkIRMayd2dU6S1XUO1xONaxx6GUq+6M/
lsjabZL0x26jpZ6ejQLh0pv8OqoKgtMTdMsg9flUeXw8WOZIZxUpSPOrZyb1zuRC
FsfXo3zlvLBqljj/kLFh5ejlE4zReNA4aYd45rfpI/HZ47HeCt+e6qDcQhiJnNIB
VnyA73G7bTXLbCS7cqPCvfejdlyGNanGJFJ0niJ1zwsFahfq4o5foFTu7mmotit9
zPAF/vODfPBJKvIviC7ggMf+Snx4A1CYQm7nlgwd0S8Nm55XXjcqg+zgy8h+2Frk
+dRsQzPjUZ6E0Faa5rPBIryF0L9HK7b7Vb2bdrnqSuDEwDxvPoqk5/Fp5swFYc3N
fuDfCvaeaUqGej0LIYNwh49Ab4JWsSvE98GGKLvzv7DoznQsDixDug+u2jsUqEjM
8JDM5OmDVkAt4T/upANvJO9CaW/14HiOEahBg+7bC/tcy6SeUbl+SvUbVKehb8l6
I+q0eY4ks87Y0oYFBjPXOcoGXfQ+QTz3WIwuMtYpWvKYEu467uFfKhiPohEviQxj
bGUKjJ6DyX6wn2r4aEJfNhb7y53vWZiboIzk9xy6bhfGhSaryTLCE2EoDHxYEGaP
goNB+zn1iB7E6kZQHbRsObPTkFlcoX1a+OB7cvlBtUL9a9w2G6W75YpvHb9e/bBm
nb8ak3TOEUOclG59Hhd1LB5lY/MRzrTYe7nKPhhT0AQLM/7EGldmbonVzZy9AiC/
TvUtp1uI1chweAaFWY1n9Lh9cxXWUp6coCxAmRCSysgO7gaHT+QjDRKw+u24pmFI
zloBOATm8u5yoTHn5cgOiB/MPZq7mLmhBzLsUHj3cQsAfANJCMiZa+PUZHAJZF7f
Jk2zURY2jtcRbbU7B+S5eyOmzN94Lbilw3OXb5u2zu7uoVemCIQbIa5lM6YBuhzU
ixt5+I/E+mlP7m/2srs+UrpFgdVftQowhq9lB+lHMtU6gGsGSEkVkafUq3AFkmVL
SH6b6Oujs0J2P5LZDspkZaqEQG9TKUH2bSgxlY00CBGrayfPxWqNZyvB5kXNM2IV
J01/pm/lo02PCwTxDAiD+cwFW7QU2+oeWFoXB6Qt1GkP3qGZ6AOLu8nk6jZ1o9Xl
hlhszo1R1vxIicDmUfYhwQ==
`pragma protect end_protected
