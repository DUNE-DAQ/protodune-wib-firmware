// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tiviKaAzWucP5YZvPRY4e8pR84UC30WXh4ueGNC1QRKpPnVocUJed1KuRMBa/n79
Fe3en9L3arBak1t/K8WoQWMQchTNhMKyAtIEYoDbzJ77xtzcvMG918j3kLO/Bq+N
lsCjJAbPxCoIEzKuRIrEbYf0k0fa3qZBx5RjBJA4WQQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10768)
hSwh0vbPEazvi6j/M60jVx/oCPsrpdCK7+3G7HvPuigv2OWzysKqDg81SmaHCOwL
proqw+xdQ2WXzss5i14pNCAiUarms0ny3vzD6n006+/KsUXpq7Xdkquo32RA2Dkt
l1W6HMQMy8VtUIBD/miIpvaG6jqrMpExgGHldrqOHp+osekKmMVhpu/LrbFTSbDn
pKHoTggmYGPB92kziKVVpsGM5KJ+KgQ3e3gmfDCr5QI0jiqMIja0HzXMyxYBgN/1
VcdmFR3RifX0mpRPw2QAcyhpVdugr8yvNF41YOEw1wCRmvFjZdG36reAhArT++V1
70SfQ/5hV65dZLo3wLC9E+Gp4SZGlsWkUBIovSzjwqe12y0BY3YhJuGO+pTV9GyG
LcYCp5H+swV7dtfGAnwrZgr4KH3LdTUW5IblKXj6R1RoAMSqZx/O30POfZAeT/sa
EUTTqVhwiRuFHBo1PWoBRjk5pfwOrs+f4J1SWfxRTcJ0offP1uv4119hCzNtYQ23
3kjToibLJkiQqsd1l4KL5vWplkiOW9hGFq7zIzHjI6QvNH/u9c+Nllx3fQOvkzBm
lrHKfFqH/oqsY1QljIypIQFHYJbQIZ3+ve5G65nZIs/aW8uYf2THy0ShlonfFgMr
5DeZOhOxZqBnmNofVqTT9KE5UYXlwdxVID9JVKB+htI4QCq3KtosmNTQsWkbHvVq
xp/eGUgPpxmwsIhneNU6HixZWPwmmaFLky+1CWU432+ABwRNSFKphWGYCsFsMlaj
M+Wig+LecVJzcz7T5S5DZdk1MZmQvFakvlU6ApKZ1sFiBalteZMTx1n9lBqPnF7S
t1O5mwfS3Ypqa1K7vpwtbJTJYCIwpmF7uZqopapcwV5lOna78k0z2JNc4MLCLYK3
Wi89zeN3zJN1jA+4UGszvWpIKIlMTEN2hAYm1a3MjdZyrtSO3RG0f/a+9blMQ/mf
klpJCvashrmfWKDlLTL7PGxi6ZCWjv+1Pzaf8WB6pc1ZVmRXE3aBXkTLGhccrOCZ
uNdDlOIvE5BIGU0FNlA6fKE+9l1bndQIURg0vWX5Dgyl91QHnOImIau/YXI5DISy
cElbCcEu6Se1wJHwhtvZDpnoAg2iUDZsEn0lXHI53iYQB/T6S1ZG5+xsOVj3Xi/1
Lpz0NjaimNJDnBNoVBo/MXt6FtA1xUzW4iCgmWwmdBwh49+lWDftK5VmReph/3Zu
PShZVxQLu8Jad8tLMCAOAH8koWL+hyxRMh5WhdjicPMObiQcg8EQtC0cPIMdlTGb
uJBbk96ppXrPm3w5Qf8jk90yyYfaV5V5fS3Gk3guWevrhngm5d5AgB6WIoZ5k4uA
LF+T9/F5wjup72Z/n2iHxMIpXz0KfjKKaounLICVSdoak9tYZ6f8br5KpmU0P3cN
c1DqOF+fiTnmMsj23Y3d2L8VshhPqzYrMkNl6Q4CKPBxm4zxjG7Ug5WPRI0X3yLy
kjA5LEQvZYSXw+V3X7A15scpSp0Ljqrh2AeckGUjEkeZYskXcwffPP5P//zS8Dvu
YH81UgUi9yQSd8/b/iCXm1KZncJiteUcVsZkV5MjNhR+eHyy11bF/CW1cxy6JjsU
OkbCdU9Rypo0XCJQQzb4wC+iVlY6jVDnoqGK9LWbDNQypopsG/95YqMFwxgbjrjw
Q1bf6Mj/x2nG58jYSDVKZQyQAgRi1j9SzrrJhtpjj4GM6i5lB05B0chX/eLWw0xt
YBhTHSYEroY5T1oMyA4wWBPO9sJZNNk+uu+A104kbT4aiScCUXM2UAxn4/8kiM5y
wo6WDYzBJcCiELv5dy174g64UiAVwNQoOiIIseeUpUkBlLax2f6yZN6dSbZ80Rmm
Vl2yW9LR43qiwuXLzP91QZcy+93/7td/xNJzSYmC3aKPyZ+upyhy2Ng4wOqgzLc2
xLPwHm+fiYONIvJ06A8JKJvyOxUWOabmrCqLT8WVeAd8K766noo50fWaMHxbcE/+
qvzkM/n6rJ0D013wSZpiFeZOBzIVtiuxZJxX3s1agT2ndlhkKxV0bm7Io7xCiSzf
8zSe+q4nmS69d2HJ4NL7UVTyr6rubdX4jlksXl9MYa9wkPOrSVdQtdOuElAITBTI
lzhOIKzbvg1VEkDbjEFfDQdgGQxc2/VOyaU01/i1LIbWN/FO0UZ8HFmECf/+1g75
Tdgv9Z03Oj/VCSoLOaR3yE/5tU2TKbMBzEUVsbN/fwFSYVjhwUvgEDzTsEmhRoiJ
xM5dx/ZG9oGXb2W9mMlW9el8wG5QflzBuJF2+xO7FXhSnmrKruLe8FBVmnpdVS5H
CudYiBs3+7VrcfRdvkMIAkIDA8fgHZJmG1XYmMpP548dpvCMckdXb76zCvQtXLIT
0+3gD02xKRnMXLto09ConAIdipj8yzIW4tz1db1rQUKQ+GHPmgesrXt93ZpxWyjs
LIW1R1/hfR7HdZnc14V2gdxg4QSNcB99d3Ti4WnHIEcpoAt+4k71PILIR4djgTyt
9uoq5p9EyGSb25BpCvi38VDUDd4T3K1xl5R9RVlk6fIxJgQ9se1skpOHMaBNJxUb
/mG+kx6wmyKXUUODbIjjrnbZdvPaOpajP9IOl5jRWHjSkK80GInV/+XcYlRwkiDH
BSd6nbEo9IXAa13TL1mVJ8RJe2GG0EKXnv8chSIg2qFuDbDjh0PwMgEUcDk822xN
nItL2xrLcIWohhyRwFpb3nsX56YhNuD5JL0p/E2flBAg6/VFjCCveZS9I7lySNE0
pDvG1uRW1DPoR13c+fNjOrYco39k9nzbVbib/JNyp5INCSk/OB9fRgoVQ8mrsvgm
ltshaBhIbjojxmU718zbX+9hK9/8UQ/1dO1oGbPE/03HVIdT4CMNDXLjjsAEUHva
ISwmUAG7jnysFS457MEKOmi+6PcGVpCy1yGYIittVfDth5mpcrxpPzwGdMoxP3nY
Ne5OT+NpKrkXsi9C4UGaMZodJqj9vp4eskiQWA2jphnhMnYco49AuMRKBMMO8FoI
X467+f+NLwUMohaEkKM73/nmssQdN9XsUsBJCgponMj8/98uwXFco2xWDhYMd2Yx
ha3j7gSJ0AtmcpzQ5s8y/pxONFNEKI2/4nbRXYbwEw//Yi+06ypzaTpwdyLhcP3+
8BNwBm8+FeWYeUk3g0ErRFvx7RhhVKX+SuaUR+7IL2RuXEODkXWAvd1RMmR2sfwl
ahEFt2XVRl+FzgxkrliVLUZZg1lnt1xSgFYwviGLKk0skXqFRx1eSX5oSV1qbDja
6WKR2OURfGcZ5pKYmHaB83tPJ68ItihUIm6PJH/UNY173aROBj6qK3VUWV/uwHzf
yyXT3wCuKe86Spez7JAQSlgBpBscPaL7G8TGb6a2fpc6GwkLbRknCap5oO4DBqfn
pCTmcJvAsQIDCnfoXHWfJOZ4MeEzIiwIHT5BNEVsiX/Sli4bRDgVB1kZ9KbEnE0f
MiEl5V+HrVVlhs2zgF3q66xOs+HyvKyQYcAnS+dAdezMldUlSBSbbQipMB6IvNCF
MBYoyjt2cXE/dCoHPtZvd8bucNY/IqDhgnwGZyGCeNDoIKoQgRYuPJAx4rY0YRzm
6kmFE7S/V8P85SLP7J/fFp8/iSXrwwAPLgWxvFN2jprwg9q6lUmTkP0x2ZNGBq2G
XY2g/d1Muc6WHDQyVZnpudP/0Vl4qsbhJ6qDUDRqYzAtowcJiXFNyq6u4WZKEgwE
yYpaV58VUWeoPC6TSMA0XenPnSW8T8fl7H3gAtDdZDa7WyZ4Sr8J1VkUFOf+fylJ
o47b/mvI9N2EmBZOmZNSuxt8mcLFytAYdATQC4fKwFUDFlbAD5IaL7KhO4hFaqqg
uMqD4PRCewbfGANHWWq2acBo7x749dqfUOCG5PewKF0A2qx+xxecA8Agx6zvSGtR
cCnu5hSjhC0WDfUVhoTshk3jBDmtbKo8xCYdp7WWVTdu7JKAL4obGZUmuNra9KMG
ukZp3d9VXjkTEAbPWywYJkfZYh6nlwFDDPCf89cUd0mFLxz2Cr+E+3ocudjA13Fi
oc1QQN7FHCDfcCbgHytXUUgVdGwakRwb3V/EILifIlTE2J1JI47ghYiQAE/nfhEg
RHD8umme3SWxF0S1hHyUI+5Luy2aI8HXVHAoRdY6RfeRR1WwkWUq6c9HMOCzuu50
vmCHAUtOLBaPhYECCisArh1NgarKFb8x5bDRXs91Mn1IICh1qHKrs0DcHedeAA34
T4wHMqYrMvElzVg3PeRpL4a+6iHTgyhQ6eyCwlsyJe3L9jKo6ji/2XXyEBisXXwx
Z7HOyPTx0FrMYd6JBFWfAU24YvgVGTnAFyOJg6WDhRMpbE58nz9uVBLIIczPMo/R
Co49scnNhCUaHKpQMc/FUI/WLwYHURLqwKpELJv/uKJjlP/1DaJMz1g+O6+YCT/+
A3kY4pPuun4j+KLkrGsnq6MwWgDH6BU+Xo+yyl6xr5y/xspF1/oai2etdGsA/I/C
XfuZu/JqsXhKAtkazfC7Bf8N72zzNjV9/rXCNdP2j7NmEeiFmGPOT2uTS/cCMRCW
xs7PNwqm7PYEGe8AfVAGwxa0yb1ltNqG7ymgjiknys+ub+JZ+dxUBPz53V7NgNS9
SpUjzmuVw4gGQhg03mmn79q65mTvs+98uCYGT06mv+eLWSCgPg400XwsfqNKXdIz
ThmCMYEPJ0V+WbTL0h4veqyFcTnBoA5E36cdJMS8jD3MqBznshfL+WgvDcubPTXf
0cVcPzTDqhP9M5vxgqewnAi0LP0zIfRf7rjQE9hskO6KJ7Rlt2s5Yd6TQA8tbF7x
4xh8fM5xHASFNLdF9Ih0Uu2gPKqaLL57amYU2Z0slTDUUkKpZclTe2aTQXoIe52g
mWk+vdNY8LJCVj/Xm/f95RN2G7SpvyoBBPrdcaWl+Puvt2EQrlUPU/2Xws5AT8Le
zddTuwTzqHqRNJhTBq9c1pt5sPjHtmdAwxh023gJsESQRVsqN9RVVyjd/tP5ngUP
kEJXzgk7ZOhNJw7INZMeTv0L2wYlyM5vagvdK6VRc5Qbio4SGHwKbIFJOvHucGzF
ZdvI/A45omsqo0FWtbIai4aWRJcNtVEvHUe1wvb8MCS2bl8wCLr93bj9aN2d7eqY
VwhHKPt+k2seSgdaQ99U0/fHEKy5K8mLQm47MUNOz9ltRZu69jU3Vzx4Cw8FF2nA
kg0HCHNXt+XIdMMwgDaxEg6DWOnYfTl/5gFGm3DJ/kvi+oM8YnzWjhQDGK8SH89D
dFvScjpHtdL292Gh2T88upgns2a1nmaNtX0hgtxxaCRaiVaXwt0Zseac3ghsYKSy
z9BxsD7AmZDYbTi4aToraZUFN/RQvygViJ9M6YKREGliNPv++FmXxLSq5X4mwc4m
zcDGKqHA4m3vFLfkoNze2OQ1om4xSCwc3u2hVqDWkvGbLgO3wPJA01hpRwyit9gC
5LbXFryiFhfUmA8zvcHGiBGe7j+dkWihfCIatIwZ80nVtyoSIcN34JagGGHSSWJL
9DNSRo6k0F9w9g+cwASIm2vswGfqzmbBZfXVpHHd1JJ53n1ob44f6Qo3ttpdEl2p
9HIxhpdfq9S3Z5eIVawn36dpUnvmXEo4x3L9hDR11hqj55HGLP8cHx6YR50pw5pQ
AdvSc5uubx9w/AUbzpcwIuQIBUjXc+MioFLEQfuVEPSfy5E6pUsOM2gHBn+FzBAe
FYnTRrushmTu/EiaCRyiTNtEHcBCDXaBsMzK6D88jZR8MPElUESCFB2Oe1qaQDt3
9Lj8o1aUhuxJwGJOUe9cNi28xh+XdMGLAfqlCcXkxLuxdc6eVPXAdMOxGhkFCiHl
/Et9WJCmdV/qn9HU7uknNZIWGmoTYdW/dUDkFulWMWgyRmfzPAP3eE/lv1C/naKJ
FXKGHKeWGsHEG+TtixZM9DP1hrF5KGidEsuBwWJWyVr4z/pPNxdjjz8SoPIU2VGS
GOpU1xo2yaxr2Qb4p5K+gLzQTAruMqsVGT2CWLzBH5CpMs8BmcSENwFUYbZWfCG9
xP70m7M4Qk8z8KRT/vHN5oi+SnDYfFjm9QPxFXUhvWxCDNf4CsZK+qMgAfaxm4G+
kCYk7bEQjSlfSue5xoWgW5VbgGqPvoqtFVaintCZrW4phpMCt3m3zwu5qJyLB6FG
dm2fgAcDwxZuZEFlicjpeym1Rxhv2QiEepa/raaGwzXC4UD+2aOOUqgCoshjgq63
EErYhi0SfYpx3/ectuM+/2JHnNlF0E/4yoYQEOxK7TjhygrbAAqROiJvAzDp3spy
EhphTUviNKWb6eCDykxZuoqT9MVKCUyw5Sjm5mZNZJRVdl4Pi5+ED2yokVwmOfsE
I9p41ZR8RQFj9zJXGCrYuRHeR+WoPljkBD/3yMKNL6DGETNQsD8rGFgTOe2JNTmf
FL+aoKOZAJcGmi0bJIeQ8xwMslPkmap3o0A79z/ifq8zLNBQ+uB7GCTiiiFyUPcS
E6rMUctkIDA4k2MlJcX1HW9b7WTuiVhGxRTRG5QDuktBJQaojU9uz1l9suGi130j
1VIWHqHtuF4bh+1nDjYE3V011OYrbGE8UTPOAJNT2Binz07ZTyacclQkSav2ZXOc
EmEB2zVjxHfgVKfOrucODhPGi1D+DnY/S7XtDn0wkE8VPnG4DkTnOnF3UsWXVXoT
qmQ0FsDkbl3WAxEoMLQlNua2KssTf4YCuigF6qPKI5Vbf4lzCU/CgtZ/giqf7paa
vD46v3/rxO91l5lamlIJf3G7PetfIXoVkJlmYJoVSFUq9ZnyjYTNpQ6Z8WutzWVB
TBrgN66hreeatnwkDDOaLoJRC0+rF7mIbFDPza+ZL2/KASTE7mkTX7uE0pOJwmvW
5rxm2FtE5xL9Q2S7O4cg9Dfn+tEWKpQw3RNHjXy0Eqwb1gkVTb6ejQrznb/oEfP6
W82/ZyMLnZRgWhq+Y++W3QjSReMJCMs6qbo91yjlHVLXh7r7rOQHQXhJpiBVffrv
bPXrBVcwsLavEfsWym2JNfXdya8D6vneZGtg1NCQH1Y879sRw8OUJCgdd9/ILPZ5
Ar0Q3bxYXc9hqURFrpdTkL6nnibMIdWMRkMvsnogxKKAbNmNamsIIor5UXiFMSNc
YPypjZicELhbzOouCDihT2z5+7ZVZeDFckWDe26c5sjnIeUVYQZBd83tw61hdGLm
BXO9PeW2SnpDeryCjXsHWMeuaj1s40w5IRmV8l5ODnWykehscgQnA7dArRfS2cR+
rqko4mpP9anYmj8Lutgb0T6AjhuXjCua668dUnNW+iADJd/N66ENKWhbAv+Wd+WT
R/XSWqDBCFwSGpZg5G70ZOokGVW+N8KpRnGVetVitROde9osdv1LGkY/4uaJFlwv
8mfrfOKvXUmcaJ4vmKtsnUmNofTVObuzK5XyqiGpIyMqdSlAS7nN7Ex9wBKopJe1
0SrFGAQfMowIOMhI+ZPDcHNd45YhOUTV99RJnWKDbQdb1ATC+vcsRBNmd9j7Rkzr
IVLiOrpSIstsjHTTha/ELkwj24RJu4uMu4C2cSrJUyrE93VXHwDTCKreUMiU7AgQ
vEAjUS2faeHG2TfNH2HRl0xQfkAXgN0Al/XkJeYc5Nk+aNm8XGY3LoElLGVSH/KR
y7hRPjw62DBY4wj3XtQBs1Cnfzh51wzcA/pBA9lsgn2TMHDNB8UAT08RfWLcydJ7
+nNioP5DLrBHgfTY8uI4hdTQAfZUGfxj//2cKljuHZuTiKZYg3Xq5phx3C9Qs10a
pKnUtvyxUe6J4lv22JjZ5oxGr/33/nOnSyA9BOq/deNhEFw3kW3QQk9/UB0sTx7j
qqXtilRGASQW56/NEKhgK/FfFuen9KLJQvN2zmPw8TNW4H0dGK9MbQv/tqbBSktM
rAXfsRGpjF+XWg2vgsuEWWRkIjR0uinSalSNg3X5Df08GKOIAypesSqKZs8w1liG
t332RklpZaQ4VaHXpcsDSKfgjoQ9btyImz5uFwWv/afONiJxgq8HHeYRPLYxdrBD
qB0M04p0UUwK+BCk37hMiTapwAMy90TGBLZRkoPWcU2QLUer99EvLsSXRYMIZ6F9
uIW5YtpVVEW5/cBtZGTcGbozK2N4av0KVyMZz9AsnqK5eMh8/zROWHeHKbzxZicn
0/oYWfLbLejaKwoX7amcdpc06Kp5jtlAYUQjORwGjcc9LW+9rrK4+RZS7hQEsShC
dBM9EZ0pXL0WKGHC6vQl6OV0zSNSVJqa4UmEEeF7rRAHP3vUa36KhIbdsTUPgr7K
VDLTzAoyJLft1w3wqkxbKxuHPJd9yt0F9tCdcRXoOHX8uPRHf5GSU+adh15+OCsP
L+LOkWjKILqfN9NnYvAqw7Fed9bOM4yPj8BXa+CFgKee3Q7Yc+2z5BpajNjTsGaN
zpRMoHvzA/x/J5/IJcElFodhLYTa8mCRpbSbl6hM5pBaOhFuXr5TeJQ+Bp0YnRSP
k058WXDxPkDOdJFLblQsLxeiqnKbCoqZTN8FHQymUh0baGs6g/SMxo0PWooHbYaL
2Qi9AfK/eUvZ8IqC6DKckFhXGRocdVhjVRzq3wuUgDy7GWVT82rN91dTeTCuCWq4
Pt13F2eIBg6f9LYmvM4NcfxDnO0aRPaaii6QohOCkjxHhEQfDr1JaAWEsGhj76b1
eHGXLhQ5mM09cyHbvHXC74xJn1Z9Xc+y8EVv2Td66/qI6CkDN+JI9e/SkDLh5aLG
9tA+Lu1hduc0gHiMwHiRD0h3OqT0vi+fs8eEmZ9qLebMf7+lj2URSQGxdEHkrf1c
VgBQrBlTJywgMH1YX/pfL7Whu7SuXuLVmYL01iWY4jeJq2pfuHUVuquMniDwIhMs
60P1KsvT4nUUFSymL/eHOJk6qmzOpc7bPsygaHY5opTV6C9qmS98B64dYcuWNsrh
TTXsjM8fr850WRGLbfmKIwvtveNpiiPB4ktubiziAByoqHEVVGa6mwLMjynOjwrA
sfqyjYpakkT7k8+YUNZf4tUfbCJwfVMe2rS6pEDhWhA504IFN2qUI/svJ35I0Ori
BxFMxOSKjU865Cqr72Mp8fMEhCA9qe4BaeMeFbkWwrcFxAPF3/EDCCDYOnA+xjDl
8ocRpr89zwb1uUyLlvh6WgcfNzqg51ff6yH1iZh0GUaXvNQPyr4cGB8cAh+e6/z9
+FcTcmb1UoE9l4PFlDyq6a9k/Cve3z4//te+zMQp4qCb+dfw2r0Q77U6x9cQqIuD
6S/u9d1lQQMqXSO2qUk97c0/HzNRIaBw3B352hj+KW15cQzDYbdu0VFeMBWpZAMB
+hUXpFH9ZpSKPw30wgak2RytlsePMPevd7gNCYQbOzMLHjiEMT7/McLp0DnI1lFG
JVAWgS/BnaZLPxBevBgpIrXRxzD/B3HbrxYOAWMizzWUtOX7NwcD+KRWW75SLCDz
Op+D9TrYz+0oWkoVI/Wp+2EsXAwaH1NkT+VBIaFqHk/NAG+Cx96uVPRlJyD97OHQ
Z65T8R6wTh8eayBGjJtspzZbn5LV7GlHSOY/saSpSpuGJqj5VfUjxPUhpk44RJ8Z
UJ6jY8fS3rg98oFjFBgPtgfVV/xPZZtG8MwKoDCQzLzlWHCXy66g0NH//bhFli2B
UOVBi9If3NsO3JOzj4SMIqiZF6+320zvX7AEDCMRzIA625BE190ZcJqVFaudLnNN
VJjrLAsf4vUghxv6DtTF2LPHCtQ3lBKPU0z1ZW1UhY9pDeEh9XTSXGQkLyobUzdO
l7VSyCpP6WRpb4/zMHaMBE2JxH4V5dSuL4tbTQ6Y6HphWileLU3zT+9LBdrL+2jg
CIDLdufQINuXukWmtnJhIIIDwAZajotBeoXbuEDfp2i64P8FX1q2+PcIzy+34FX7
x9pgQyLeis9I36BArKa02GPybMcDaq85tTu6dobjQRRHQ5tiaC6lqhhH/BijEQcB
tRQE6+l4nMTkA3di6uDbb4D7FHPeaMaRGTK72jc6zZmP0b/GGv9Zpa0dq4Qj7ToD
QCJy3qJyjxNmrrE/Bs3Xo78Vq07Y36DGF68Y31BzCHyZEBhoc+atiZ4YBkhs/zLo
cXhj1Gxvz9n/wfZ/qJAy8T4D21OzpExfzFroYiWxRBBYMbM1g2lnCAknD0qqTR9N
xKx2tT8k+Ez3ogOQujyWheyMxHQNPagnV8wqzZwRU+tOQzzAjA+MxEe/ITDhdeH3
dY3d32++aZrVIF0GwXXQYB96XhmFQWWrbLLgFoJpuVOHeiUoNtPndyaICaFPQbus
9/iwzUGczRtM1E+gxNuZjgw1g0Tp5bAbBYKhx5LMQiETEe2VrbVb5tUkhdfCasZu
YQ73Yv/8I/o30ukRiV51wXBn7k/SD3RB+CNpn3Gp4F17Cu87cWFll/KMkt1C2C8M
LIZyT7MiMtA48frRAbM90QsrXyWhOAs32Qf/HIXuKPw3/5bUt5BOXDvnVOcw7R6b
9GZ5rk70TZGAtVIC/f7Wa8WOwAeC4Am4gdoJmF56q6eFx7vLRNIjXTMf8jbB061p
mqs1h3WCYsafdrA/Jqr6NuosaePKolLKJO0snZlwPwYkDrFprLsZl5vDb/E99tiE
gkFd27r5iNwK8XjPalMntUuec3LxLhXItEf7yt/6XPcYBWO557k+l5f0MWZPNJ7W
Mse7dpt/KdU9fjgPWxjrpWUNoPYhT1zLu6+WXIfO0iGbzEhRfIg4Rzvz8HM+m4Q2
E08OAqPbAmYIP4fuiUy7ajX5NpjewBe+liHjwcmZOUPfxtV6xfEu7Bz1Gejk2kAK
qf2yNHULA7jh7TZ/NqTf912/IywUq1jdgGcxJw8DnbRt2diZHt6V+p7N8hD0wTIz
UZrbgTiykiua4e233SHgO1fIRDeR31HmjRpBasuhC6h7yo4vaEBW1kEAlc0mdutV
gFFTA8WDEaDN8LlWiwKzSMsmMsr39NhtG0Jwlt1qrmDOTBeGBc+2dSmEXkReeh43
UVmfLNvMRMXd4UwBchMjjlpMHwPTZaGrh/Kf74F4PIR6CyxtksVnLbgq1qiLcmK8
UB6jy5mr9bx6fKW5X0JFtPF7LcBLFgw1pOeIq+jTedtZ6kU35hfrxm8WaI0rnOOL
TISsz7bGNsmbh7C/5fyVGBihEQfH4wCfSxzR4yicNCxpCVbt1pGCom1m+DXolq5Z
6/oendHJfM5sn4XVt2llXF/XLWznQ8/9Un8dbvOFCpv2qBu2HC9vxibFOU1Zl3JW
jKBA5MK6RtXslVciFHDTCCrOo/7PLhtosdLIuaiDSUS1Wgtx99J3OGXsT6MGjky5
/iXQa2Y6KJYFbJDnmJjuIv7xM7f/nG1CIjUTa8bnUhgJgdObefhw7revAorVgY8l
EdVx+mySEuK8e0QxbGdzfs21sfBTX04clJY4DZXslG0K5c08rr3fO63wTJtNo9Jq
c2P8UdN6kChfhDjPTi8nbAnV7z6G2jgnnck2bbF/kJD0CXItqSze90Ct1rO8mYxG
XG6EhwoLbB6U9a6tjq5ksKOAwuAV7KQGr952t+mPBVLbKgDvVuRPMrPMI2lUEPWh
AORXeHCsDgkHYcfyfV39M0pjlw2CjFqI+A/p5XyPueW0uWxkvpjomPfatVj2Bu5U
ieExFHZZltJzLw7/XD54UmQXAMzZaDU11ehGUmQHh6h75qpQ9C9HDaXGW+jMBwyx
yG8bZ+KdjCKP1ieOILR4dNWf4fi4TMT/puNHd1q2wP5j70BGCpQrGZYuCWrwXdJY
1M68r+O2Zf3fNVcija6SSSqdHQjhJszTSHRv5WYp90GmUH+GfVZdQR9RBX40zgsM
vERXWmAE71WhYtHfWiB9NYFx/HhNwrMaQYTnKjxNS3g1O2bPI5Gd8gmlBrcbkBEv
iKh3TWu/tKbgHunmUp1VKRmDRNLOKJ6AKor17z2r0W1NLLG3uoS5tQQhPnySFuCr
7VlBRWws+kVAYNjpteBBZCu9uIWTiTvmR2bUT2VTVI7jGt4WTBQT0/lMxuvZT+SB
1XhDUc7Rm3WJRX+KKqe3i6Ybt5pHbZp06snhC7nilL7lQ1tWkxsP+hlGwFn8tsCQ
0jbIIU9BYXMsICkxQoTIJiM9Z4D0pqdtEHPHEqC3I0MP8Nkg5s2cMLa3rlryiQBw
8a8mM2nWYQt63ul3z6jxa36AAnBrC6xw0jgBZAwO268o08tgl3Rz3gwfkxZ7KIWB
JzirF34YeYieTK6L/tbKgrfhjELybJI0rJrOw5V5JPghJ1K0Lu+ZdXgdgpmPJ9Uk
YspJxL9Nm665KnT2dUqTrgqdcGyUjy/KfvEjws6aeZ3BJBSg7s8169HmQnMcp2CM
fKI4bEROmv4C77Kz4ACjxueOEWtqLsHjR0X1EAmL/VqP3YDL9KcmKMZHkvY21fMN
kWNj7IYn2cDHchOY6Aha/MzZMUzeFqCsYd67HN+giq2vnfFih+T2wGtMOZHbhmut
TDjzPyi/KDfa8xJMApv2q3cAJeqUBYTh1/O1ololiUmYJ4ML/a9oDKov5hgiaJtS
mgdBFTau6ZF5KTpGzjio6W7mFWdUTz0mOvLhgMkdzTVVT7RIFmIqatpG08KTjwsR
Ipu1YmXiEHn/Y+MW0AWegFxbQFMi/6z1cs1GWJML4+uYkhNhorNvEh6RctAA0aRq
jevSbYC9PbxNrvXJWUIjVA4sy4adxE6yjBE9ynUpaptI6iKg4tDcWHVQ4C4RstXI
sEdYpjQf9yBolqRUFE00ZTQaxCQqeQNFbmiDcJcfAVe42k1dzrNXViZOSOuGyB2K
bRW91tdh2eMrN2U4GLzSPTFz0tv8EKG+IBTtlU3wS2YX3wYd52CfKIFFEkJsdTUW
bWQk+dnwc70QYSL24/YRyu6yn/UasCEM+AOsgJ/BGYCMt0gm0Du6/sHGDr+ebSJ6
cBxDnWvNP4OGd0lnWuhMSZ9yh0AK/YaRv5tCQ3syrK7nYQM/YBU1h7pD2EdwHp6B
deI2xKzl3GhWC3YD1XvD9Dr2vqaMNwpvH6g43ZeqKrLz2BM1rbQQYY7iqiKoYGoC
tDyjd+iTiFrXYD8HBoP0roSYVsRK9A9+A5C/c2B+8dKZBaNSdZJ2LZ73hIksrSWK
Sigha4gMuPMflUp5W3sV0A38Cm8pM34+tNMd3ohnbZf5NnZlZKdu6OVPaRIJNH2d
bA0HbyKqykem/W6zQ6hFpg8QWdWjlcnIh9k2uN7HGmtF5b0gcFSbtAawf+sft7vh
r0ZyMuVVyh30TA4NfeLlOgwlH89Nwp/bIy7In1ZwxzaukiFNqXWpN9p6o/dqndl6
QjYg+kVkIyr66dVpZKnjhsi1UBzpMl0NrvOtPNAyexAwP26+B5NYRrVEalBb1AMW
3csU9o7Fa5w0zSwWGrYJBM+Te9LO0iehzrJXwuvdsb0mj/ZBYYkb9CAF44qZVcqR
nuox/SpDDQOdk2hFOI5vUFqo6wkx6mI+8Q/N2sMyDJKgZlaqjrk4Pum0aMeTV/me
HEIz0Gn69ZOx20AQnfQXAkCQ9SZFTMX32Q6l9EBFjk/sNpwJKdPTmmtD7sU/rBB2
yUnPbAhCLpKU8yWj+qaGpoY9JmnOXnk038NV7ngz+atxfJVdrvcv3cJzhNFNhRng
Pl0veqcPsf8x9wg0zfAzN+/5/hmry9GX7kPfHhJX889tTwC2X899RpZW9mr9YUx1
6onzCVJvfgdyuRg0jM75DlPJM+e+gGIh9v/tn6cjeBESx/OHtl1Rnda0O9LpCO/6
fskUnPuQ19lS8AfRehUEk835DuN5EdLmYXdaxF3pFQd9A9bOP8fu5X8xAeoG5yLL
K9AFc6NjxWiygbL+BVQzxAHs0EmJUt8s6VoNgq6U517oQZAj0gkVE0jczWCFVfZX
JTXGksqQIcLlUVHH6B8Ytd2JS2wvxAn+K0WtbRuxe1u6ueY67WoR8xONb5a3MF54
milg0C0PSgntRqOuV4W9nVBFAQ8xXjzfTJzDp93oBf9050k6Rg/kSkEJga1jG2yd
hzJb+tCEGUz8tSG3Avzeb2seFHkjQ2OqYYaVLH26MLvP4u/7gg6bbzUOr+TPnloj
AE33J//uojxK3hyHN8nDQmPBQOyZe/zSFFJyJECJ4hc7jJW4R8s/5JTULl7/XVok
Iv0ox37E/7IVrxPQq/zwDxwcEfhYnNxmYj0yXFqYDiW4uvR5Jvw+fgb/0fA/a5ZG
rWh6CrkKUwpZ41IDBqIoY9TRa6Fo4zoNvLZPVAhOWeBsP23jHsZ40AufmojBCdhZ
l04+R+rJ63sqUCRwiE1tNr6tnRDP3/NucvCPyXFfFUvTgxxP604SVOKe8SMt1nzx
aUrgyH1ptx+k4G6dy7VmDYkKbrCIcWuI5ZoVa9rVlsoatvzlEG5VY54c48U6INZb
4PdOsyeizM5NMYqnzGcDSw==
`pragma protect end_protected
