// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r7hlVwfFJdxyKgWz4PCHeeh2+qTUy48bjmHYTOrOsw8gnFdJe9DX2FwiQfxdjBtJ
lLWJ5RTLQZG6qQT+8u5raXja4lp3RrtXgXaXY/cqpkxdhF3OrnuOXciJ6DxjyPqO
93UkKdpQjZW/bXan/DmQqhHtgOiAyFytlJHKJT9zafg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15616)
NVJdZoRMhHa2f9WmORKiNif3arA/BpvWys8k2xYbO92y2Hlz6P3yt3/FVc0Le3Rw
GFno14acG49M5TuBy0qwZIaeX1SgyeXiBjdmI2DVZp7dtahUGvwOzBAmvzJKS/8N
CeaeUgyGSsrxLjRjXlvRQeFMobH7mZmBbvN6MKRycyzikIvYJTclun/243PsiGmW
rSzL0iubJTnU/A4epDFi/rcFRAD84QadZDsbrQgGSLR0ftcChNv5MDqVEBrLgKsY
WbqRAEjFxiA9UFak0SkfL1GDmMJ5Kcw8iX3cp5NFUPV2uJozP8lVPBY+bMz5tq1m
rpsSPVHvOcELrVdFvDtg6Pm8dKJAlpLoBgVcYEG9Zkpc7NGJW0i+BP49tgkkkjaG
yrODAobddj42YpwTRbxdnFh473oIejx2/MeivgjOazyLNiuv29Q17qX62k11Dzc2
6yDrh9ciylH8XKRA65MueWtuWUP9Yb82CFZa+Z5SAm2gr1OLVMzbXMSg6cnl5foO
zwryeM3pJjOwX535DqIWgsY1+8L28M/LvVi5+Hb4M/KS5cDPYq1vxj+pU5QpQ3+n
1PY+auoRNJXMwgix8x9bT89zjZhlb7vC3ZfRi/QKlo+uC2Rj5UkTtvh9kgyQit2p
s48xL568jQI6Vja7FGMzSLzMVNSkjtx2ykV36pUGoBCQLWgRcKAkQyuBNdK2+Gjv
dvQnB0LxbyoJDN6FaDQt4ALj54hdR15QXI34bgJD4vTxofnirmN+Yv/PvityMmgm
4+62JboWFt3mRQ9M5AYDDC/4DH7sKbTH0t4W+T1EJkZ88oWKadgZ/Kg7IkbdcT7i
TPG8WUhCFBlNNi9Tkrs19GMt1XvAYGvcH7DzsdXqyHSVtSAqk04lX2SUXMhrus+6
8dJjGSfF4CWVU6xgptpmWUopATzeAL/KqRBMOoGaCUmr3nxMxb0iwn10ojjX+XTY
pCFogK5IDnHClWSiUtNlCXgsvzgqclLxHHrcHkCfDvzA0LIK6eUIAMTsZHR0wsyR
KyGjKiTcEgo0ij6BHYxmCPNVQSAU7GpG6F/xW8TRvVK8pf8P0rFbtEC37XfLWqHS
Afv9n8Fn796Usw5udx6jASrxhPVG9kQtS+DVgoN40qjN9XThB9+H7guruWjHjInB
P1syXYkGQjVGumHYMowsOQPMfDS945yYgpiV3XKmXIYcnQMNkQzh0wdI4rdzUove
mvcyum4n2lsdWvmlc22JV3S9RNzeDQPGxr5pGubFUqgcWEDX2EowOUGwQdZ0Gp15
4gK9IfSO6OyIskPSgEsTmLPYW+zBmX12Mufb2L1ulSFZMLogs82jfGtdaO4Qc0D/
GpH6M5n43JXvJWee2fbi09zlJ/w2ihMGa6W536gTTlemiGM6uxyXj+pDPM6NeViB
CUVF26q/OrOWLRo1awqpmQ8pmOS7ar9aw0ndU/SvbiiJL/KiJlepFfmL7y77ZK3i
Ghy6kPJqwBayudAaGbIpATlS7FEADEl7VkE9DcyaLpmTstpDDDeJrznbWRCmiHDx
52N4ld0fnOLk3aiNsHIraHzvZ37W38U0/Ip1QCGE9SgNsRXxFxb3d+WJNkzKYv61
q1eJSvI/e9PbW1WFk1/I3QgsLMa9WUrpEdjXl1fckoH/mxr9I9ppR8ut+TA61kFi
9E/CIxgLirSqHkOQuf2cJz+klOlLfYTfCZLU3iSc+yWgABvCcHgQc2vzUYNUYlFZ
CCuHinvVvqNtJpI5OP/xfE87TC2SQc/TDrpZ9+u9SAYFAT1f7QBHLSQYNV/WEFwV
oieCIH1e5LR+tU3N0A/ueO09ifMhNul/tfxhDK9YMM01JkgwrbDH3qretkfUnKx7
MmaRaTdNKu0I7IiOMvaG6VI1ZSKpyDUBuGLs5lbmpS10CkYeG1qpNHF/7Mg/CKP1
5l+qEYEfgzARhzD3yuRK5U9Jx/uW6sqVklF8HJ/uPMnTtzjc7IYR8317+LgKCPtq
mRF6EMc30EGfQ0tbnULp+8ldXZgddSY+CWZiYVI5ggiH56x36cbmBKgMvX791ryU
4RYY2AQAi2vNdfi4qGhHvd41FW4bU1BneOjlXVKToQWW+JUTQ6FTr3pBGUUT/rtp
/nvW+uOCywyr4jP3OgMYJvry7fzcZsyvDtNmeH4hVqmmBmN728fEwxJL18k5StIt
gZDNiq3w8NbWZvZoan4kI8SGwmLCWVglTSYoM7wM0HtFDwDtRg6TIj29smDp/ZZD
iWgYxAxvMjQFXUiKodjL4e4nOQ3OJhPTtadj6XNR/uhAPtwHStVANteF1RokoH6q
fO+sky9EKmTDw+tSBaa6rj3MkekzmG6SR+4zREkE5XfyuxtzKAHv4/QzeTjsAcZA
9YP5vx0Zg7BQaxQLmDKjR1TvamDzNN9KXHT7CNGfXFt1Tml8yXwBo46LjsMycpPn
Y2uedswrabFlrqJiWK5oWAgC6Nd3vmqCaoM/8WgI//yRE70zWaAuBgETDKN+xLC+
c/RYEW0m+xwQ1ktcYRITj0g92Jq1sYjXf1iQjjvAni3HMVavtIIyiVWLR5JwCGy6
qf8h9Qppi4T+neBPcsrW2h7bTqsBMLNWfVY1OYlFnjBND/ulQZnMGCiVSCjgWAnR
0B2tN33ZJOr9HOOf0waHJnjnuoghJSzJscUXeI232WltqTgSiJXiuGzW47FgfRN3
aDY2O5RmycqGKR0IhAeCsdRBzuEtK431Ht1L9e1TCg8bsYUnqcX1twS8pMveYE2w
gMYz3G9jtlQfnd0futg8GLVYH7WvWkF71ScadfuSAIkE4vzn/KyhNERraZuta5lw
C4swGCePDV0a69rC9hp0JXXhYrt9lTvz256dy378ej4DW/CForPtvUZDy0OJSmW5
sX04hWsyB4kNKBcL8Maow+t3kB0OEB6l0VC5fN0U2FGe726yuNT4uz/lvLcOC+Bh
SrHzs2sGnfRsMe96hnalkAyukoHesCrqWgmNgoW9elNHjFXR2w1nK1ekDYhg7nTN
rxDh3QEyDvqn2KcrDUrYRIqRC/r9mHpizMKl7yrfRsE5fi6A7LxlvskOXZJtGvJD
08kVqphB3gqFxSNVVb3VYBI0UwWr7aUjhxCulku3VyOvoFtXNtWKk7gij8nQunIu
DiqmVtbU1HfPgJ+ubpkiKMOm+bdZ6DEpIaqUzO5VaIyKtotxcCBp9sj7OInge6sa
OPAJVAR5zjRK8IEsPkPllJ4Xs+27x1DggtVncA0IjVxyRFVwq3Y9G/ZnkP4w3Axz
CLy1uytH6o8oK3qiWSs7LdUVWGNWdStJtp/kfazvfOBBCb8xrZ89H+wmzbRggJT7
7Rsxu+2SX6zvMCGWD0Exj6p473VkJDmCJB4J5nEiJFjjA7ZJzMAS/d/pd/dg+C6h
psNoocF3f0A8j40WPogSaIQc/B2tZqfijsZQwfK93ldXPPOIXLxwIllg0ZU4b4x5
0+zNpPOYwEIuorS2Z8+yXuJ+NaG636V2tGSuYoomTayYdrlqLy8Ci9M4HG5uQhhH
4XdGQXCPIyoh7M+uTpSeJL9I1WazX/ILHXpOafWJEuOq6JC7s2JQbVZTtVNOdFrk
6U/z9py5fmDgC8P8REcIPDHwYhNjNDjw+ajacbeheGVgvzpsr+nXhMghfD9z0E2w
a9eEbPhd6EMlMgx923HqD+fsaisJIigUR0oWLwDh6iRUwoy2EyCeKNJC/00B5/kh
GPFQ6hk2D2MccGQIfRJsuXi+qOlaCenVizIhUmIHeWBhlEZZurne5EL9Jo6nNUzR
qY46oSvTT8a6jNdWHFNiVYVZ/2tny/1JDMVfr9JUzKnWnRQxJxT/jRJcK/psR8jR
sXyjWttKwFx1smYSkSeIZ91nJ/N+rJWmdrdL6ycX/PPG8tzFlGpcQ7mgdKKM64PV
y+/rA4i9JN7Bcfamer+VsG2BPB2mmIrhCOfhP4ThxKaiksncayQxwE22pSy8+QCU
svGjDh/zHranH8AeNuV7bod5R8qhyfPSDPSBCGSizoPvDR7rEYVZQp1WU3rIGoWx
i1ThBvWnWIcB8HN1f1ueMauG0Fbz1WmshsUCgEOZ+Fz1zppbFFYDw5Ch3ILDwnF0
uuZuT13006qAT+pVEOHe2jjKdJjHj7S2PzoDncJdznORxDuyaYXX2vUQ0VfMA3U/
S24ni2rsvVtUGfzuQeOyALqk3zE3e1R88cGpqOiWD4mvhh6Zm6Ns6BfNDMU8k9Ve
xVM9PIHekRjMjrC/VnwQQWoT0rKLZTotIKvtKDX+mt4B0/nLql/9CgnJT3EvALqU
H+TeImOoBcyh7mSxDQI3PRfnZFMWF0F8X8l3Qnmh9gzGU/yfjpYDWD36ncc+rfwM
B6yy9Wlx0dkFZCIcXE2tBeEY14dDl6Vrn4NOE3sNscIerWoLm3+Vvh4oKj9xkuwv
p596pJGjYkpVgHwl8qyGNC43GFIknCWRzwg2oh6sezVcJh1hUF5vnWBXQyxrQWq/
4Wd0PFX3qJFZFgUTtoPJhhnH4K81rKx62CoP2eyIsBtbtZxiY0fCmmgc2WMhR1aw
zykHXPag3XDxVxEAFzUezrAo86rYOcneRxZvZZvBhjMT8Lh76X47twQXUhaGhIEB
fOeINst8Kzq4XAAlPKFyX1plwxaI9d5ogChO4h0Af0AtpsydMNfy+PTP6jUA3PWR
AvVKBACg0yublEqmDIxIci4LTOFjTI4rgcOtntf0rQ8cLDo51/g/doYsQWhQnleB
6y4yRf6U6b7mhxm53zwGwc/v7RTmtDIdoyH1B64J6dDbLLFF7eGP4Aj/sOscz4Xr
3MQicX1WWxO4sgn4RKzVb0YX48ld8V5nb4tFBs0n+HpLvh1f3aJtSB9ZMM8Xylod
j3aY/1ZcM0QSA0laSEiuTWHVvAp15hg+eynIfxByopw/Lynki0vxrbpzPl1ddbC1
46H9JaTnUYUx9/6rsuhF9C/4Xb2mg9CA27xvGcY76B8EwcuFKcgn+FRu3zzrDkAZ
9tS8RO3OuTIbTH5HBq0HMUxDvc9nKIKl8nZh9Y0E+/+YGj4dwUVSortvYmPak8bv
+G7naSPUwk+xmS9fV9nAn0WUbyhJ5QSby0L97heLzj48j+tEXa3+VEGuNhut/zDG
nHYCoC1eoI5sFmGHIs15vZmKgXQ881lGUgTBUWqLPEb6FVpWnl0pFFGJf9SokunR
Xl5R+W3v3/m5SfX2eZPeCPZqSMYr+UOZvyMjNXbK91oQ5r+n8F5WZ2qGE/iIodPB
8yviHlvkuvuWPFOFKbrXSbO/u0kT+3JE4Y0vH8uEByKTLffTl7M6++XBwqoyKq0T
qwG8uzqexToFTfM5rNhNb9+ET82RsML4wTYbkxaW2kQ0eM16dYOEI8UUGdp+54kG
RuJsz91J8+lSIizl+rx49wzj5fJuKd88KL1x+i4xnm4HkDEOVDTNbA8+aoEJTUS2
0RyK5CAGy4pZUDjMOmt+PdCRR09WzQR/31QSStjG68NgaMXPxgJSELuHP5Gu+EnA
oSjzryH0p7JfetcZYd81BT+tiHuzkQwZ6kO1jaDlje7cqQkK5zwJhQ001UE/uwDp
gbC2sS/wV3MsnxXqVuBICPFyGrzgEdEfkemEXPfaV13b5MoaP99llObFn6rTVLbS
ezHr4Xv9Yp8TiqXe52k7sMqN0NJy0VPQy62TROafIqJg2otnduaQNjMTg6LubzYz
hvE+A1AB/5qwLrFrWM3F2Y5TCxkQhS654uWl8WXEv2GTlw10bpdu6wurgzeCIg6H
xoRSgor7K0O2+atlLlqLMwk3V3tXos0qqol6xJy1xPdkDDNrbxdXVWUtb+CWiRSk
M3nUNrnfdXX7S2/UHUzLAfMU8T5hVcOCj2thYniBKc3t+wCalL3PXMmIC4txphgR
aEXuP//efqO+QE49axnlGHhUSJ8ABPxebuPB6PHg/Q4X3lw3YQ9XUOxpbmuPtLBP
zn+R1hUl9PG8cmRkHuEN/fu/6G8AeG0nerf1n4EsNNin4YFSrkaFkf/mJZK+3EZ6
LP7zxR1eSo9vehrWciX2GyHNrhY5b3A2AcVJS6FnYia45wGk7Sf8JQJMAfTNtdnp
9jmU0rd8QsmqqXpsBV7In529ndeyqTJzo3kOY6LmJUbk9Dxhcg7kc5OyqfrUqtXk
1OaPTb+pSo6MRVL3QGMnmIKDVNiInB9o2Rm6hmCNK0sNnIArV9Fs9Nx+Bbj2CyRG
h3jmNlI13113Y3DfkaXev7dFQkisKPev1i4J6lqYjK2kn9X5U+Aa1vyRXXtg/hUq
VeDZ6uzYxDQdbcjLSojW2If64mJzeIiBFQZW58hasuM3lV423kHjyiFhDngnyzgC
6YxK6Xi212ktTzXSyl5N3Sad+qFc4sfU6pqpEUZ4/+ikRj26c99+3Q/WWxOVmpDO
BUZIwEoMNXYczmY95VU2EGRrlPJOWO9U2Gv/qgBBnR2TYwyVDy86qIhD2rt7OJ7X
TD+2KXdnLA3RAea5owF+mWCDMYUFsWh5T9hCeQoCW3LWZbW4BpNJo23D/XcgTe1B
xDzaZbXDBTNRwnKWniznzHL60gh246jqjG8sOoxtObhg6mw264LsDnAA1YJS9+qo
UYqEZ2nFWKR+XOdES6hs0VII1tUEz8FIgrVZyFUclaAKr6+RDM+1KCL/bUJJL+hH
5F5AaL7naSO/+yU2pfmz2YZ+xsr2qJe1xZGZGnHghBMWzfnFxlCCUr/rr4B3GgMp
sNIUA4Pqla5yr480HDDcfUXoEHADDRpONII/9g+S/SW9s0FG1Zi8wJF0eWTdCGJv
K8fZ8EZoRt5EQDON6Ze2NiEgKvbFQij717Ijo9J7Phd6cvATTtCdjexjK12mxkJB
GEAllOs3ggE5q0lewYdIxSzQT/zU/TOp1KUoMlp7N5s1IrCOlJ8KF438dCK9WR9U
zy0TCJN7dxUK6rycm6hJ7hToAHytUfg1FqWXmZ1iHGm0owmEMfE9O8aJcA0CLDFF
DBB52BsG3mc8sRXjytMbg3zwEqbEWmUluZid76XIKylB3CXuF/0444zw6xR+DX2e
BA/92SXpsWJGi8g/26luyQrtd4Yvm4PFImFI5/9S6OKShDKl9DX5nTMij8ngB3jp
ERfTjzrirMsiVGTHDWgMKbBb7OvUHJbOmpTP08rUO3WaKbrVH33ugLcbe8adnF12
L+WNX3oTkTN7MgfY3/ISkG3ea1cGXud7rTeVonaU6QkHbWSU7jMAZI4JmkKrYSAl
XTuEPCBWU2GqNyaj+9Lzhu8z1kUWVFw6UUZ/4EulL7Z8/Jbvxv3Sbp/uJXX+K0g4
fd/Q4yfUksP3tHLmjmQhpujyw9e1HDOMN4AaWaOvTXua7HG1egqrms4eFkgOWE/l
YR1R8J9QqeyBNbhKymLV3TpwokU3XvLXJTZMGwgLTp9m5xezBlKa50iO6ao5IjVG
6PxHpRABarVC4cIxhOvZHMhUYmgCe80zDZaljWmVY82yJAYlaluXCNduMMQt9kPP
OXqtYN7ULnhioBX63ehdY+5MboZNv14gJgrejNgQRcg5sA6DSkqUq/tVJYKb9Sta
30QW2MOgUCU8S4AUMlhV3l97kAi+WltQpiFbqCIxhhN5+xzfsgH7pVK/xVI//A6J
oNwMBxUeRSbMLwBKfL200SLWAr/OSK50MgJbWE7cfjFCufRlPkiFGUzA13Pgp6Xi
ko0dLSnBk5zjBkwzf2EppkNEmnvcON3U9O+xd8+Saam1Yz8I/+pOi8kMQ5xetcuY
MnnfwFtaeszqKjIrU0TFBRC6EiA6l7yPdHa9Cd/+S4xYclj46LWQW4SZ/s0+Dwyc
1OU03zUgFNLhMCp9MF5TY8hAWzCSZVcnhsIKprVoCwvREsKWw8lW/OsgPx4TEPWe
eTyat09W+QIAcqk6HqqQqFsL6CboXI7AAp7Dw9Gj5nV5smjR/l+9WwY0MwiGFtBc
UppacNTl/C1sZ8wHX2y0i5jw3JLjD2qjxD1hk96jOUeROSNjX29pVSdiFW3lu423
qwFbvHDnm3xa4yX3N5UY3qsAzzLcvxfMLr0RN6HAj7wVsCfqwQ7FdRbQQAQ+wgpO
/j9YyfZvbiY3n9w8J3IbT9rSh7tY46qm4cptC/D6d3x5YHMBkFHIwtbuqEqjP2cD
MKWhaptgskZKpio6JGy94kuCB++fWH65K1B9U8GbJhPrTLA7YXho5Oo/25MsLRsz
Z+3MEe8ZvimhgvJ6t4M7PRH9ngWbOZgdzqLDyA2+IrPQc4YYeK5VTnU5jtDSvXgS
sPEDg1XTZjniOppH/v8fC919Aa48ZV3h9R0aA0VoFn3QvuOuwSU6rJi1A13koeYf
GeFA9Nv5NB4XZiZWg1zT327O+0mdeod32h79ZqX3LauCD1NAxyLPtsEbpIccIWqm
leEMFewceejAcPWX90nrVkwy4xlBzMCNN6YdREc9S1gj048QMOsALPI0CU6ltbnd
Rhpbl3OhCdgTrEHyJtQ2o+G5tB+8vScVrGLZ4k7AYqBUSOuYLr0R47CBV58LaBEJ
wALsUckrvGyO/uQjz5vJUwQMgPQda5gCYyc/4tY1BGLYPHuFKZwSHtieZAWtAg+d
4TDUrYkF0gFSqPrzmy1+qSJb2DPq5VvJyJZgx2pfvfidGBbjR24mmP2Tm9RijVKW
QtCM1zWDIgCFz7dU4smNTZjtU+3ZZevYX3L1yA5qNz7ccdJjOqMEYQ3bBaEXyumU
b0QNoLUj4cuidds9qP7du/kzF8g9Ghk/78Bi/HFufSp3TlArKTJ9OJGuNbrGchUY
JnNKWOHdprEzsaHHSonZ3UgVw+KEYSskoFIeX+uJpow6ycz1cYZIaZlvrS7fRSkd
gf4BgaQB6skKBTDOY4hDHFBXkW1yr0MEl+jyMbzGRcHLgwtgXKG0Qq1qg0HJsAuk
uL/yJiRt0ok/GU9mHmkXT57JvkLW41r0x4o6t+8Xuxz2GEAjggomyDmRLdWffAfb
c0ymIS66HRT3CpexTmNvmCU5s9unhkC6IlSwDX1D5lBiJ5GyKYei6IYgwt3UVLid
R7sOQ7fI8g3ySFTUOg5T0+nLc4DqWc9zkrmE2Fw1Z8SSTSp1MplyvHNT/dj0jYlk
WynPuGFAu8bWCaNqiN0FR5wYsCs46YwJJlcb96Re9CO/oeRkJTjm1NWUoq5S+tgr
b0zKoq8+IgMDmKTJFv2jyyUU27Hr7x7b0VWFrxhFHL00tVb8ZIysiYU/NCI6FSB+
kXWFqicVK3mabOjSiHClunGuIaSpCADkp4AoYpRcvbyIn6q0o63p+7YXIzp8bqY8
WjkfbAcG1Jv5rmUeeKP1s2fDei3Lkx8EmZZQHujmhopl7CjFjJ9cKEfTz4W8iv4H
iZs5bSYSjY5/e+nzrpH7vbuZDsPaG671OUm4BAc39P5/Cpge7NYErjkN2K7FJ3+Y
Yh6AjMl6pKpjxrCn73lpsw96Q0JWXyL1T8V1OGXnD5VjymCAaYa8G+5s9vjivxn+
brqbAb9q7VVuV2wmCHQw7ZGE6C1NN+tjRgLCLPD61523Zus8KOJjG7VD7dtqeLB4
C/b28NiIuwltO64IiPk1G05+pyWcHgqPCR8tlGRA3TCOnMOta8O0CX7hD9ZG4Rag
aEG43JnYmJrSAqZ8belmrQlk96QNVWs/C67MtqCl/JPmb7yOnXOATHQFn7N9V9Hm
/VYQsmlX5BLvEnvd9vQtJ9RDK4ackz7IY4WQMhh645vbcSx8TXHfknsIzgrvHxoR
f16OM0P/335McwrxlS/doekOvEcDFpIY7NPDjWVtpppxCAdTxVPlZiUeqaqXWSHu
hPbBXvGrsu5NwtihRDL/CtmT2ZfDGjzdypp2JuwwJUliGkah6rcqFPibvXJNTaih
cigBH4T1QC8WpcKjZHP7yyqK/FvtJUFL9rDmdCj47o63RdB5Ai6l7ed9ILbTFlNa
QdeF+B6F159gJiDJm42pvpUdgb/WF37SZ2lHH83zh/XjlwxYRiSGsZ/G0CMcQR6O
eV5VIci8eLAz6eCC2LA34KhFRKfNaZkyFOTFZhUPUcRVTG6vJ5Vq316mVH8F9HKq
IQ74iGI7KhTIgFA2AL67uJNXANJxdEXm5vwPpFn2jcT8Z6fJtID8cAMT4ieFHaLA
1GFMrWsm+A2sL5gn7knINvcBjWUepQXR5gPx2M9+GuBJofqr85UOUIOm8MJQYFw4
uXoZEqNdSJtaKFG0iZLu5OWPrZFjOUtPNqPSzszfHCgrVilYQRqh0KQ+nvi2mQ3p
z7yuVvsPN+eMs55xYMwoBXSZlNcuZ27XYVOz44QKsWj2fX3hsHodEpicsACEf8w3
Ro4SFPaaSJ1rnkc1AUB5VeDHV716Nt7Ht2+Kb7nqEN1N9oiEOEgJ/I38iz4ImrpM
2pq8kPqzMCuzV/hYkmKG1uFAgdS8QKNYCLeqEsw+3+SMz30S/RFqUKCERCc+TAYj
WYmOMfL7iiVK4NAGc+8g3i+I16Ec7OPawbmMKe9G7mXzhGwZMlwfxqmUYvmG3jUt
s0Fwu28iieGPRdnD/q3TC2pGRII2lNSxKULJszh748G21IeZVWg1jOUfsQJbXicU
AqFbnUCexTrJvbnOc5ekkPUCtsic0lU0Sz79FV6qt9ujlbBUg5kRXoj94PqzXlGx
Oj134sPSKkHQOHWHGwMZBO0lrMEA28qfSFaL6lqMXNx8GrwnPKT4j15dy9Vs5ped
4wEhsX6q/9U1+jXUxqDY73+BK+a6PCcWLwQU5+LpzeCuuByiQzdEum30iEuoqBMt
zhkMvzjLoh+uZJB9dNyU/OalEhgRnubSI/v3u5djVb45ekQE0XLOH2ZvzIVCJAGt
caLoi4xg2l6FIGZCIFNvT1BKC78lRmfheD346/VZaDhmfT3irqYQjhIj0o1xnCO5
/Vu9aF1oX5zcrzsf9Efky783FxE+/2GzsmdXCETC6wdINwhGTido06oi+/7hlSz6
9Njt0Wy/5dX46yUJ8THu3ejvwTyT70rRVPpJJjU852bJvVybfKk79+MghmTwQZ6c
oQwIc/FMbBRvUVqEgDD/mHqt78JcWV93PpMfwu0dcnW0u45mRM4J8F190UXNSvPm
2u9Vyg8v9rO5fq+B8gKyO0gIoZXArSKLoYbd+yl1zoZUqzxk4OakBW8A9DRwM2WS
gu09O3xbrxf3zC8SwYz4PJwQ68SLDoayMU52sOAVcId7rJ3A7u3XU+5N5C1J2Eo1
Y/wIjojac+4r/SJOaXJeQwFPbNC3tUo1fxnyaMSUciRUpNwsHd82s2PZT9bZe/uh
D13BkqQjrvaD/UJW6Mfaca5SZbhNZlaVCLa1tSLHs2Ylx4M30cEwT7Zc78VB9IOG
Bf6GFL01ll5g0SAP9ikIhOXoQ9za8QdbSClIi6OU65vocd3OoMl7UjkaVlHzS3Mh
Vs83H14XaCICFz300q1CyLuz1Vn1x4HIH1wHVGLws/Su06/XekMQT3U1KABr6JyR
rvy4QGMTVd7aBBZ7VSTKKz0jrinrZqxpJ9uk8HTIcMBm/7y2kFVyGi7Ld6gAbo2T
+/E47oG7jh6RoCxvao2rpJPtr8hwiJIBksUFyBEVTv4kCwW4wn/B5ySAldRfrCZV
z0f9g7corsuGtVT+bmJIAp2IOF3yuf1GgEEoM5C+cZRtKGEDSjBNE6ILohJFYTA5
O7yapdhd6txQA0Qrs0DIJlwCgU51Z9VRb8tXa3J8J9lUwRB19tJpExvPHf6YX+IG
nSEiU8WEK/aeEnS8LQeXCec3rUMgyXZPjB4kvs+QgPVoKVsWrYg6d/4uQCBECKQM
x69kjCIhr3pm5N8ebPriLyIC05LqvZPZSTiHGVci3BFWRZccRugO/ll9leAqthPp
FXBdPyp7wkNWUd03hQP4hMdG/T70uvfzIa6lKoIdRIjBwuHkZZu+O28+SVCQU5IV
q9zIdDyqdM8NA0CZAAnuZ2g8iMz9W/kZKfUYXb6oHbPwYUq8RJf2y7552uj96PPh
Iy95Sfxt5TtxF/H9pCg0nbc7w9gnfY3qus0mDtCKOdqPqrGlhuhSNmuzrZwNjKHe
cuWLL7WXotjwGZNdKcVjmSRwjh4HfiFWl+2CMd0GbXEz4Llyz+RCEllISiAATyT+
ytJYSiZdGMgweFVRRvoPsS8wherTeywguzHyqtIwqdLKFtjiyQ2uTwTgXW5KSnZz
UECmhwZpKiunf9CHDVce+iASdbqscvka6zCsD8ENlubrXjiIy92abd67kTTdptV0
/3HaUahJ66Xoq7DYUMGH0Hl22FBN4JKJLE6MoIwoBdxHIBHBoTCNfqyBntua7/AB
szblp6GCRs26i6pqkdg98g467mzNvY/rY6Axeius+Evh+U8/1sznjWhKORWObe3c
FOyT3BAJ4kx4x/xLMhSsrUFht7E7eWwGpj/SdZt/cWtobHDMNSDuSmgEpDpUAvgK
wCBtZP0QmeVmMYmsScDYnBFJCR48WADjokqmvXmP2cYmKn0+V9lzLhRoYaoR3jSx
8Fb/ZFJO8cTc3RhLpdwsqDsCJpRNCuNoBhK+rvcxknVZXCkhyhub95rhEC9QwN8i
1hMi/tMqzGmZ8VGbuWBdNsd2snG4YBO/RmdgGVBvoNSXVzhXJzJWxbEBbfY4t+Ex
gxRzl/gsPHxohr4u0JPdW6ja5kcNpI37FlXaVYP8yh15qOoSgwRq7nybri3omAMW
nUwdNgGna8EoewFH5OqySGa36IYoBM/74qMMKP7GHQVEVNB3csa4sfh/7QFLgMxA
RF96qDRCXZlvVMlYbT1BJSVWNk7BrWkJ6J26ptE8kOsNrfmZv6GmYynAZA6ALRbA
voybBHUu6sOSu9lH+vN9fE1NTlscDtQRohjbF/ut2HE4rckQuQOqjwn/h3oDDDeT
lpr0Wu1UKrtY64iaAWTPyBYGKb9EjkPSb8I9JPizirTevkfROAzipuanOpPnfUCT
+CLR1cBnsddwZ5vGfS8ba/wf+sPVDn7X+to2KcWF4UB1nlu8NzXbNkn/xrUhu9sv
087W7F/JLgp6Dbrt5MR3Kmz3mgon4mkzsteUC0hPletYByUrERFOC4JYfAmzTZUT
7skQrZouyvXqt16jygey3BT0hiJ5o5OH02ZpXpo7t9a3hNp1aQwGnztieeNDcwkG
3+XCvI63nw6JVg6W42PNVod9jsr//SPEgt2X4+laavhQBPR0//2Z1gs1VttEBkqx
jwCLrp4XeZc46NOTEYxeV6kkedrLCHTLBz8RTNjkb1yqEE2U62GhBEGDMkLAxPl3
Ts5SZAO/UPL1omiWaw7/cIlAdfll0cLDrWr2rnx0LQO3Mui0zokn9a4t060JZsD5
XTPOLSziPuwGbCfl7BdqNOTSTHeWTFY/HLAVygH8WlqTt6twJlUtWJv/S8d6gtzl
mrVl263iWbb9Qa/D4zGIQsgPOq536f0a6MoOS3FRX8uwx0NrgBRuV6grtMeIonYF
FETQvonEEo3dM3Y1I2vXkfKzzlXj0ATYKKUn5qaAMCrlGVd3cCoKN98XyNiY/Obc
UZ3YS8SW96I4nFmI55BL8OUJdDRoEf/cGiTM5F6ncMqnMLntxSbj72KtRSjvvc9X
NzvcyOtiHWPbuq8pQ7ObwQKnwvLe43j67i7kOOJZ2QQnRlGGBSH72tuxC+aK/pNL
UydQa41Bg5PVphbdZXMSlXMmtFZpaduBw87LNVLFtSRsH30ZjNKff0DQY4Z5ZjVB
wzy2RUdhAi2XmcFNaHKKKKMKnjlWCnaCYTgGgGyRtCAWqVBTMnR7d6jG/vAAwwRW
lGvBSrcu3yUJJgsIVuhakQwIIGHMI2PEGWpnWzJpxWE1Wh8C6SgK/KsYn3+JyIDt
cvdguGDmIdEWm58AcLXrPT78LheWqgbgok3CckdfP3+oJyU5b57gdtBvbj7Nezi2
4SFhKAlV922Tqa1KU93EP5jkba7OsB4sWIC2iojaWkAWTV8+W6WRov7WG/oGdRGK
bqBj4LXAVOVkjGj+z1ivjz6E1l9026wUbP73cyZ7drgmwpizSCR04slnCW/TfJzL
rsPvyz2/wH6a1L6Un+Hi/P403RtjJ4zONuwVy3EfGm39WTvBTDQKiMnNbbhu0rV5
nQMOBtU3jDUkAJtew2/biyelxuDuerMoDXWhkyBFZcEBwGVFo2qpsXPoqE07F3gc
GfV7AT4td1xzMhrURGr4hQyG3d2sDahkQZyclkhVVIYbVAEo/gTXkuHCcMpUB2te
rT4f+xugi1vbAauehQOVeSbr6gWEqEJ8HSXeukidWuXWXfFTuALnLW4CVNNtO4ai
VZutY4v8wiDIK3Ym04x2TCITpwbuo2mN/sFJkGYmpAu14ovbXDqESyhn+SWFOnE5
nRQHTqemBqavSa/jRBYEEm2Q8aMrCGLF4QGkfe1CWxR4nQ4bNeLfcXjTU9tP2gzQ
pfsZAgrBTZd5OYihwYWG2rvm9NzWdAuxO4D03IH7mfG4aqIRyvVndmIt1HDuRVFC
HWA9JCPliu2DITTwX3HCBjfs5+Mh49jKk6+4O9r+m6a+h07O8ZBAYaT9pjlgjJyP
oPUegArKe/QCXdLOmCTHGswM5Wg6Ln01/+cDycAvcOE+ov4qB+cTzS6Zyigs04gs
zbqg8v9JXtmOZXJrNbWBqnEGlgVTQCSjFzeOrgAFsm+ocC5TRh/3kjVfR7xgSgXv
ZCdBY3UYBM+/i0hilsQcyVvqlrkNgMUGt5tauhsdz3LsTqocKsTwd11bICUc9QnY
moSZJ1M/Re4R/3uvtrCoKIJnyn0wD8HBHZRefQQ3fbJOjDCDWvBeSC2Bvi9zp839
voNyjDyd5rs42ruVrVs/G8wdjIUdeNdwhpXxectVBiQz+CCOIIfnr57M0kaifW2x
zkKtjY/Kt2Om1hcxj6iDlxHNmNzc4tEXQS1iup+bmxjFWmTJSP7OysKo06xFpihN
Z4sjn6SnLTXsAk9DP19mshjMgGoWjZmMlh+FH6vImDB9p+/gaL47tP1KixY/q44F
p3WvHS7dRvZDRkJehxAQo9LsVzHcbm2UV1jffm0dhwJxn3BNfBe/9d00ZYy5jqcy
wOfwMZ2MJNORAlFwLr5+e2uTlonaiklD9V/sQ3g4nbhIq+L3tGosHqRDpXplcyaU
/WuCVmWctF0jw4yLp/bNMuOCo0+iu/dikHZZDioTWZn3zn/EB25xLyXMLrgBeCh5
lgBzqR4ZqYLtXiYR+PJnLywogZDd2npyCtxiqjb/Np5gtz0/jP1DFmaILTYl1GwL
LCEuB/1BRJqBYeoyU8chSps6Q0tvDazxg0cPy2jy4/zJmi5tjsof3jubIyQMKkUU
g7qWyD8fS7oSk5HFDzw3EY1y/zxd6gKjY/wN/PD9BNfqSB2sM+mGM4/TJ4sXbEQ4
ConCxPoSDlcK6zn6VuuIHLei46586cT5vdxrJoHvuSLWDAF6vcUWgXhKtsdCb2aZ
t9J6ZnR8UHnK4jP4MCHSNKZpR+q9rpzG6DKSxEeDmpUUhQdmoaPKvHvwo5zoPsDj
FMQAi8zElcMFQZIN0db0aDWn8xt2lyQaGids3sxkCqlJxDWJg9ZpOD9un/bkj696
0PDzd4kV6TmMJcgLxjra+aFpDP3qP6Mvz1HLHcnkl+tZnFwSDmbklKwj8y5orFts
wDxhRg1X7vR1MHbbkJP9E/tTMkWoaIpaRggJqJLkGE2MEIoo/bSjtHKr+aCCm1s/
2lkNSpZISj5hcj6od6ZKcgmfP2s8zdEYPxLEqd0q4rZeHbYe0qswWS9qT/U/Cf2K
9UywZiGPXq/SRJrSrrPIzj+uHyakZVWdPaIZwomNUy7iCWbJyrIMvkMZe6KlX/99
oPNbtoWviAP6z0AU0CqiAS2iEKwGmzFlarMxhOsd2ipowQmQ5K2nOj1f0ZOyzRkj
QwjKb+mX5bep1h10dNhKi+CslIP7Wt7UOYESR0fpAFmLsCgBum1FJ6IPiWITpq+K
8cE/2og2uQ6N2x4MVJe8GH/brB/NEESWSBAaZAKOOv8F5ekxtaUjBGWaoPK1Iih1
/a3crLJk2Jj683ZX/AZh9DY0xe4mQeK9i9y4zAuXpCjpgNNcZpT5J0IGz7KhDy+/
Ifjt+3nQG1TL8+893TsmdV1Cr5TR/tXWNpeacz5hChDeXNozEteRygAxy7Q1N5SX
Dr+NOO5Wd9SU/yU5VMbl6Jo15kviHFBxq5CP+nDzVlIwKLrXKvE+dOtMr1Bc44rx
GuxAVEW+rZMG3D5fxkdP6n8qbReU4lLgJPWBoM+67MzVH3B/yP0RRkv85gO7CgRc
Zy/53DVINiMFHBPG0IHdN62pQjcOQ6LzeC1FRk3/u2MaFSeFClwkJCCmC0aR2iCt
0vqxZN4zrRwNb4yFbZFUQwB6yuHW/Y1x/kaB6dR/U2BywN9/hutrQT2fWseZ4Ybn
XDuIOUj2ljHmrlieuEeGDxpVJhnHBEn7cpDp6nKK4hwpADDLGP7sZyJ9ndqgZmuI
NdWjNng6JO9lItcgrfKRk0OV83sQbNN/kr/T2tZgQGu1nzAGmgXlspsHIWIjwpJr
QM9Xv09y9R+up8UNSSQvlFUC8avC29DIIqao+T22C88VdV2I0KyLBNnauZVLFyfQ
Z9C3aehYIZnz1sq6YmnD9cP+q/+/lxli4iTwqZfNo9g01uUNeUWDro+1k8dp848+
xsKMDmjcRot0MgjbRDEUCyU8AztBzcB0SqFHDE3j2ZsV+668zCPecRTjsdVx5nxG
4TGWW7hmsqpVsZaSEgrBkw3YFm9ZUehC+mkDMD1l/7QUxuYDXqtJlWF2PyEYcuA5
HLCjCkMivfeD0CzOQD3sClXCOmChUyvQLAIaeOnTYLbEKyb0SQkHDjdaD4kIClEC
PDG+UXeMXd8CwmcG4IJlgt+K8VLmqMvPkhL30EsU4rTi5m3aF4Qx0fUbkLN0mzMo
GhUcM7UjFNZptloJy8vf4bFvyS4rZ5yx6j0H7QVyT2CMZRsP/NzPO7asrW0NNXTu
bb8aZB725hHzGEBs75anvdIv7ULaL+TWZSxl3H9PZbS6u43LRy0SNrhcpogjPlYG
rJMC5NMc5hhbayyzXpwvnGg+G9yH3wiX5Y37XQLTXF4qftSYg9OWBYg7b8khG0Rd
4MCrUoCLY/7JII9J0CPkYKo1kfAt4PiImjNHVe1XLAXYDW87ACxxOdeslKdBdtzU
4LGnzqGeraApKICIdrXa5Yc6uJFazzDGnznkSX9NIPapavoUJaT0+/9khC3LHeWE
jzaz7Ztw7VxqWHeJP+QZJ1YhsXnr9YtZxtvdPBrAvx6pCjJgRDHK8Xjq62DbD4HX
vbsYfzty5PcgdeMXAPlQAqeEZMGHQM2vEw2cgfuSH7tslibK4j+3pwQ09eFBySEg
COfhl+C6g0MMrIGo5CR6GN4u1zMIQrDLBqICTKV1RZtqdoMLJntNo0rg4LSqKxIN
ad51ZMCWIY0SaSM73qlgHKeqDdFf2v301Q813KmdTsJtVbiqZ0t4D4qgMWn/GOPK
g9WFSd0RvqT82hkVqK3JcoUDb6WeoCvZ4YYEOqU/Bgor+JMBLcyf84+OlPQ9TtY2
cn/cB8ntuvEqIJ8qDZIkNjyb47TxtwYa2wCmO5JL7x6qDsmta7jcMXYDldua6+QR
eA8jzYv3mwibCmmzbtCZeZZ7E6o25kd2R8or96hQzTU8I0ngbpD5PQBQX0hxbRwg
VeZ43+hn7naLypPenRUWa2pkE1cqWFJUSPZ/NF5jAiMLvFSaW18wBpoF+hy9lky9
Jecotjg46D3Q68yp4HR2VV6Myk+dyZlUsJ6aq3ktoQvIuunBuJ6ert/DElvsDUrE
xZ5wRZex+DCOeN9m07A2eh5cahyQPWXM5obPPol8t1XrVKmOotgOpODkVgLMgs2C
jbO3lLYDiCvSqfYGpHI5qoLZL9IeUfiM59CvjTNGiT/aZ37WYQo+/4PuxG4Nd0vr
VU/bhpvoneFzW7Dsz5eH3DM6tMR1AicVQsB70CTy8bbMkIuN7ACsX00C8tXxMnU2
xImcd56YAGG/fTyamwnVu4/cUxOPpOsgooYVHMLq13tPBcCwN8m59RmKBWg0CAh3
xT14vBY5G3JR6ogIqYhkwR3q+RPYWCxcWnUY0Hr29NzmRxAr0qkt3b/6UoqOGTXN
XJtM0fNtjGlznefpzIzbQj9b6yBGFLWeYE88xT4RoFkoLNoZtdlfc06eakZ6Dd8M
+pMfAS3qoWMIoGO4PlgCP978G2ShgW52qZAXWZnz82Bh7HN1nCfWVGll+nMUI1qZ
VqOYDWO9WdY/syBjyzezV4UuypxPhZBmtBjUk2UX/n7M8TGl8WrF/pjLNH0Elgp8
4nJYjMHlJdS5Npgi4opuwrKVOuY2POAAEXU1vDCMRTLhPTuFD4nbRQ7uDqWegNoY
ZNrUPAPSooCtkpoV0slIJmb+JEO88QJ1puPii0GC5rIDvqjsaWCLOkStCgzwfENw
V8yCLcR53kJluwegry1HSm1P3VJ5AtQ7sS/4VALX3BpuwN1/IKbhh5iO+SbeT+JL
flUOQXHBmUyBzEw/zzBVgoRYmqW0Puyz81doLfADEw9n6y0ngQlpCEqT/nRBheiO
tbufWNzvExY1VD47X415LhqVMyshVS6iEc6D0avSHS5fpHxUeaECvsCgZRA+K2YJ
zaijPMkZEr/sGjd6D7sVywB1Cxm1M/jOciDH1b5hM2/ZPkGMLaytmmaGj++JiWhn
UWcy4hTDSHy+XosDrqznLLOGE5A1oNCrfnuZze36JEOt5G/nK26sTeQkjbbZU7DT
O5tATJqIAXA4dPmBwS/gI9wHEv18L8bA1SGIGqyked33YdHUQQHyO0kPTjJYuQJt
V8CJc2fqprLHulsguOAdRYNx85Ne19AbPR+yMhwx8437M1j0kphe8Ux83UvKttYX
pAEHWBiHqRXvjU74L30KF/V4Wu/nJsecd8bXQSjpjnYsIuiq2ksoX+bbwxc9IcLP
QckDrEc6UCVWiN4MKqy2ZTIOkyVbuhHU5080Id9APJdlh741dHD9PUvBI/fnSCP6
nm4GVN9MQa30VbdKpKz8LmhxnaEEfrmRoEMQDA9XWvbaLAFgkg/KHnk1hkvZZgRU
0YJdwkaUZh9zcUU1Pk7DFO0/ia1bs35EplUoFfceW0W1jfonmgmn133fSctX5U9B
9gGQQ0FWs9bpOG7uIikv3fSaEcy3KC6ub8ApP8776m9v/5Kwsv2LTpjNAoCW4hrV
wcdn8SHGxJ9zQgIz23ZDi+EIg1/EwA9kj3G9vQU1BMyyubqB/z1GCOSMp4hglU2d
I49xgF2LuOIUr5QqiqV2+06BCNwxNm6Rs/cksCTVcYA7ckv5X/2jKAy+Fnz2uo+J
HGpW5DeCvOVuULmSrDob17+oJWyagQXi3jLwojNh8wy4iWZxg8vdeID/OyC2WTAX
tuNMkJdMGd1tur6Eh+ACYi8Yan46D40cAujvTJXzHwYW4QyLEQ811xGJPVKEJ5L9
OCSwgzlgM5D83EubYpj/LP1q97hyiIpF4arErwsn401ap0A2rD3Pl1A4BeXoZKro
7jhSKNoxok4LQCWKvQKkpnoXa5dt/ZIhAKZi3v0+g1DByXbWYyEi4DqF1G8U8+Ok
pa5Bgb4jbTSW/qUzwEtDsLukBZ84rmKYiPqRAPwuX5UXcg1IEJYS7REgpnGngLvI
YpjlQfpRIHVOwoHJjbLjiuE5z+PJIkpocwb+Omi/3xrmQytxHod3m+S90wLghuRo
IJ1rVudWlN/3CQDpHdTvRJ7/oTAPlM/F0aHT8JUUrUT16g/Gcs0QrgUSNo+Kw1w0
jpvoE9egmJm2PzkOMtLAyV3Wy5Pqf4kCo0V4+TylBAfaPBaJbyv19PiB18L4nmKX
PnLGZxf40UuS99UQbR2PHqHEZK0jBuZdng7uR8rzMSw/rwBPeNUu2nFuimHl9MVo
PnoiiMfHslZwKQlks3EZKW652dLFZFYTowRgCtxsTO/3RHCora20MfE82qVoGYk0
jOmQMlmj7iWZVmEVP1N7fbbEb9s8Kp6sn6AjqpPZLAfL0T6juPnU6m4AxP1UT1Y+
HgcXmv35a3/K9wphM9rR0JXuIk/6I6gOK5h850/qPpeTvYkAbSzp8eLeAY/AxDe2
lVWGpZDFu/wvKtCjg9dejbcwzDoyCn9rsxW0T2krY5G1qxqk1KAQLRyXJ/Gz8CWq
FRTcn6Uv/mF681jIsWkWw1h0DnHpZIvyG0oKpoSa6o3FIxh+MyyoW7g22NXwwGGl
OYur6akxMc7v+QeOARx85jDTRLko5Sc6G+XSqDWCt17Ko6Glc8R+g2jhC5ZPL8Zb
yL2X0aEN6Gjlnu0MEEOVERLpj9ShGob80T3OeEtephft4+pjg1ZA/gFR3ae7lPIm
CmXjns+QfHhgY1gWsg/ZvhbCJpCevnLGlhBhfrh8lWJMbc8PCVDUDQoqfQdCTQuR
5n17iVRgZ8CGlG/joQySyaP/WH4i0qWvuIWxAAYRPa+vB6ogwF3YV3f2J/4o9d+U
lrKXHqno5BmE10V21z3IZ5IlJwQoElrzWZAABzjSNe0tzsDix8FoDUsCl6DQw6Tj
R625+jr4o07Ex6hX8+Sv6j83XwFCIEyy84xcVOQ7QjWwJ61BVYILEgzjfMlm6MqU
OG9GC9woUA4Mm2aqudJwQxaqq/0jWZn8kj1tPYiC+wOBa124PhUn7s/gLMbaNf3j
h8WVUZQs1HAjGK6860SKEovFyVb5BvaHD6GiL1w+oknDYwj129EOrF2Yf7R/bqoP
Jz22qA3jz2x/vsw13SCsjb/g2laalcYxUrw+4SJmBksk/63gNt+TMOZEez7WOHPp
LUGNIX+haFnzD23QvqufoQ==
`pragma protect end_protected
