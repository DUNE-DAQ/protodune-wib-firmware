// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
t1w8GUqnUjHaDJeYuu919HU2moX2I69+mpQWpoOfBRK1mfhZ/vXQxckiJUdcHWBS
VXJi0oDBN6Jf5rm/Vn6TlUthDKTQubobXBbu7vAR2tILjWVM4++dlQPUh3CxJuxM
nmEfXkDo/2NWK25CfOj2OtEAj8JjqbPH7jMCZzKrxzA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6944)
kQSd6RQ5LFR+1H6VzQNCFoDEaqmBWeOeGolGWHhj80vklLMIEUwktCLw5RczOxvR
sXaPI5M1vE/q7d4/5TmSVDOpwTUeetCX9HdWnQuyIkuDx88ny5XiHRWOUzG0Vd1u
2aFpQaBo+cKXRb6tr6p9nb7I0auA8SOSj1hsCdcYTMte6Dwik/SDIDormbN2Y4w3
gCLjIQ9VRrEcbh4HeScRRf4D3gC699+bYL4fTqc2TlYdiL1+S+RPOBs92a0HjXDq
yKKs6KkKtw8q0WP2yXCp2clMjQ6SVQRhVrvli1/dbTC3uKS302MknWI4TikbqCRn
RR6gxt4UxbGXUc5KIbbesaUrUth/1hJNpi4dByEgdFH5eIhLzOEWIy+QLkbAYTEQ
N1V4PIhLTRe2R37azh3j/mEI1WPDunebKdG/XxQzg6iAOp4+4DANaeC1WVGFB1OC
cghSVqHl7L+jpREyCCvGHjynOvEp6CiXPb4ejM0rdbYOUUCnfpvybeKuDVfDxDL6
UnHby2Bs2QgCQlp01UUdg5KgCKtoKIf6MP1BEx1Urur1RwggVC/JM6oH6ieb1K/g
9Z0nXvUu35j7/Nygd7wN3gWrGuC8w1UiKw4mfcBy76bGb1bb6+v2upgUVvvv9Duq
YzlcIimvbS5e+6qMCIbNZqMQTZcKo0gddSQKatpgovV8kcT3jtaY4oNR+gxXxnR2
VnU7eHKVtrNQxr7jdVlthsIsn/FTYXkUKTOcFOFRRL+8uiRaEZAurL99GaFn1cf/
PkRj9/tANAR+nuI/FtU9zxw5hOsyTQeTkQV2GwnyDjHgPVlytmec2ZQq27JNLa6w
hoCQ9PSDIwkyiFf90/KSIk8kPhE456Qvr+KSzQ+vHAiu+4ArgspGOxevJKv35DBo
5Ox08ztypvNEbSfzepnRGnRh2wQLHkU1+RscsC2WFWhJWv1CSSbxfsoHAA0UXZCv
OryXYAGHXJ8Kdn/UFWuAHB1eXFxZyfysWCD64w4nJyjvEfoamGbcIoAorgINZ1GW
NtZiW3kAc3ZhTDwK1sHxWKptJfonrGPsrYkN1iszugWY53I+T4BdDjNoxzAXAjCx
YUC7qs1ItOTgT6KlJKXpakKaLVOtC3t5unXR7dekJ38IWuAw1NqtVxqArFbBBJaS
8buUvV+4e45a20kHOGE1BlSJ4pTIwsrviuDuqJLHdy0ujk8PypczAoCWF6ULaHwE
FwwjGYllA1x/GytITo9N66HHw9OQASHztcP+YzH3oEupbQdsKN8eG6M0l80sd4pN
NwlCO0falB0PtrmuBLt8+r54AQWPrW+BKF2c2450PXO/MmhGBLNSYcF0AM7d4Q++
E63EsZRSfgsqBxvGYXRRIh9oDVzV/ZqFdlt1OqwIDzSul5avZMS98Ehn2+AmDUzt
hmp/NsgXfBskRubVDgU0iVsUTyIXAJG/6Oll3QU06PgELxGpvy2TlTN2AmN6pZKb
Bmb3ipqqg0KaHcgeh1ko47jZ3XL4L71Qk5SkCRnQkAgUCIbs84kk8Q5x5/e6ueaR
DbDoGzI7/+tAMC0ePWmRZRwy9vEpt9F3grlEzkDoOYzU3TDj1wc21aXMzx8z+diz
1w35s0TpoTwtCP3gCuP35vSVYE+/MDZOZ4UNtwOGZBE9LwJWVpKBOI/3OE6ISXxd
FGrTtso/WMdODjm9K+GbWpHc+lejiV+EuH8PyHqvjh+Gp/fHtbGZ++09y9X73wQG
NrzhFdW47UBNLxXwfSupLNVpCAq0MY4t3WgolOGuxBz+hvR+7gUqBxyuLJcrtNIU
bJ9g9rxDASWFKTRGsQnNM3ZhLDhvG7lXZeXPYmlG1hOCa0IYZ8GCP+8HVWmEFnxX
WPP/No5Gu0JGZUIupqeHb0nvcDpJDYBTfx9Y3kz9t55ti93kUraw/KCbI5WC8rhx
cCeqPccSbiKSyHaoeEn6RZgHNLFrHLGBaPyUfjYViU2+K7X0lB5XBp2MAJ5O8Bjc
duGGBTQBcvr9pYAAjXeULFP92OgfB5P39gEHcNv86JfSfxnqirpDGHzrk1ME/aXE
tz4vriU0QaOPTabAeFbrb+tslL//Tz7a2af8hlo3OJVa8kcuWbYmEU0L0OlHxT8F
gU/M1qbykRGlfA3W7VVSr8B4cXKlO74693eKKh///tUqxf4925SPSol6jzgO+edH
+vGS7Tw3SuLx50yEeQ9ojRGq0CiyZaWq2FW+h3n5t5kP2l7q7dKNRxJNeW3stgip
brT/Te2x3zkbPIAn6KvzxXBEkNczrqlzk2FyFiIRXqVRVarWv+yFwRk20ZRQOrmC
tdmOX91935+6AJESK/RTFcjiU9VgNN2Fy4Bm5d4O1eFALJIZrEn/3epQfdlE8vUD
qINmx4ql0mnI+tpR+qtzm7N4OdkgGZ2p4yUk76C5ie9uJQX4fqdS7mdSSB+Dxg6B
NG+j5x7sUkrEK1wivZ1EsegvZ1znVYzhOjk86f2+Q7Pe6Wwi+9xop3FIAcda63s9
laPHE/kRzhdLn3SvymITL6Vw5YYh4jg5bo8tnwkQNjxgHERYYf70SVxCGnZ6ri13
K/jymp1VftbC/goOdOiuu4fNlhpBOc96TlDtv4RwGnuqVt6Wm7FTvny2fe/i8TJd
nj4UeM+OZYQLDd75lqCYeL8BcAFmkapbXwZKYZvWrR0/kNzxNjH6gkoHQ3W1jzWB
OUz1SETcGYA3OFKymF2bFGYrl8cl1LMZs3u4dNPE/u6k1bfwL5HZ4Z4FImyhiV4v
INbZE4uUUorrwGQL2YqizPF1FnpT9lD3hFgS+Xz9wFz7PHw08V9xHBuVSTOL0Ryl
rQAIvg5D4FUV7D6VBgJzCHlv2VAJUi3gJGgXrJSHxYQPs+eT8OROFq9LASrtc+Sl
Iwgwox++yNNE6up2Ximcqx8L6UCnEO0C+rPyhhN/SrxRcF/+SrjlScx2zmYpKKVI
FZgoVNbsG95aA+UNiVKELjh5CS9YN5AzgE2dIBH08LXQu951fC9pXrbZirUeh7RN
R1VbWQP1ebX7u+HDl49HOOgJn4dhbMC4rOZgU+bDlPU2TwsmCBq13H1OqBYlolpQ
UyBF1C0LzjIEc9BSryNDLw/f4RDImOScYFB22A87Mh1mUW6fmO1LaYiFHPG/kp2M
C+3Z+rYpxRplxF8jonj0mw068XhfaoB+qxg3C1HB+C6IGA/PCA+idUp18AQk+mR/
snBdWRTCB9ZVlr1QHNXNN9uFcmeAD27nuKfC68XyylRvPMx5gxNnMkf3UIJ4W+39
T3GHu84q1O6hOeA6m+4h1hFP3ch5sKSeDRv5qt27HTAEVzD9+KUViCsopJtGyi5L
7s0aZIqqNTA5fBgfpphKBD0TAnv6wnSH3JTFDns/5P3JQ7zhf+3MYyeHXxAwUHH5
LVtuhVNTZrgPNEDEoq3Mm6eXKJEnyYY4EJ+M5ekDJ5d2ZkSRe9SDtC6KJ44Ii8t0
XHEL7A60sdX9hGyEM96n+RY8p9FWghXbLW37SSZZgMi+EIiJUAmmfgukJmUE5TBH
pnI/hpCVGHWtD687ujSun75L9HX0drrge7sASFKQk+66i7fpCuD7zKOzQLUhzgin
vITkA93jJD2yhvnd3TPIahqIJyc7WnlQKVbS4k1veUerBgO8Syr0EyGjUpQ4d0Va
d9H7dyQqnrlYzygi8JzYpeS0+GxR9uhHS/HbzqO9ZEPGZFHgLmorHnFgGyohqgab
nUe6d2MwC379ntTNujzdJurKVJYSzDtrZiL2Fyhbmvoru4+uZgbEjiUYiM9/Xjle
VVCv181ZjV0NCxMiOvBP5qVjnnlhZN6FoKg/9QU4CCeR8/PbHmoPFwZNw6NW5MzU
2r+Nvw6sTejjuctTloGd86Smsu9n6FC6/KxZhePuEmJHJSct70Zb0+RC9NkUKZem
d1D0OfscStzGl3P5HR0nX/paXUmHJyFZodpZvQS0O06OjhZSAhw6ki+h9SPfMzJz
Ni6RWNqfdwiovVzu0Ze3t/HkXzsWtXmmYNey1SCHTbByygcgHv92aDu2mXwqQVBm
fWg7BsUPdpWN1AoJe0B90H8ywUlAO+q336rQ182KVY352e2GtdMKqSjhr/fYOAcz
9Hmq/cM1scuMwrF47Hco9O5LtKxtAr/zXJAPI1y0xHfpCkszn31Y4TpREy3jM72W
fxOz6L/+8ZxooE/tHlDPBfyGOsG28Q0FJQAcaRVFWuh1Cle8dTAGkbS9uXSJB3mJ
k9tAj4uqXixIr/2taYiIeYGbSSY0ZfXpNrhUVR69SHo0oJldN/svX+jwOB+77bsI
JanlRbgfgdhIP4Vu5cpfOyQBxQxCMH2WzH3RCJvUlSmS9wzjW7O9/pGdrAfBxT8l
TeY2Dh6Em59ZAn/QOGnMcBp/1kA60bOlpd5vI8B0NjjMByM+IGJw2/ognpH2dBlC
ZqiPKMBtT9hW+6R4ZqGGtM1qwlvBqsKtXnm2vonqq9LOBCScxQwXC5GJpVoBU2YE
oU1UU5gIfnRTBPXD2QFUpKgErMl/hLq+wyYK/LzU+FrZnyvw1K5enLzjqeZ5coCz
OtwdE6mIR6614+jRsTAMQH0LcmK8s2UrwvR5os7WMyTxxqsMmz3oUOMHT7CtLf+H
MW6EIeSXvOK130c3//pqkB4B0aizAkiZWSdusmG+cAM+bzrBFKK204szT8xL3zt1
YHWlibRpxtrpHdFt6GKQUWT2jTVSG6S7puPWXWm76brKFQ1xFr07RcjbC/p4ZdMZ
VL+7zLHe0UqJtcVM8ndY8vJhb5TX1MrZ+TsDfmAp4esgw20E4dBuGcOuJWkKHHZt
eWdn0DhDYYQ4lhO347dA7RiaihpRuR1CPXLvd3//wzQaBHK94gAEsaZ6AG0CM8+n
Qz8CcsaEBSWL5guwBhgsIZYZhmImaaUkjk/auPKGo9n8y0NJ8BkFCQ00Imriqi+e
ZgSRIXAmIDTBUyWRdxMsHPXrDyJq+77nzhU9ZKz1Sq7MBNSe+DtdgITsIgollH7g
PRjblJohhetJJFB0DRxfKJvrCIBSvQhBXxLs00INiN+lT1CbzQba7kh2vIGm9Hzj
66CXHFkwFUvUBOkVVCNOVIX/EFvBCNU7CG6kZJATchUVbuqPDWLGGnOs9Ffv5Y9P
/N0PEdBPFmKjjARtTEp1rwxgl7ajEmQKeL+uJBBS2ZpelWXfCLwcjntwjkg25Enp
s6C0Lk14Lzof/8pNL9DRrHaLYpZWnIpNvDvN/xhcNJ+wWWNM/eKziBjAJLGs5Q3J
loDuX2DwH9veMoexrg1ijUDiBmNWUqEvuayHlTzGk1ET+i78NYNT8MG01sUqAS+r
SF6jm1nWKMRg3yJVsvXnsNNljC8NKRKXh+lmk7UAv848GieZn2vxqDfh2I/8jeGK
7ZtXMFHzW5Nd5rmHR0euoBVFG7aSMho/SeEur/obmFLZn7cxQuleQYE2yiN6a7uY
XIfsKd46VG6ncNluLFZEdZfDP0Aekh+6Dk69/9wLJnN9JugMf1FARKiIv4dZg1IJ
Pjr2n7Mr5cxZWGna5E9rCkycd7vp8fuaLaJdGTDApqhXNx+aoo7NM/oO/bFWja3F
ffvp9bchN1T1YOl0kRnC6xMDQ37b3MAzSyWImtBkfF+gKYoAUjnOBGaf926rqCSB
mytyhylly6NSp/LW6tRXErLAFA3AEm5QG01zaqnHg5BsdybqO5RRDApmj3r/EZ7B
IQuAYVC6KLKsVBP03v6yRM8qRkH25qXQjVUqFF8lLRKfa5YxIBT+9c8xhovmYFhz
p//0GfVx/W3QxopEnkew/g2p44TZy5Reb9kaMliW9C+pMxnbjzP8fzkGBwpd1ngb
l9sRfXToH/OCSx0cYVO699QZMtxJOYs+C50afFpa5dex2tg0afQ/TASbvA2NWrqy
RYy2PkPkgt3PDeFhChj6yUmV1CvJiGaSiFbOzb/Ma+CkXAPVv0DPJrAsQBmaSqCc
HpiEh0SVbrBxFEge5CE55Q8AbZGQBMVlbF2fliI2Luj6sd3noiYwYCuApdzal/NX
6C/DyZ3lDjoZogzuXbDQUc2jILOhJSHL3mZSqbSOioGlseXlT/zQHKVh144UvAb2
UdPzqWZYN/KmaK9iRnfyun/mex44IeDjJ7TqrOHOD9NTJJsFj4TYLo6dj6K8uFRH
gHl5MIqB9917oTeMO8rkwXD8NsWA5hYtYtaeKklM3pHOkLtnf+iwKrOcI2WmPy3n
0rpeVzOP3qXdLKvMg/9qeeNRpbSLNKPP3twjsLUvSNXOPkxgIZFRoKt8w7ATQK6r
2FDcTLPVS27gtBGafTx2VZtfyWgjLC65d/puZ18Qqr/MUrG9x0zWBxgsawGuzZjR
v+vQGog9TZd2DiDhh6e+/2mRqlet3qtqEjhDAwD0w4K3KYi9bDnzrvtDRvc6SU+J
vxFZCsgPUu/lk+u9pBj3TELPZV6aJmfI+Rx31AefxK9Cj/aefk5kDBReNJqc+j0n
tCeQa0eWV79mKxxEGbadrxnCtpCkp056p2GXyarMAdVw9LoT/nWqHPfblD4IWXMP
BlYSpG+N8ABsNv4cglbGlKlxeLETNINYDAiV9RORMJKgnyGSqDZ20DsyJ5yQrOBb
11Kwea81p2R+8rAh1coj2NhheHDR5RaZHNSsDNgYfujBKCfoKAJA2s2js1vlnN0t
R1dAmahPupR15zeRkaz28/ZYOkpDaysI/5bQZ8KX/S3E9lNBr0nyVE708HN4dOd2
EGxHMgovQC/qcph8hkR0l6rF6ScLLXFO6Do5pl87CN8WHK6kInmldNREDt3Ww30f
BsI9eqyEnHiMxqX5FjXSExdRdtGqHhWSuXgPbBd3yJ8XjeAEmVucFFdVSARf6rN2
dPlQhu9vrbjxpQE898apsUVsbkkCAzYudLCNAyei6QpXS3z11TRER+AcAOrzNfLk
VnmFinTkVdEZwTBeX+7zLNE2SM7/EvcLUHGyiWBXxeY7hKx4Wij6WmekFJxTSvO/
WNBz+l97VZlwbw+0zVqg46Swb2cPelncu4AKKqM1t63eYgiqIELk0JuZCzObBVrr
NN+QQWc5LXd15qJPJLttsYrYQWn3Pp8JwV93zIkVWCJ0javI7z38+gCRuB1Tg76a
BDpWnq8gHGjfD19HLaqAC92/JpM6y2gSVSzvahDqYD9kwMyk4zKT55BT/0LG2uQd
6TNJiPnJZpJOKPwyfyGsa6VUKAlrw3BfBv1V+JMotGNNNCuUNavlOLh8mzaYUKdC
V+ofQdDwd44D/UY98By0T9+0ve5FvmtXJQ2WVOn3HJSk2qGB6NUPmO9Uyzcee/+n
PCbgp6/Sb8ckQGOvElVaeQ2otSny9NGT0gGUEhBunaavdh499wPXjmbMdReHcIED
/CiO8FdC3t2isphOdtxstkURI4F2llS8Jo7MgtcaZB/pVAW27Nr/NIJwtuFds89W
0KW7nl8blPNT904YM/Kq6T3eFiyxeqAHVLOojpq/v9aP59b6tnUdHh57lU43inFx
nK4y/4PoH1HbQ5wVqsFAerK4sb/0JAiPbaT9E4Kzi0KQU1avrMm/M8BbzplIGNWh
oVgAJwzr4QlgqkHbqictUvpJ+hmtPv5d4iCCs8+ZaYpK4KYpu1ncOJE6ib+ugtLI
9Nd71xUt/symkpo1UXshFkFUUXgVTgDMpFnXOLYbgQTh9z5jftwXJCEBewJ4DbTJ
n7FQtctZEcxgGv4KQ89hJwjuHh0ZZbw2kQyxf5SyauuXA0rHmjyTb9O7XXl2MQZH
TXTU3gBXTyOHpvLDG47oXXYfg4OPRbsmg4kV3I86aFINddUXSteewOCVu0+Iv3NM
ITqKipWBMqNimE3Fx940ZaqoljFXNOymda/Ges1aI/wZ2dlcHDk7Plvb/ptmmzDI
hiLtUmgxTVNPvmw4zchFBUPK7sr+MU6CVnGCRxFobLddA0yhPdWR35G79CIGQIiM
ZqgUpCoy/FgdzaMWVBbsc81Uov9vFToLXEW6NBjgPeoABNm5YtOd+zRR9PBKiqso
W8nm78Fd8JzIUjxOmMTL1Rv7/8BW/qGfBxn4B3CZG63PRAzauwnjlvGM3yZNkyzK
JgEmLy1oCs8AZ/CcCzUe8ZOP3Eg1Y3m2A9RXL2ttM6a/HcEnD+4hH2/Qd8w3QhIL
Gkc8YeQWbdIlQH0E8Tw5lzVJvfzL0dcqOq+O7uyRQZe7Jzsn4eIpouAyRkJmRrHh
uuT0/tfX2dZVzxKapqb4Gglms68dqxw0zsl8e3XOBqPmfJHb1kLSm27T25DHCC0Y
IbxQ15FYw+Md5eAHkyw+5fyYR8jNP5y1TP4MWu6vZEClhZ3VFRAJ7xh5fArt2eo4
eMEvKfbMsn4nftrvZOqzOt++kS5zLFa5hetVoleriTKm9q3fpLje3whYZfvFYD2W
/xWJhkXHW26rIQYYW2TRXPEiEW+K6BCCPuJQLvpK68X3bMpMAL8OYoidqxJ32bnC
pXqZ3Svx1N4WfzIXQattNhs8B0mmx5AZ6QnI0eDNmyvjcMuh7hL4/HMg+6ER055O
4llp963yZReiiKokTKq/foaZVWtKYbWYdDunl0Wg0jF9Vv64RfuTHWjliRVz4YRs
NITdpzw4H9fd4DoSUjYedzc7S0POU8IEihkKAc3SRg6CEui+jSgnGVHFs3D3/dtJ
iokCc4PEKxp6Ml/za5S/+jEAQYFj0QxWtPztYu0OouBB8RGRxzQahDDG2RvCpLOM
NWEyeGPpIhIQmMqDWqSSalg9L5e0HcHZ5WLnC/1hBDXM01UX0XgeffVvzoe4qMVR
mvEsZn4TiGDjyknGbaIjLABjeF/TputXZUhCxway0CAii6lXlxqJQhmHQDlWqkMw
NG/6uzNzS5y91R87oVoNMYQ8KGwBhmj/CWB/WbPIq9bSPqloxF6y6CWN18ZxBMwd
MyGYvOF53jQ8222LCcpln1xnSXG1rA6/mNEY3TSeMiKa9GNs93NENl0qVxo9kZx2
g2GgDHk4LknuC2qP1/x+k5k/v4etYb3B3/0ktOBYaS7IjUpX8J2nl3DMvremirzH
mkfNuLBowzQ7HRozZ8OMqcgjPzGzcMnuQZ+uNtFfZ7xHFeu7qRwSc7n/A+vbmHKV
6wdT3dy0DdpGxI0qdHmlb0Ae+xiLchqKCNCt2HcMH8q/SlqMzYnSGTN/nOjB9CaR
4skJwZjTndK9z7MkJLIgXDHZ/KsDo7Vhyp2+/9JUAu34Co9MSHj8v72IvRssbev+
6CZ5ZyNdZyC1KCRB0i/j+Gs23MsLpANCMQ9iIcH2J2Y=
`pragma protect end_protected
