// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eyNEkJ9/k5WoXao9bC7foNqvUcerOcfXYjYxAJmnPuhL/cmKwPPL3d5f+dUjLfSa
ZyEsOAunSempCdJ69d+Ei8gWXO8lOimyI6eBmd4QW652Sbvd2kTEn0RwurwzdBuy
XLmQNlpfjcwaCNeX6J/klIdDLZWXRVYymG9fKwvivkg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 103456)
NOiVcV9hr02G/d71OYFaYtNLRsqXb3WT0ShYEf3agNMHa/jS/1USqfQ7ADRaUXiO
M778rmIxbCxLzZfKsT8/z/ZjKhfdU9Uc49xrvH/5OPx8DUNV1ez28FhZOFjAXwGR
Vz89P/84+O0OgrGRdGmuqF+UleVsTg427RxbH1YeJvROKoDVJW+w0ys7BjU+gQ4r
GZt0WjORvl60YODW7wBZWsTmixvO7z3YvGzeaIwoJ4hIvo5FJVv8t9Q3+1N90o3O
IVXBKiOYKlLW1FIjbzSmN9xNNHiKliuYg0+uFH8aP52FTiS/+owvlq7g0BJCWf0D
xzXXmxa2KWPY84pN1klh8WdMdLyPetUoij6yEJwv6eitMuVdf90u6o+xP3rIXxEm
oAjbPEJbypAuiteivd27YS0F0Po4LAZCSr2YcJu5GvzPDUbGCAPYeUhzHVWeo9OP
YdimzrmIeHHWZtdzCL58Tb/sAP5RSf6hVi/Av9sFYOqZ7+8r5KJL/4nalseOPp0A
1xA4Thkn7+NYUbOZcf/kx7I+kDpo78bhPvIveHgk/Cd6UTYG/QZL8obXgGhObIsg
Tsq56tDZ9CUt4+8/pyK17xz1FyvmSEK5Lof6YgMFLWB1lVLgNgFO9QSMUu1qrAn1
eBV6sbUUsq+40Ht6iXt7GySGRtV9ouLgNwyFDpx5/5lrHgSiPhmbx3QdohRHQPie
M3CAO/2XnBGbuaaIplPHecp1zX5WHpP4V2AAIo6tfeYZIzvXGPDH6XxiOmzKdqta
5uBrs01oqIHzqHOIdjG/AzMq/S4I07SKpsQRlw3tGVvKZbS9Hcdh27/PcO9EruQk
tzWPXmdCvHbsaogQuS5PUSn4Hbm9Z4aDXst99fSIUriGW1Z3KtPVdvk4YvH7fACB
SGOrvcY9SWg/MbRfJRdzoaDtfQuCnSKLhmW+7jlj1p2U2VljZU/3heAGNU3GOanh
XIuugYNNlMCCYZwpYwJrHUk168J0va3URY++tcFJK8rU++zFQ8+0Dp8i3tHwkjvk
nkbFxpPGrwR6xG66LYy6yipHuwcbJQxbmE0YAqYTbSqXEeNIEp5AFsQYvak5SKKs
oHInnKKaNyRxeeARkr1mH9lMDY/sc0D8jPw1lIaZKxzrKH9Y2AXFV0Zlh/bkLwsC
P8rJgzezWjyRKYN7pGG6ULL5oL3Pfqc5+PFPUQHu/3NRWhdZ896jGhEzKH08UkNf
xkVZWT16adzfmmOhFZ20sez3zHnUHpyyilWbDvbAbt77eTyo41mfNAyPkRveZDie
QTiKayEoqMR/enrOiNJtlcX1uqjRmLlQWBE8a+dzYOJbxPc4PN7GMGDQo0q0Fq9p
ylr5V4ddwiBc9uVgvbI+FY2N6O4FTYb0JPVpuKqVNU4GPCmzWlRq94Cq9klV4nfd
kFaiH8QwWub25A+titnkJX0EBapWrBO8niZW8fU8iCvEve1PGm/Uhqq00yPl5mZa
VH2+xXL1jpBC2EVU3JutUftMM0PBp/LVTB4rjV0lbfq1r6QJHd1NvpB1SMCQ+tkK
0o2ZQ87k6i9QdrQMyjsmZuZlk9YvIFAKDsQG9ZzLgCZ7qajByQ+g4DzC9G1LLgUt
JBCqkzA3enTOqrAxTTetXNNGTfi6DQpgf7/5fHkwE4Qy/psuT8GEJdTRKNWzBbmm
lt5d2AaQ+jbSpjGVizsH9lTmy0aTs/hrv+cG3oYPBYLw9G5cpPNrIS7+TktooTQ2
J4UsaKqqpsm3WmHGblkv7EsMtetrRcyeEy6QWUn9d2nHlEGFXO38kVDuPKLGtpFl
/k31ek/B6awwe3hs5u3MXhGr42AnHIvcq1KYJOeMvoW6rohRVeEhF9hO7YfGdaGv
k4bptcmiaOgkif5w13QYsK+Da4SrRACCMY6KHPMlPhFWFjSMiKjVg8z8bbGVGRjH
rrJnFXhTzOFqE+fYu8JfkfswJ1WK5NLFcMOZSzHZeKW+wCVQXHbDFePOS6cjZ+2B
B0yydAWNeNYoxlNqwxBW55dJkOaibsS2jQSaxJ6mMk1XOp07SIRju8K8qucna9R5
XtRL3H1CFovQruvZ1n3kunxRGDwdt8LIg+gN9z986Y/9nU6yh12gaHeWfhd8bTXb
YM7104R33DWkBFLe7LMMpG86+Ldc08tlGcggmVPxnqAJmRnUdV1DMNUjjAa0BUNJ
g/MocImc3Uchc9RKmklRBiIxNesyWIjCX3lEvM45f40Cxu81++rvTq/uU5k4DmWV
VrQY/vNz5PiaadW4++l/Ja8t7KY0haJXmg0NSFh55DTMkP8B/T/QFACLWI3+whu5
v3dKx4gTOhG7ahi7Yxg26XtcQfFqKs7VcclZ5BVP7eHiBYf7Eu6WcxdVRzb9rneD
3WRbs03xjHbrf/eCcmLla9+sJrucsLm/hJp61kbOi1u4mQIZ6Uu3kbTuvZffkFLz
zWsNRLaSAbn6mCCBJvOYZifSzDKNf9OFSVLy/bKwoZOyqFzUJaIbGqZMMXzlzAQ+
TSXOAnd6QDgaQ/4b6g+60qi/8H97rrq+id6R47dwAIFWs/EOpNxf+0ykLlqdi4hZ
F7r7AL9S6bkGL2M8oD1xucIjhwP1FEEg3WHU3gXoB08SY4V4PXiahLv3Kmo90fAb
PDEspJ0SufkcmAL/0PPljK8nd2RoHKATjkJGjnXvqMjARiHhcCQ9PyY5nWxho4aK
nUVNoBRaWINWMHP75N6QT5jgiF8SXoj0qwEdL+HF64t8xzqqJy7oHT9bfbkeOtfQ
bQgXHpFZJ1BuT+ejTFYU3JrGGsxIyg2ELUoocrD1YcPkpH8y8bBEeMoOcTotHQhP
BYnBPfMrspKg3ieG8tgxagOPay5W7vyk/NDcaEuU4m9jhsqngkjv+SEGm7ezxs4y
l+Kq/Vo4DDpFPedVrZ9Qm9w7vB7mQxL8V/0VKP9UqTcUlkDW77b1v4icybVf+Qcz
qn+y/euaqoVe1fAWr3E181SZ6wXROULZP/JRW5QWVedqpM5gzNACaWb5M/O8e4kM
Z0x+5a6qdm2pZAJ2lNHbgOTZqSaNVgeMeiHfzdKmosLKe77v1A8o9gSi3O/v0HeR
Tkkbc3zWWheckCtqo42fzXbZy7r8S16iAAuD0kPgntRcimFveAkVOsP/50OCBUmS
+JZzHaB7q7RnJpCrZ+Hz7Zr8bMJth84y7HeJ7QRBD8dhMAXrAvUj+X4Wfd/raL56
Z86lR50Cy9UZAx7ghFhvUrLpfm3fZDMusxSN5+oXGx9yD0zGaPWJy0eO6sw4HKBH
y6AsgC6h6rzcr8xDmgdjpTc7dtmFEsf7mctZ5dSU4KgctQQvMSb0NjVGz0/k7H13
gJPzSUNETqS0Pi0Y1rqqtUVjF4tKir+ZlZ2QPQx406wa+b0jbXEgflY8ostpSpHs
ECo5OcuF5UBpns043MbZxJ83OnhjXzPiN0fkJUzA+Mackx1+fARZEngRmnJLMzQj
3xu3kgjUmucurr7ltsasWD59F0twuUz4qw761XLkVdVAnYn2hLfu25ThFdoAcOTw
HD95BfBM0QX8715febM/9t3WURX1CD87wnccpHiCxtqQaHg62LpPOXEAvQ9rDO3o
g1wRWmtnBrbseeZ0M2mK2rhS9A9ak+B8tPJcYp++43Nz8ySwLTGNDMCTnVsuA4VS
QuSK2n0DIbaSBysNTeshqemF6oHiAnj27jWdQYOGVo7Hg41dGbwFeDdUgSkIvijO
WyUywUim5z84zZxe9uGejGh+14uML0cakr0F3tkhJc1Q5vUA9JCyHGFiiSjsuNY2
wVH7UcxIu381/YQRu5u8JFZPp9GmfbqdGtXnLx4AhimT3RrK/n7vBQpwESOD1j3v
fS7XCfc7QBDJgpksDlGtUFzYw/N/7HUjA+3K+A4N7sFnL8gESXzEQquRrB+b1EWk
XFop7Kv8JYezowpOyZFGqSO3xAh99MTCkk6VuIbZPh8I+kppi7JVaRKYUuN1JSXQ
OyIupoJ1DndovupllDezaTVbgBuz0GQgQz4CIcsp2J3BHGiKJPC2Z0r13VaDg5LK
jf+d0Nl5lwwd+4quYK9jJWPucjsuZf1GL2H/+k0x2dCYPxvjrpyRl5TJx8z6Ti5z
nFInu0Myp+Fq2CxSddpLg8MsRm3qkVHrNbCNOvwL6wP8t240qV8/vYJRqISv/6QV
WK56zlqfIpEQVOfsIYg5tV7M0lFZf56YzgNH0tPnnM8aHa1NjltE0ytJeIw4Ojbn
Pb7ovGhv46JLC6MTHFoFDzwgjquJD9fMrt6N+a/P2IOsdO9iTwYUnptm8vlZj/jy
tZbTDrnkouxIvwbADkXNsiTvq1o703w7z7M3zoqGMgwp/LDvpqPSM6aa2w71wzJ3
H9rOgjXuAQL9lsDjELn92g3jvXHKZHxbrFpqaF+HCKAtpRy63qdQObzne2gONF9a
YQFQMjYc4qcRioFfNZ0vvfa71Ov5jgJfPEJPO3A184kSYnJKGfY9S6H0D/BA8CZL
XghYQDNosTSNMoGV3Xjt5SCYEePrYWdOApp7UEOwafhS55yEF+eYq3iI5qliTlDA
YlereZDWfDBZS/4dp4cKpK+JYB46WHGxucVP6GYJrnRQ4tXbn2gPIeFze0LcVu+r
3I9mAkJn5nJ61zLYWjF3mnjuSax5AmPfLBfLISTgTxHI9wk3RjLgW5+sIKsAfERD
gPQHCXIcy50T7KaysX8SAcEsTO2N7Ay3SDU93Hhvarp2DJ/Jrf6r1PoaNjByATfb
qCzntHQGxzHtXoxxBEZim+RrEqCSmShM6qb2fy8zUezc7Ok+7/D22tUApoXFALwX
+b+kx4ri1/+Xm9wg3V5uhEuaJBrGZtP4axH335hJtddLnvAmA7YlHq68+giEekof
tnWNc/j4Js0eaJi1NU4F42ydRb1CgP0edGyAqnWhKnuGNQXQxMyuGsPkLXjFHqBN
E+3grkT7bnXSDgGxvWiiKjR7+oL6vD+iA4yNuy7Vb1rI3eymgLT+/qilm9+EtINb
ZUAJwkmWYf7puJKaAlXRe4sxU79fDVHBklD+w5KaMr2maybMvvU03j4fcMFVwMzX
xKKqoEgEPZE5Ca11tUmsNDJU0pjx1NyQaNsA8zLW4b2dff+on211cxpQA9z3p0NT
qg4UgwLL2LyEU4e6Q8VLCwJyZC5u3nTB4yxBxs6cxjZNieNeV+aDLKh27UseRJGZ
Wf42mtvE0XessnjX8Y0CR0IK1ab+sGfncPkqjEZMjow9NPF5I+H8Zitra6CLkhle
opwvCNwTIhJ8nAqnw5OxP7aZ8s6t4DdFhljC4MuffrznCe4DelDIbqL9BPN+Jh1W
tE5VV8N6VC2b4tYGBs+mRYP05YMNN3de0vUDCUNGeNPpa5fhBBMBjUb0QZaAqXHj
TKwQwWTyEF0tNWoBBNsgbWiYL/+WTNOtKheiz0/XNk8nZ3iI9rWv2IpsqPV2oTjv
K8CuHONv4jFk3RtCuoExqDL2lrkZhMq0ZKyEBtp4XmrdkOeVG46nVouDu92TDwS4
FKvhGU0/Q3vwRVVzzHzkp4gViMco7Yx96WL7IdUyTc3F1gJ0x6vLkR1tmIV+BhIr
1t7jBHpu9bsLc2sNBPs8yQ3LxCj1Yr8N/ZgHYU2hP/H6rW1n7WpzHhZpdXRrPm3E
VgXlLeZ0pzwvhsqzyySWaYBCQH/gJRq6SwubC9opqgYF9oqd3emyMG/Dy1s3TkSX
T1NVqGrMyjkOz3D7ROBK29Jc5yG79h/NNVJG36iMeVNcbdaNuvnipXsLP79QaM/H
Df7Oz5Mrnz0c6FY3Cl4Mp1B80PmXIfjSpShEDMnalsRSZdlRzuifUmQYatFlefMs
uoVvqVXCX6Pdt6+fd/9gMOC/XBZqh4kbMvHntwsk6ZbVmynsd1xn83AG/BKb7Tyt
W64qd8DN0EmuuqVJ8n9sz9UZTzc9CyLVgwbsLLI8uV/3xOC3Ig6fIabcSR8iUeU5
S9ml5Owt3exsMejt0zFuj3I2Jybrny5I1aIfA2lwjnr3uSa2zi8c0pGWx+YHxobM
0n3TSdGTelaWzoWkRpqAuUSlxHGpNAsKb1K3hwZk8N06Fr1b5wc+n0LYAOru8/gF
4kqvfHpiIEZfNwWog/GB+4wr59Y3IIUXnt8oXDgBDztWLnSzrhbJ0FZ2xZqgi74D
lAJCO/RXhFM+qkPDP5wDdXOKX+osM6w4F7Nvs/gKN3UW2D13WuhqJjTizO27/5BI
v0wlU8vDZQrLse7i3r1WG0/5jOsA4EiaegHaZ7WioNEL2V4PniKIMCvYoES3JtXP
69w/Qm5AEYW8vDiaBkUaH/vjmGL17eW4FHlyOXM0GhW2MpvFXZV5dSwVt2AZ4kcy
WNNdqJ/g0NHmHgHVA6TGR+XABVimtGmAoejZd22ymeStO9P0y1yAHpBFge2cUvv4
s31ZrDfeMu2yRxaplMsZcTQfFnslZsVVqqwa/JXDoSqLihCVQUtuCTiyjL48gGdD
UEMrCyx7dDig/JgPHgNySkx/JXccGiGHQ1UbC7IRnHMYP2tsNhHJw9UFoycLoZHQ
eD9V928D7+QvY2m9rMVCZumPdupqedVK4IS0wCP5fW3iwz6hJEM1O6sldtAa0WJH
aV3HpwPpaLzWeNsGoorFri4KBC4s70uuc1kfdsAzb0/wj0l5R86ua4DVJKuvHJyG
xtFeqH4NY85QHcy/emYFIIqOg+ZAcaWgyh9gLKfVdPFQ8jGWBV3Kip/uJF/M7UTI
TJmv6NZ3bzDQDFtKlGjKHkgUxJo3s94+ZRgcO0XyP9KK30Uz34THx7GiEyHrefPk
4GcfXGQAx31LJUF2yCuMwKC6Hiv6cySu2rA0eMVgLBvG9KuU5NdiMrSRDsqOt0s8
Qjk/swWuBoG1hg8njPi5z1Vtz9Cg60HZA3LfZUNMK3T8Ma7Ce3aG8znyl5coQBXo
daczcJzn1OtwVdmUX7vKGuiuFqSwsftIYCQqA7qFpfptgGQMGFgO1ZHFC94FYDs/
erbZHfR1OndY/dlZLXgH4yyULyo2BLnYALcmzKl1U+15QIkMikRF+JIl7UMt7eWZ
IbUEAjfHBm+0DLssp2T0T7mJRFU7B4I6p7PgzBOC2Xm1PhfYRFX5KBIOvXB+eVcM
mvqnL2+2qUFmE1VqMpwFuzBBhFm0taPH2s1EHf4iWZRRDpB7QUrL3709sjCKN2Vk
vGml3ZLtVzvEFsGJ2HyE7z2q15F9OOG7q8hJVRPTN5Hw0JAfi92C6LYK2ZFmb97f
EaddeDhYBXiTxH1tErAAR4lAupqh5fYYFroqPAtbnkz2QW6tueIxLbkYnPfuVOUY
N6MXiX1hcpTi+jlfteMvKCduIg9vuK7qQbkxqnqXFeaq1wL1+aQX9Wdf+Znij+Jy
Las9WgDUJTIHBskMJL2XaXgBgR1PPjtqCv5escWnxqjRzVpSgrO+pE6nZf6HUc19
SDSYi1DSyTYBoVphbdjzoRv4bth/pXGLHN2tnv5AEBQlcLL/1u6dGlt/R8JI+Gn+
uscKa+1zUnksT+9/TvuGYT0TKmUMhRL8YIIisk7zqkBAYbktMGxtx7I9n2njq1av
8WH5VuOalMnihsHwGbB2tGn9O3tRi5hnGP4+IjG+pim9GpAr++QHmVgtjUsLWv8C
dsp7lUH1qzI6KyJFnd1MhIqDsCUzgBcTmLMduvimRw+Z4hEng2Pg9V5jI4sduChH
p+IViZecpjOjUZdLle5ML5XBdo6MUG6enexQ5SlYLMECKWz+XoG0ola4b6WB8Rau
EHt5NdHrgg7T7kENjvxyNU9KkrbIB2z6ZGbOKjjwPfEP9Xb1oyWAq3BbLjKEG6rN
7PwurK81/agUzFdD90frsoFanAveWeli9HI1rxl6SMuo8abDsBcjz0tai5yz91Fs
cBG0wsdQ8O+oUwgPK2Un95rNGtcJlZ+XYGg6O7ViPYmqtk/fXQPYC/OWVPvQjGAJ
3fI1YYcuJPeQ1zWPCRnsITODOvBztYzuAjKBqJQ+fdUXQQ8tJskATEji+S0z4m0A
PNChfy0NBluEHGfg0pk5qdEcOY5VfC5IA7vpUeWN6jm/M0ihkDRpkgLn6TXyYIjp
+c7kgDun0+mITeaTF1yiWl6vmCKnDFlWJU3MBQD6b5z9pzjmhpRId48ta3XavsIB
9USPiI5WeKzaxbbZIdspwddcsflSbFp8+P1hKnxMFeRY+B+l5hKCzOsJ6CKV38BY
hzGKeywhhzPAIV03XqmW58aqukJQGTKf3ZpFC1Mcp4m2Rw8t/ekFlL28Jh4I8YgW
xLCjhWzIKdEan8iUtszb3AGfNkiuXMdzIcv5cOXmNjvpnOQHZSg9Kkmom0T924EH
Rv8n7VTfT0kcJPZnnOJKxLQ1ryQILx2uVcPI21om5GPf9pKEZzp86MJOzs6NgzWx
DyfMk73Swzub91E9ZwtHc2YJJoUOuW3ZEtZUbG8QP1EQRnwfl9+rBxVMnoUZZKED
27+Fj/vhej5zNIGpnabTlvCKE4Uda6jf7ZgKD4+85P8bhtXWoGAYo15fBdu+jUI2
8UBUvexVcdDyPlUVEwBPflIv3T7EgKQUJCGvJlx7ESV9eeXr5kO5yuCppjT3aPM4
i7ziNhv2jNJZONbKN1zkWUAv/gsG8Ud/I6n2pthCLnpikl5JuXW1XNfOUh9bpA3J
wX12SU3OONP3J9TogR1kWktvolRdQVPT0zIPe6+cStnZDKlKrlq/8DV2q3VKwVCL
HXaL0tjbNv6KsiweW0maAHJfT4eKgrfbYLxjA/NVgyDH/owIY5kbkPNLOs60QGp1
dT+g7RHnP1uvwApFy7Nx7x6M7zwnqBms6gY7OoEeZNNry4mu8H1mRl+PIX2gbuyq
aBEXPJ7yWWvf5fX4FsKjct2ZRAvEWkDAnYxPltGnHr5hqSeSTVhNW3Ten1MKmFEN
C0i9QD4IYH1xuM1fuTFfJnIMhhCrQdlAxS7MnjAoTIokTt3JluhOb4X0Nd7EsnaK
AmClBu0A843izdOvBV8Tj2bGv11BCd+zqyJXC+uOOTPKx/XZibYjYkKRAMwJbGIB
JQKEF8/n/NCEb58ckY0ZOY9K3Q7erRxDwmP08IrtyyGUrIBptnd5RD/25qDpLUiS
MuVmFw/mKXOys2RPCgrdyOkqIZQkfoErj2IIZq89cnnKx4ERNWEbOAW1/MLwpveR
lNP6qBYHGkvXodknoRrMSY7M9+/q+PTHpuYsgAwNW8cHU8GAQtWKrZ/F2pEbFOCC
b/g1lxehdNP8yEVHXV86o6O+tiH9kNRr6syhxR6naudKiYBZh2fI9HATmNuifFg3
eqOFGQbRgmmDfnxd0undzVNlcpS/0nAqHVcmb8JOR0IYf5fSg86+jChXPZ1rhDEw
RZqCa8WWNU+o8bDT2NeBamizS1QvbKQ3kLc+zGwqT5BdJxSO9Cgke+lbnbez2QTB
E7AXmY0KaNyHAPgeXUvyAopQWvnyEGQQgckWb6cK+FmK+VtzPQy6k87hcVBC3rNJ
nZ4QS8p7DRTbjWNhXCDSiG+Ay2DoV5WFK7udlzncaMVf4EIRWnHaaDJyJ8zUgSoV
cjMpCYVrUWceNbmbYawWW8gXfCaEdYwE9aMGUgDLwEdkxuuF9JgqxMqCratOsoMW
VutfCi0SNwxAOAtNBjrZECDf+mTItP/DXg59DKfXMxz48CTeMI/klaKDHP3zPiTy
+0F8LHCgJAnxUAIOuV9Raaf0F9R7OXHBKOcnlU+SuC+qtrfik07kJG6rRxbwZ5iw
h79Iavv0xVLdqsgkMlDYxyAy9VoKJhjASekMfSp6t/FRRF89MqTbaHAz6kFmHJIH
2cJnG0O5bp7UG37C5krJ0UmgMzbNoi5lARzogY6layWRQp3vuokqbPp/4eTUngBN
xOCHMul0Jb+iwzijsgYDOdpvMpnDDCjH0iRAkJRENPXEtMOKAp6sd9Lg7KG+Jte7
BsPccFwGOzkCgkrhCO/LMuTM58pxBA1or3ZAeZ/7VkOncwjgo0byOI6Ln0W/cXi0
fQq7bXYoiHnkb/yohSUkG0MGfEnI1xzAEsgwcRk4FA8UyXBw6zYoDN+SnQgNuWyN
58J4m+rV45Rvx47Ul6ZmpYCm6ti5DQ3RcbeGAK1I3Qj6u6/r17YXQp5EyZrCzHBM
puGShhpxLRkRJeYbxAf9KanYXlKZWLz+crzWX355Vo6TGYqZ+GcaV7UNEoE8JMlf
I8BmCC3EcACzUZvXsuyLqPZkIuxjvhUGDBe/S+bfvneF6z49+59YqNYYZEoUSpjy
NU5wAFROJEyv5LEHbFr8iN3nYiyYX29p8BWTsz8soFlVDCBabuxPHkyrQw4LGBY7
5VxL7L/oe5DPATAyDFVZK4a2hPCnzzSeeKgpYNJuwzBwItmIuc1ocvS2p1nme9T0
Bi3wr3ihVaz+USKstP44Bu5YbNMDyDaPuAczmDFbi42m5ySZWimVDyNLmzmxQAKX
1F4aw042GEGRIoNKm4qdrhEjIKvUpPP+J1Gs0hlVPMe0aK2Dr3/GulseDpsTaspR
vEO1fzRO8kl81/FGFsKpZ6QSM8+WVT4q3o0Aye1rPfNZ1bttctPUNp/fiIqKnkT0
xAavf2u1rTwUURuRqMFclscjzqvC/yzqgK2topr8/JH/N1uSdGU6yyxjqunRFQhF
4vuMkc7zuy3GjOGJo5YQycpHsuTPhKL8BMMbpNCkyVXVtuw5otVNC7hcLh/KBkmg
Nk5zKgF1cQljPVWvncJ9aHCzLRi8h+QrSin9TYVPyxxh1sFE3zwxEQZDaQTMC3mX
pUPSjjXtswc3WN22SVfixMdFAKiPp5QaZbYar7HTir2GszLtLtn7P40/RR1jocJ5
x1XlFV4QG+EEyvcHjwt7YRMSH85m9jWwJrSE3C/K5MmADwi1iCsKNXc+pG+KAD3j
dN1NvHxSN0BNrHD59t6q0b4fO8vmtXWk9MpVd/dn+Jgp0TcGZ0G8V0df/39gvEJz
fUXitglC7c/86UY4rKiVI4MCrtmegPPU1YK089ftfd/ZsZXNOBs3PcWKzzPhqVYL
9ynC1mPaWMgVwaKqXfVQiiRBpeJ1H4ycZB5d9+OF9vn/8mby4RIVCSHM7KOygKh6
ktU2BxZLoWAKJ8XndBX8/+APfvHJR8Urp0lMyW/0XTuqKvDXiT9ZeCbRf7xZN+RL
wesvCrzEMuVfJbmrcN02Et3oYUViBNDUmokrl98W3VznkIXUgyXh5YXau6ZPTdud
bYcBkeWsPbuXGC4SVhGRggNMFVv0GwIGNiRNPD7+5tD8JQBuXhuxMGa9mvcfAQVI
2fe8ntgdHWxaai7y2keEOTgFb6uHDZM+/guW1S3lsu9xVBLwkpBSbHoohusTy7Kn
mTE15VdI2iGeGwewtiRMKiUZgIzdnWO+uAx0aRkLMNq4AkXK36hJ14bQsBeW2SHt
HEhuX/nmX1e+XGPNm6Ru+kvOpRVw/WkeDBQUskY5znf984HjIo/L5U5mC/kF4mJJ
zrKDxyz79hoDGWfwOKctj41Rz0g8CT9q0N7n8ad1hWPjVFYXNdkeU5o2Jk1XqHDj
hwRMmkokFh/mckqXzP3JkWJUf7pzM/+55BaPlLF71Igv5vMMYpgeK9BjZ151NCOR
5kMWXEG+8/0+APCewmmBjQA1tJE4d1G4ek59MJB8TmHxll36dxv0NF3CZFRI4yXh
OMSU7D9SvDUSDdn8M7rpabKQDuP5GmrxGbExF+5eYNCSnJ0O/TiTJ7lkRupQpuZD
On4DE+U4vDZoFR2nwfQ1RANXfhTpnf75EBaGiKy/lXO+ENvJIbHBmLQQYgZmoahw
v1AC9ezWwZYWWsak9FINaD0Q5w/KBIJlhYs5G155sRE8uMcAHhz6kxellJbWNjBb
lT9+hE/c0gAKhz33zFRcMed13Dis1JDsNXAj42rqeroVYuMuWfCpkTNpT497qqw6
XT6TLdgyQW1bnBsUV8Rhvu6nV5cHjzOuVA1zyefw7c97EylDoA0tgbpPF8xBvM78
FvjJlz6wejZ/FCwyhEZBm7duPg0XPqyWMPHBaN8JvM5tfb27ZdWbUfjWp9SoADsR
qAHbzjT4VYgR6jLIFLOS2m1O/LR5SKesxu1XLPIvMw1QedDt73D6pyfclN3ZcLyO
lVFKqqnqrbpqnntN9U/6dwv0UiYnt1w72fLJxM7oHPpPuuKn3CIYMxNm7GDdYbNI
IjzZngKwFGBNQ/b/29yl9M/KahR7eRpLmpiVZmYciebUGzuBO8/0JETWHk/8eX6u
NQMES4Jleq+Eyo1xWu54++WYOE5nKUJc4iT446WbCpygNAzQLouzFrEVNG0a4pXh
80QcGQxx0cTw0Ewy6mCFlHdjHFoXmt8vAKUxCdHuKly9YKhqQDxU+Hu7uHvf6Jeq
FiACkPbmUB4ThFjIXHZGFuEqoBq3FySDoeSS3keL7LeFUkLMWJyMSsonHpPEvCbz
rdkF9rIS25C/UGqNkLHepcUT+82Id9lvL5MdN1Zwfm80vIYXguT/2rCJD4sX7jkf
ABJtmpKSpJDe2kkQsVnXnO+QnB1LLkJPj86xA2agLlhaZxXrHS5JWqQVZKJw6hHX
JBFN+VxuxhqJcocd0IjbvzJycTh0K92nOatDN3Pm1VflpNDbMM7BrdRQaiAK7z6D
JCH2EExDJD3udDoXZzjDr8TSXeGLxUbWxonCNtoGDk7VIGVL56FVDb8+EzI6TrNo
2LIL4i6tx7lCLoKwzcAwzGOBrLeivptMcPsxTwewwOHcGBwcnaxJf6jUiUFm+f0k
B/2M0eYBt2gj7SO8cZY+o4pQbKYy5turWWRbTpnRGxnkLlbowTIIfWhyaDwAhc0q
+V4Kxizu0wBvq13XTvqoD0cw8RwqOf9pFOWvd3rUi/gHD7eAizOsriWSICgNsDQ2
/iQpk2IZxzdjLfeLhY6l4EILxFt891KkVZB85NBgSOInf0Xp5SohubjOlZY/F4vH
2XCZc9gY2Vos0g0xIUELOQkw31UGF2RsB+OQXZ9jNvRmWpEU231qCAr0574TVvcc
F2uxcGmAF5d5kCis9p43YJOGJla8FWs70b/91kvUrRQ83LHCH+VluI7NSrw2Nnw3
d7Rwz9tY0KTX7b7WPJo7TUYDiBq11n7mzg/Dd0eGPKAuQvkIU+bA/bMbbBhoivAT
eVB370m2pc4jIzlHSvkgL2TSLwv5Yl7K5ojtGZpmSnwUYAUqJAi6wp6pRhXNNudc
rFRuip2/60wxR6FL3NWhUXEBRAlQH+ZVPciPPyMHVONWdl41D1vGAhcB4UUyVpgQ
fSg/kUpNwi+pFxsLMYWTWgdUItdDns+pdddL6I7U1SoTV/fh3HVB0WLv/bo0ziwu
/Fq0Y574icC2lZry7qxABoWQzl+C5R4lBim19yaj6zaZxmVgBOK0uMTAmQ7iwCFt
Yl+tBOeWJTSLTv/ZDiMQGLovHdHoP/L3YFf4ZQIL704faxXmnBncmKlWDMv2FU33
F2Xmh5vdaRy4kI2i5SFkaB1JSZ7axzDBrMeORtbOOiQbK+0uJnx4IYCtDL7kvse3
VGbY6Tm5tq4QDHGjtpMGwNxUDH8lmt4wZ+seq4ck9zPw4mhSHRs+4iYRvsvhv0fE
YRjYZFPyXV2gxmZT7WCgQM37EYIOc8nakU5Kt/6oeWZkB1WMr5FvWVHnY62VSmCJ
aKpcF1sy2uKd30m2ZWnEUFT53d0oKLAtFSHOAQUE2peRLqNigZAfiOAvxsXAkC3I
OMAVpfATGRwP/ykdV+tXgyyrVp1pyaLvG1ElgubF2baoYTE6xgVzxndfVXgXnXBw
46mZMP594KHkOVnCrTOuA6+a/Osu0RE1LronS1zUtj6vCTrO2X7P4Kd05H4oStjf
UoxWGpmPJUGv/DZMql+F3jWHs+eXgGAVBxgkSGq7Va9sAA7endvwZAonz1reugF4
rMVY2V6+9LCc3BoqBSxqoIQ8+FlV05domL5HyLHGsMkkYtq3mhPvs4DcGjHpNdvK
VaQqU3nNW64N0hW69WxdY4bR9ED3GVgzf4xfjL6mSGbR/CJ/NZkynko5kUoQ6BIy
3ji3NqBzfXyicKQAj98o0uIhdKnLNr7GEpx0Szq+/KH5DEoi++hMro7hInsKYKPh
tO9SAKimiZQqOWretfBhsr68qB/0egzK5TleCAPSKxvGP8ITmenYQPtZfqT3qxng
DCagOHaLf2FzKlpc0WH07WrNJTRX5CtR6ru+VWII/k2wem8VyYYeBj3noWGnRfjh
UsDFY7wiuNM9hhKAu442JZAOtLJcYZ0ym57t51WuqgeFUdVevlQJ91qHvip4sgzW
X61niDKHy3UBeZN5JovzKhN3JakepqRkato0trFXUpO0IoDibxDX177DXUOehBx8
bzxlTQAnz/BxrCtMQldlIMaL9FefMzLWW809VQMkgE/CMQrVcLI+cGPhoA48yC4Y
9furEXZyp46lLk+ND4OY+pLx7ElYO1P3gb+nBa92oKPobVVEgFrt0mZqEqF5gAKx
TBlT3IB3a/1K0eW+HG4j7Qq8bRsycHJ2t1ypvyZpF31wyjM/ZUIJABADRZfnkWyK
nvauiipXximYhNMho7wZK9kfmC1YbO7OEDkC4CZos6zZmXUtIHNfIBa3xkuBnF/Z
ZF5hd/qO6OMk4eAfAEZ2GIiTdgFC3wpEXnS3mFC70v/W44EbnHCv11CliEn46fm5
jzPaPLp0N5Wu5k2+Ys51ODdjbIR5AyrgXn68sjj0H+TuF3ZKVTuNzKgkqzHDsaQj
rrLmThXRCh5023PyPtJBAjReCeIAItBla/hONnxawMMYQClkfUVHwjvDohk97Jrz
NO4dE6BMfypnWfnuAW63x+XYd+f/4eCNsCPIpuqheJUq5rpo5DHtQyKg1s2LUEOd
Rdu7Ot/PToTvc0BqZSTtdJRda/SbBHViuxybsf6A+otYYLOUUnQJapReEmk+VHjz
wfn2Ht+2UhaTtDCQA4HW/JrHcQC3qhligfC7m7yedKhukn1rhSdfRA1aJ/Lnoltd
7RgW5RWdvqMDTfaaY8+fIgh9BQmhAAOUEWuOec5Jjqf4RZJj9Gyxn1kk6ZBgR+5P
M+uWafnqBPL/Oce+DC8T06opBKXy9no+ptT/GgoCpI9EBBIpKZK16d3yR5CKw3q7
o92e/S8mhssQCE7WwJtxgYOPTQaQMaLEMx+IswBNGGCrpXQkk/UAdjmxPJGIdayH
0PlqFaGbz79lu7/CwKygB+q14azxarl8BDsHoAJLY3QiokDSEJY2HbJDlKOtHFHA
1GRpXYEsm/7Dg/tKJNytIl+1ji9rxkW+f4JL8/pS5EYQJM6csRvJVb2ifxcmP/p2
nvvyNiXeU2HSQPX7PZOP58nr8GQ9wg3WH5YTK14YHzms72fAh7xNXlAQrpiEQp69
y457qhToKGtAh5chqKRcXwJDUd6/91PpgD9800t1E4W2Cq3uDETF1zkPM/4zxqZP
k4NtSOkNBgo1rvSt0PDlqvz1eo1hmLwGA5smvw9uIPetw8o3WVx4ChoZwLpRmTg1
XR2UGxFAeTi2La3dNEEuVEX2PWpKqkZ0ndDt8nPmpXLvoXXI+aDhXMeR2oc+mm59
dUsv1pfyqgFRGW674d5gUjH3ig2f5MvO2NI6CGrFckGv7FYCl1xYiDcC1d/ffyqW
zPEOonn5W3Ymyl4K6vz9wlVZSdjBf1eiA0sWX4gHFb/JNe7kXq8uOtR4naivGz+5
CtuW1XN4nZlpEsWlhaajFzuhmLVySLCxxdA+6y9/8Y49zjIS10J/Lf8YtXyuY10C
a1Hj+s4lqDPwd9d3cxPYhVRHN13BAnIDxhV/vvvl4waW4dEDKHRinV6YHOk5GH3u
Bs1NTC8BptsJo7yHyjwBVtxExTcX0FLelxdHtoIbvR5JL6a64V3iNUPoJgfvp8E3
oJ7elVUuOj3/9FDpz6ksmIb+UL+EN3iGq+iDHEs7wxf5QOO3PVDf5msv8ERjaAzZ
wtw6YfFVsIvmYBMwGq4ZmuktOyXUoYJZYCJZW8tvZ5yomNbaSpZTIpB7vvcayGil
ZBoap2Jp59mjAKTolIqd1mgFz2dnZivRM9wUpEwk4oW8pCG9vz6S1+Id1Ft56aG/
x9X0VgJQ6oRfGnAzwIFyc5fa7znDB4cuV4sNS0MKDIUwMAsY6jFhTlUDUh35jHUz
Ugtf9Aq+n+OBnMq4P6uvVcdIGNQs9hik7w+80G8tqqbEsJmiRnMpVdkQyGulydiN
ZIMyPgXRKc0E5GoltMNQo4l7vyA33QSTLT0Zbg6VvU4yLjWTkiDI9jChSXJPwr9F
oRhTEwCDKFc1VrgNSSCbP9BjKCEng6TSM1Yq1AIidqqXTGhJjsblzK9BdUo2GVFN
Wyq7LRVm6kO+EDX2vc4Avv05GV2CUsFZYWtreQz+BGlAt/Nx9yw75Q9aG/vmS6Xy
v5VN9aQspZSPfgfv+nbM4FgMkkxBUp2tRci+NqNWMTdQGooLLQgLG6k27fonavSB
2GNYs01WUVtrSr19AuXoGFZSGu4U0HRKxGzXGdhfwkvkqBfW3ypYySRms1bPhLiP
e+5uXNeN8w29dFvdCmvUt9hSPR7nAbmyeqcoILdNqoW0UMff4lCk7bHdnM0Y+Tpg
JtYBRKU2rb2YER16hrylSTZWKxNt3sBRuZwJ6AM3YHixXCfkRaE/AbAqwGJiv+nN
trbrXemVE/wAZ9rzgXFuVekr78ZBpeMudwDiEZwQJ9nBP91W2Ai4PaAWJAyeyXEP
t6NX604FL05+EGpvxbueJiW8UsvEYmGoMjTTauUCVYPeDQLY8PnuZYTAvfcF7XmN
vL6jobx2hZurb2sWTTawn/D/fVISO+00Gl68wZLxm8yzVU0O+IVwn5dA5ep5lJCH
mB+Ph7pfMsp3SmyEgzRO771QF+FhHDadFmQ8Z8KSct1IJxjBTUZqZsCGhTOSJMQT
U7HzsFjHsEuwl+3j6EGznDKyTakJ5PD+tUAf+jCnxiaZCGQ/xhA5xyiP7SC43YrW
/9vFTJFAUOg/zZBzwRBj3GTkIvmvVjw1K7JRwQ2+BKtB++VKdZ9XgW6UPHNiszDZ
IczENtz8CwCZFpETTWhUiKuYflnQ4qGBMJD+M3okkj61WAozCli6JXmL1t8FIIJo
WBjlf/Km9J3NhqDm+AI3YlZDqMeq1opVSlJ8JQtntiYe/dXOsKJUx+BVevdbcHja
B8Xd0J9+pGqoKMujtbwT83wvHahYWtSU69EPziUSwRR0osN2I/a9PKoioesbF3xV
oHn3mGQTXPLp44lEvaUq6VrtWtuQOJQbs7jAJXGUX0wbtUKxcD9pbj5KhaUWVkxY
jwhl4bxzjQtSKlz8Fx724t5NgD8lmnxngoRPjv7qspDsa/R/rloPhgEB4E8Djl9h
lc5jm8t0jCpjiBGr5ctOSHTD5i0fzqmCxLCggHcU8lTUoSVm3dGHRnelX8DcPn1N
KKtDA3CUz3c39Dk5knqq4+SvS5PsNaKmfM6bakeMoFiNmp4wUZtZNmDRqPnx0Mr9
Wi2J0LFsoO9cSuXwT4ehs1tpG+MXgWFC4rjFD/N6d/+SotBVVxKTP5OPvEcWcxD/
k4Yo2ZaNnbdsMlneVeS+4gxDKb8FhURD+nNIgQcZ9WjJHv87DjKhYqjePL4JDz0w
TLedaoN84M5H1nGtjeHbpEKQlGm9M+Tp3oEN7pX7gSt0032uIa4kW5AqmuQ8REnz
5I1EGzeMrHSVyKrsTRRgmcFCbYFmwtZXl/vyyrd/N0sr41yacAigOVnuBE4KtFTx
jyzidceQyMAwZi9/Ca++lbmDqBK0OCr5P/e+RCZsJUt4qEeQizkspOwoAL3FEGcW
tXQ4TMxtTjhPXx9GWhR0jE646aiD/6Sp7epbLbs+NZtiWcv2miQ3yswvgmfmq4LU
+b9tFlGIgT4qgfITQ4aFCNavLSFPw8jbRrXqwnXITK7oNcEmyZXzyOfk6mbsj1+L
+aUSQ8NaGHuC5WHnHFEoPlE7iH427Bb0ICcCk3JnyTHJJ2/RZO6aWS1/58cHfocI
4uZjuPZQFSWpQ34L3W+/qSvtJ+iL0QnOr7NqBpOLE7ujAOsknQxMNrapHTtNXFwv
nGTajifkMyKctgzSNiFV4/FW6nQitGxc2A+ATIhSOSXH91qK0wk5or7E3HUrh/Iq
a2Pt/FCDfmLGQy0FhCGHyoXM67OxNV2Iqz2bLtQgJoH1tQlbeShOoN+Hz0p90nYQ
iVW2o7hHQPNtCu/biYeOIo38w7w1pGgfrnxVZxN0t92VTKvPf9kiNeh22lDfpyqL
NiBG/efIKF5InCqEgci2ajSPFkeIk+pF1DVOlq5s2f5sCZcPLZOySOyKygNsoLC1
MeV/TNH/PTI8hACIX8AdOdHnupv9ErSe71pWPixKSXyzWvEBn3IpVBEShSJ+vEma
kwFl91KWOaNZBDxkuasWsO4g5aFVAnVh7tVAZwNu86JBpHGzJo4paiVBkYcRG/9L
qDbcxpPMnme8sHmvVzuezTLQkqi+w4QCydCvgsSRM5uZ0whTC2qjEe9QSSv9sIuI
DqDJgboPNtzFdnbycVFJPN5oYZ5AUoWu56U2+ukvn15lLiNpFk8zE27vs3Xmm8Rq
ek99oRl7RUSKqitJ8tCo+NPMF0lkveSHY7ei0jhR9SwVBLAw10KCxhAo+bicMT1J
W3qSoEzFrZAcxYVCCqk4momO9duw7TOGbSRymsMMmR4yOwXK75+Di1EsG2fvxUua
AnApED8dHZDWV8s5FFNqWAGGUWq/dcHejzj0YUlF+3SIpbMR/loMHsmTCZl4m654
YmDI+eplwElNzBLW8cPUF6wRHI/lKJTLgDGJMJTBpsBJtwa4VlKX93uzgM0v+CeQ
bjQ69leWY8NMVq0xmxK43MKe63lqg7XKPSYowLQq1RYqn+JsQkjPfG2w6r56PIPc
A/jc4gie6UZA4KHZQq7e/dkkS+qeM+5bf3cbGbJkrkDkgFQ8SG4I5kVFDhgcRY3N
00g29WBo9O3Cwv1+ZZj0/i3dZFbqMl+EOAxOvz8YaeBil2F7HVK4waYr7Nse6L/W
QhDJhMDzEsv4VGt/UnaSl6Gop+3OvEbPKP9DzTOBnWLF6UD8f4ttjggmypYEXVWT
6GQUCG+F7NSYQrdoctB8058MVasgCVTDqypazTNs5+Fz2cIhm3b3FkITDbB/pMJq
bZlumOSlpvibFsRD8V8ZFMsqRhU5CASBtT04TGi35hT5AgNvyUMukzNbT1zOQ4G/
xpXHoZ5VsB+iATZVJ7hSLkl+2a9u3BhXvBEvpanmtWybrlqoUnDCUsXZU3brcu3r
UBvhlLM8cHkdii2hmAQo6uzG6mOjxBb70AcufpG3uhJyV/BHX96AeH8TQ3hSikjH
c30+XWCQWQJ8UAjN+s92INHeiiLSZRa2MflaaGRfHYfCFj8eRU8uc4CNR9eQa8y8
QqKH5zBfJgRWQlWpg9/Wva5fS1QS7EoGQ02HF8dHN0pE9ec/3vG58RxJTeZ7+3At
ILtFnDnMLYswLlh0WrAvNPxrJwziQDN+iAl9yDP7pOD88KhKlydldBPcpEWJgNo6
GFGzoomwPfwdQXbf0yW4P+HXOGVgf8CKbntt3cHeKYy8roQPt6B29dGf7tn63Eoy
NN0eQdsI3tpy0oLN26ik0KAYy79p+Xtq8Cmi/2PuSG/BFwiuIenGUMJhUFE4KIBL
wDsCHCEH4ZwQUs18fe6c8HCbX1A3sPbewgcs7LtznlYyLO/4jQqjR6SI4NLbMLT2
GkegTo5hwzlkvBX+snY8V5pzR+N5Im0E/uPrRdlzFqGBVeBTfu0egX8yHVzCRzLx
umQ0WsdIC2GdfyHvwlCuiMTCWTI+JIziI+V41sGwvJFK5ckZT3qk1Mh2LWCz00CU
JWCn6CVJOcxidsOzXEC3KPvp4Gig+VO8+q59pNItsFH/l8ZTH5axwQjQuJF/3snw
SJSIuGeuXDuOpqV+CVV+BJeT/CfgvPy3NQD+EZEK6J6vLB5z7emoRbTsUmEAP3cE
Smc1PXkw7llYkrYU4pWLbZU1NKE5WR81JWWHhBZh7kEVsxXQAlt9OkxrRCD3Emdv
8Dt/5spjiVdHFFIb1rmiOTOLURi6cqRNoha3SFVe0o18OILXeNIwnkrtVLTMLfiu
mx0LwQUUQdUsulu/AWfKXKzd5/VCxHDh0mEplwYRJaC+/7njadLdXJsxTRCJI3H4
bj36vESlZc4hETpTgl6MywBld8mGhBo7XjW8csWovGJ6SUgJz3LbpGZdmvzA+ow0
ysB7hzIXHMtVNjTd3bV7B/zbB3Ol3oQ59FbKpXbZwBX7u4CfE9725ORwpv/RfHD8
EIUktORg5+YGO3s0Tj4Ho+sDw/UWqyOGJ7zfD6I7pg9fu7xV5sY8tT6RiF+Yd6W6
Hf8SnMCvb4X/gQbolBDM4K7cDBmk8wgnRCiDEeBeDuKb2iiy9OXSecb8a9XGpeOc
Ir+ypbpi7LSCpL8Q9uIC5Y78PoWY0m9OnnnDyiZ95wk5+z6ix4ZlOg7SQ+mAx6Ki
ppmpJ+Q95VT228x+3Ic42gUnf9YP4yN6A5x7UvCipiXRjNdUK26QCOcaG5ExdYIh
YU427wXA9vTOdCQL+hOMOjxfhxmj9YqYYWn/96pn3dezXZiZQJ4Vh/N9otZ9BrJg
pVVr3dfsyYJmR/f3EEcQBHQ3vUfCRflL/PmC3xeNEs8ubGPaYD1ACm2yuDnvBBxL
FgjpBS8DrNx60v05nOb9E/jmRin4G8NaBYbEX3zU4kpygFwA7Jttnq6g7K8AReFN
mHTJeN1hbVHwH4rYfh8+f97b2BqO/cIXURIULlvXNiFSZXM/MU3LfLB8+tnTqaED
wOmxq7J4qGeFMSFCC+ggMTXmkNyDRUlG8pWwsQwBe5LdnC6XpQZHuJzM7IE1RJAh
UpjuYhfmNHBuinh6Kjb4bZVg6uOr8PK1m2mPkMQqzV5Vfv/pVaGKSCRO4LrofTVr
toVhXL114yDzgOIYmlAHct5bGSMSk3P0R95fHpaBjNUPYbqknUkrci+GVDEAwg0M
Tz7EpwZs+TRvzX/eGc/I/km1b19iAGOTggtnhMqAbiR9sZk0IDOtG3CzvLtnQQ+w
EFto4SDdEHN+IXvxFEw6sRsAh7RyH5nxUxUjufsAcMycK1SKVC5a/j8ubwmqw1UC
Dbs6QpUb2Ap6iGRl4jpuNjNurdPCzed8qXSD6NGb1Bt/yT6+iMV044aMyV0n2+A8
qFAngCTrVZIPZeYZpHY28l8H+yH2ACZkyFay0R8otPxN9OL5Z5/8zFCLeU5FIuxO
As+Imi+5pn/hr/txOszqon7mkSPKxWIoX93WyHDg8WOesnqLXSr909wU4g+8dnAW
tq2GjglBcPrr1OeWA+vN33ti7OKi5uRlBchmK0vhsreT2NRuA3GC4OUyHQz4Mavo
zR2XRCuzFhwrTsDshz5fjromDA4J319sH86FCFDwrETISVTDuFCnQeWX+akfD2tp
CeUk6K7TLAO+MpaBEpTcFRKEbH8NhjoZcOD5FRgN/k3dDZT6spLTNSXiVFiN0Mch
weqEjgce6o9GJH7ZhzjWJDQsXB3bFeuBzFkqLrm4R7Ba3UlbhpVVVjZjOuLbKpFV
egwUZQpaA3jy3EscK0o3FAiXUiitYRv+E9f8EifdKLDZPrjVkmmfW6YADyELxFO/
XSFoocUgjqrSqPNm0Bmq5C78StKgC/aw6vLhUHL+EaCofXNdO1exK4hp+y67kiLP
UF8EPqWCh3Z+xGfkh41e9GJfxPHIQqGdg7HrOZy4WJgSEclQFwsaUMlQ9G9tX8KW
LpzGu1WJbgCAcpZQr25y2KNCIYCuwsG4IAg8SJyTuiDZBZsvU4env43o22faJouI
YfzAJCRyXI+1ZHBitb3CB+3gIiRhJ9MFBokvUK/gs4jcSIgEvUTvlZt2Gh2sDEWC
fJ1Q8mbUdfukvsSBv3pwphxo4kWFJzF1OryUHOX+7plGGQQB8zRK8ELcF27w4GJ2
zobG/sSakuGmo4yKnv7C/PnlbbT+ZZUTERkdJfQf9Iia5FwL/yzgdsN3Khq9A5dI
tE7QtLd+1h6RbL69cUxROigyuDAGvCSgL5k5ofWOzm95a2Cy5FTW7GGxdJQ6i1SC
a2cJIVaAQDTkyv9RqGcVtWBTq35rFiE7phCQ3rT+sAuzJ5uDGhRPsSTC3r3Apbdr
4AQGxyVmB6+noHXwh8gioavuPjZuwVRoCVlDYTAqcYogI34MNmxG/+/IWu0xyX2I
1u37aOm6zjAQENK3yitbM7gmS3rQdwFYGHzYb4YM3/SloSrxAYArozY0HbCR4o7j
RvA08Whh1a7X3rGYhRmlUQOCd2AYxSPKw1zQ9tLfm7q/soVktFXyR/0pLEtprkOu
p5HA8BBRUZngz4FxbNmQvlhHVaJRO+CAuzl2ZQJ6e13+DLoOKY83Tw3z7PVp+k+j
X4YKWZbc5CWTDo708qjBj5VrIQV4CnRxswQDXqW2u+m7KnY20ifjpl+j2fXFPgzg
k0gXtZH6Ot9YAiJBrjXecx3+QEOmS4VvzaCxOJ8BmuHEhtOpWZr89pEA945M3Eat
/b5SRxQddREcGfFNRWgAK29u24HYcODSFhqxXeOI3rRy8Y3FFWP+ti8vmR0mOGS7
CzQhg3nLzU8Yk0TrDvfB7L1vqsdsVMY6TBRtwSeBQr0Quw4cDhpue1MnGnsxLqJ/
aMkf2vezCumQ2LStkVhAERVpQO661L1bNmDET0bIG96J5G2dgzyKTsGuW36vJ3wF
s++2BASgL6EVTSN6+4P0U46jqy00omzfn8j2CrCUjgoIxLMSXjYlHqt6SpJWaTrT
C3x4w5WZah3HKjSk0ua+DeeUZq3T/4Qx9qqfMNrn600IdP2v/7OK9In35Bhc3cJQ
V4XcwA39aDNTaOlNaaptXuGKt+TF7G5SpwHsUK+u4ZgLlhWVArF2MvPCyk4t/5FL
cAwHbM3J+qQ6XIIMRkGAFw4r5fxGDFWWJLynv9ArcKt4HSqTvVA2P7z7nH92Tl/c
YUixxQwDyTSdEsPtpGeg13saKcGStlOz420tA/UiyAA/JWWsekkZetZpfNLo+ZgH
NtFceuAPTSllr+idJsaA3Mu0pYemBuBWD4WxDGTY7MX9ysHXyEZxaEvLIKL+SfDb
krrMg2NHf2Xkg3r+QUvpeNvdx5zyq1nUWGAVj9c/h4+9QzVZupMfT3IHZzSi87iS
XCdTkgCWHE771xiQ2lW9/eAr8IHNM50wPdBnf7z6FnVooKLUWRm6e8uUHWIYlWnp
OVSXp7yFboblkYbNjrbxrcoXFXn5rEY2tXlT5YazyKoSKdZAawknxGXRl2StxX2G
ZrktTNtvmUMFsoXzWz6EG3UFjZYFMEj0AsSZjItyni2KXRtKa73tWDNspeXfYt0p
W5IOVBJdzSCfXMnlxzY+1qIcK2Zo1UcRQ83+D3fkghlRvym6XVfkv1qu+q5xzrTl
65u88A7iV7j6flvA8pdc1iSwXY7Iwxyec0wx5pAuJNV0942giVcaRTvI0RoT/04s
TQ6l0OkTQa9k/QAWkHinR4bYlele9j3KIxhM5i0eA6P6cNIwteoB5gWiadbr+utN
+CnzOLV5K2XcRxhInQkHsANb0Y7GUXzGgOjljUlJjiOjda4xbQZkuTBbF8qtfIHE
FK/e78uNI1iKZRssPadh5fxpMOWoR6Ib2q5ThVUGj4dBCLdp8XKl+T9IKTiV4eZf
xxpO9MqTJkozftnQ7M1Md1kl93N2mzYr535eikZ1FeQm4jbJ8jlmuCJinxCitlfh
A9HOQehg5TQq6cnly8wlaAC2fCJaTtsxfymnGA84uGS5siV4NfGgC8hcU6FuJRjy
4jCpa80fj+mk36QTx80zOUloZzwk7G1gwuDXQ3KV2Zkbsb1V/2p3liS3VwKEWgHF
JdK1TcxD9vuxWoFcXYP9gbjAB9hcpNwSMjd89xJaDnzQiFiY+C2FW7GlUnfChFah
+7Vn9+HuJU8Jh2C0H7HIiJMHyw/nes+X4xQSFVvsvc4ZfNI7kKxwY2620z9CJW0f
DhcebaaAkUZOzRww7QPU/uON9JTIsDSIEj5Q7O4OzQCeNwCT/1HZLPkx3iGKvZRG
XG9zgsqemDXzj2KwciRN74q7sS+t87uarjTRM7Rd78pwF7q6W4sB6jSn/UGJgC6h
7JoOz6u/CQoxIeaGi8E/rWUA9Unp1o5Okw3i50RNFk/BmK4QowMfylfnsbx/kPUf
Gm33Ms9p5TXBRKvHJJJgYybV0Bc3ibvzVhXHh1tAtICFCLe4ec6H5U/UuYouG2Qp
KfTD8B1g/I/AyMSVoMTbBhibzjMbJXl0ZUUDXmZGo2B2BqundcejA7/4DAGwg9RU
E4R2CQi+uCmT6PucQtSS1kNoQaKF4taiIJF8xhBShzoWINzCxOKFOj1I6Zcb9rr/
bACwnfJctI+nYbMTyRg/ouuGCYsqG3XE9CcI3MyTVEwBuRngryPOLkYxkCXNXizH
h35kr3nW4dPuNunNmN6E4Bu22x9nzUOy7zaIeIHJzY4K5ZraPHL47JsP4CjR1BU4
3fjBVcR67jPyyIAnIdbAEQdD9o6Csa5fKFYcvkNT8CCqPTRcuuCZ+seZSrnS9qFz
miYw3YhzhBce1xWFq9C6z0mkXxoWSG2kw0iX7ZnY40kB5eYs74xoFOidhnuFgJew
Hx73OjcV7+yUTOS8vhCN8u+48qGHwg1YEvjxxyJ4Dj9LdK6Np4jGNtSQXiUX85Aa
CfKFrOZR8MREBqiChNwcp1WVkmDwa8EcNfZCNZ+zUotnEVt8ZoAwWOJiTjz8JzLU
tg/cU4eMyhYFs8AwWsPPsu6yajvQKd9IvmVK5z0M7rBmD/2f4iZV9zNX/Qf4VBuo
SpDOxbVuuPAcNwel9lmOXxcTHPRiwrQxfQp3nEJzgy8ihb2zjFgDeveQzxJJieB8
xX9CeBp0Y8YMWLid+JtqW86ZNlmxFHamFwbYJeSDzWvn+6oC/fxDMunrMDuZp2vC
Gfu04agNOwuiE+E3A053jRkEkK/drC8GGJIqDlcYTgLr1yb2/mpQKvFW7hKbAvwK
DangSel8RcAlCkA9AFCtW4q5J756aRgezSbwK+NHfEMGvAsWbkUVu6A47NSF7Pqr
s9kQEyIsRHtpq+C7VvrWlbT3yv6Im8MBOOFZ8rRzt0YF+jedIm9UVIQwWr8d7EqZ
teVsiTULHtzoqHfk6krWpK/tO4wVxoP6SBHmlr0PkcZp93XbAVhGGCjw+78quY6b
v8DtVtuOx2F8KrVANBx1WyiDKvDMaBDFLHb+JaNmCWW360wQkQu0MCDJzp/op2xL
23HowuXDtyryHk4qWn16ulYj4n1t7erkyo/3mSlQ8bHbbB/tgZG7G020S+w9shQ1
Wnd5opN4KJLNpfYgh6O74JnEtqQ3bjps02XQN+IJn4uPB4w2TyUt98b7TnYMLbCM
z46M8Y64VxYppw7M2UPqzBdJPpP1+qXdUVgIFIPvK8+gnn2FW8eJJdtza9/H7Rzx
0atto3EgaTTDp4YnBGiSpzvnh6rCjqjlnL5eNDHGmT6NZY4EPCO1ph4k+9/4X3ub
XQ0TCTtem7J3+xImIKbLxBL2pfDjSGbtSIU7mpP+Yn+CUzV19Q8glPwNyMszvHLi
7M60Uc/8iqmxODuomiN1TfyAhGz0Gsf0W6w51guwMorFbb/YrEHBF/SfsHEPIBlY
ixGEZwro2TwXoapyiMSi0KiDpPt7Q/Rz3B/68gD/WqpqhanI+FXYfMIxqrbqfnLK
EnaA6Zt8AL72cKqxyNZyAmA+hymu1u6HCb9jG+2cXeHkaZ8ed0vDFWLfKyl6IRAk
l9EXfVGeTV78R+jK/VVtI2fDQndNcnWxEy9hgdnMJroog9LJkqnDH+K7KELMr5/l
7u4cc+SNVSqr8t6IPcVL9iKc7kqbeHbgCVQtS6eyv4W7F49x802MoVU1OOOLGY8R
80E7rn1nyIQQGk7OqN1YmcwycBLhYrQOtlg5ekX69EyO18gRNp4rOoMabN2/bU9r
gUWHB2Q9giRT3ZpqkiHtGTEfYbVvMeV3rwlah0dy1Tts8lMJ9ZdG7Q13v435AN8f
+qAnYr69SIhMgsmPRqFYulfmvAvAYb+DSSVrMbZp2i+mSXS9vz5OG+HbkzY6Icz2
/xCgOzu6a+mnHgFwUZfAZEVtbpWO5t8Ecxe3GuqX/45GzgEvkQRUZZIBRHYGxbsZ
+RyzsJ6SU9CDmPKhrHOEC8LnaYlXKMpnxZhMmIBQ2TxMMTug1CKJV3lFKqhSqVm3
Gx5HxnIydTT9n1W7Yjp2ZuZJpFEXn6fx1FRplD4pUZcX65uEHP6mEGCjz1uwjqQw
Z8F4lxCrWYZ2GagUwmiQIJwJ11ZlR9S2fGOazMl2y2ObV3nXlPERYnTT0LvtMEb0
hGCepk3dnKKqZONOJ5nxKVLxnDeRNcPRFVUySR8jPGPr/tv0EiNPvL0y1/VsgK6f
MtHDn23xr1s4JPNitKHwtw55WgAYxE7+o06UDk6u/Nl7c08sEqBuWT20rZF5ocjw
D9WWRQefgFBA2YWbKOrTF/KnOyOu4vyrC31/34CB8Qe5av3re/ZEQ+TBH1jFKP5l
qE6RcC8jAHcjPJRhHhNIYUNPxc6h2UsKexxsQm/xtVCdwe11yftRjRB8jBWfufa6
7qWwUwVweRYzxxl60znOHR9mHMSntUt3XMUQ6/FqxhPhgGLiWtJmeJ77w1B7SB3j
DRtiqvZg7cMVF7B6dRWsRdpS5pfYrapAyyZ8WI7F3oUd0kvscLsqZDX//ps9mNAl
Z/9dDA6cyNnrJON8tXluKw6fIQk9MwUnVt7o8BF/r4688mk9fUmL/DlEUdxK2gWz
ecqO/da8aIQi8lBTIc9Q+gbtY1FA9eBoFTtyU+mIDTmANL1Nqh+9c5dhXEHgpsSk
5P8lMjmRGQrnaY6itF/Rqws1oltR5jZBU18axgsSejRvAyh/DSldYtwnOKnoFzBE
R3wqQ09usnrx+QvBezQpFlFgJX5wQdl9uR4uyX8MjsnNXV+ovGHa3V+fbCdzPncS
ybbDoz2V9iL/A/vGLcXt6oD6rQmscYX9++L5vOB4w9j1a/YP0l7fgAyULHVYFhwf
DAKV0cZUKfPDy36fpyMDztj9bMgodu9LYB+z5shokrWHfxUzVbJHTejA+AJHwgRo
wS0gWCo4OidfnCXSSLD3b3spCqL1mG77vQHjbXq5HzDR2XeY4aewUANbl3PgRJ35
LuUdZSRw5XE0w3sUyVk0kB8EyFJ2tAfggt9hoxNMviKrU72bpIYz7txwJzFP4pVY
8exKYzMc2QHACX5T1lcT+DD+CyK5ASWQjc9ydmVr7RguSvb4yiK9pI30sZSgnVVR
vRQmVNETpD8nlramRTqD3SCE5wVKdMkAp5G12eRYKckB31huRjGgPa/6qtqOANty
9tth2RGzJEmXc1iuZz/mWf1fAH1sxO3U4/X1xHN8YLTwAtUDRLQ0OQFxAorIc01l
kK2yBFJimIpzsowCLEoqmvPjyToDPk1RZQagKTUHCFzEwb16MprxZONqazW30r7S
Pu4cJZ/b1SutkuyfUJxxZqFDssC2N8M1zLUEtkCNSSk5RK1CRcHiqLxVUK5SXJst
UajQWo78X3OyX0JVcdlE/BJJjTXIGuAzkJsNMEprgPnYnoR7FV3dvglHce+/3LZ0
JO2OtFrjuhT2EqfUwgx33E2ohqTLjvl9XBU1KcT/1ocETju5EDUdKUhe2NTILhFQ
OiRogJ6xb6BO08+7r6GPDewCA25ui8J9qJHX3YAWxcmE7HHoMj6ESiLm3j19axYm
aa3laT+dMoDnpHqtZjyKYrinDdO+SsQrCztsS3Mbex4V2TYlyjWQW/s4byQepyfr
OCDJFnhVmiigB4yGF/R0tDl5mmJeAfU+GcWyOgvzT7KMvoB2gaLikCUO1yoJFetd
Yetk08y8RE6gPo6AeNoyupHcG0NTJ4TAafO+GfvFSXAsCJ+Btq7L0bqbblGZEfic
qtKLBt0IHOKSfAcMoXwJd+lHsKvAKJ6zyZEi0C+tHP8pFtpbJuOswdIQwFWWraUf
VQgPetfNIjPk2LmE+odso77yPQQBmai4GnBCSVhvW6hM5EUgTvCKW59U0B51Qayf
XFFn6Ca2SpeC9v2PMNrNomZfbp1f/rlRGGsajQDAr3em72k5PgySh4FW4MBVWqPv
gQgW/RMtHVWBLj69JhYwycPQj7njOUKcDjx5FgalL5Jpfp58vsDsjRBg7rTmW3Pn
jJPDgHuIKsOo9Ik9vT/JfLUBRkZ84kiPAOK4T1B2GCFQOLK6bJdj0RcB/zc2gqDg
3YZaBQDzGyw4P4dVIvX/Bt9WNB5YZCCyf1Hf7ml/MrwKYf0T//M2RJVwOgyxSm7E
GLQlLUvZZKUX3mJmJHTASbDQYWHyyKU6vIsb+/fsqVucYcQdpgv4vX8HCygNspr3
ZPVyM8hBPwgEByIrBNB8HcvVCNmJMo6wwsTE+9ShHvPz6ShdtPR6tKWrZksH3PUU
uf+qVVWM3aqBxZK1+/NzuEEpA45xfR9H69FD/UcIzD89jUV00sQYqLlKPKweTZAe
Kg5IryWaNpLOcYDllj/Iwh/nwK6nb1B3anfXp7jT5RzKbEd9mQ+m2gxvCDTl/pm5
7okjovyOirC7alRHxffJq+LKmkwtU8/JQ60CA+vOY8STpcjzeeM/ZmXJKZJaeng9
xOEtbDUX5OdYl8oCBt05+GgKXOT1++ltAcqxQGPK+QHmIKSy7kuW1+EH7b2dOW0y
mA6kSeU7lnMqBLLXCsXGAuySQuFPEpjqaHjvaN0atyKqg4xojxDpCUKPbIKqLVq9
l4LUQdVsQi1MXbp62tGT/VZlN+Siz1ijYfIaQUTwj2aqXZb7cY69vdWpwlCDiy2y
oQv1+utJ8nfBeBTeVwdrlc9JgiD0/bM02ymhIktDyKY9RBKP8ikparHDoksQgNNM
SAhzRs3yo3gWj3KeqK+gf4p5oltQUbHdLM3D4AcastzcH9bFUN1EX2DwbDccbmTP
VnP0wQR/H4X4WFCWTEDewLzmJzx73ZU3cX2kl6SXryWBqPjiECd78oIB/tjuTC/G
u6f3Af1TMitgfkF3jFMOt2V8z9E5lgX4CJDcInBLP/GMnNNHfLjRXcd7NbepOQku
S07wAU/34s5fwek0IvgUPWylhHvKGBOy8jFJEFByywss5eMpYSltjuj2ipjJto4A
IOBZHIGictWTu04il4NcSPnrMg5hunV9sH0w00q/0W3TbjURUBrTi3DA5ObPQ8vP
bI8kN5xiHJkh5A1ElNdBi+Dsg2NqigxIg4qRGnT0vnyFbgP/Zftooao4iNacFjvJ
EFNvI2Y0CGBjnquUEJD6pmJoeslj6srfvkuGNtDWEnlfh5ODLs7oTmQY+sABxvBj
L+Kn0LHx/kLX5+fDnlXba0Z5NzcKV6SqKT242RVfEU5IHP2EQMbpu3iRnJLeoBOe
4y/YFDSLpVqnRhGhGfTHFpdfSrnFAMscggf2CLLddLOLlWK7TKBamqKPQg0p7lsj
7jRJAvZe8aVO7SuJTqw5Y/nR48WrsnZ86MB70CZzdKX6oDYHyIYDymEkvhaWr20w
L1fpT8IWMRrPNhLZh7MUms/EMrGUFwjrPRJL6zP29ewImH7M1xfexvRcn30HWdBg
FJ+zUaB5UJ4ekMlbfcwZgwbQn5QgNQ/7e27Hj9ocznuvSDnnUy4LMByI/SbCUqzQ
ec4dQGVhW5C7BiAY+eZ8FJZaLnfFX33R942rn5e0Y9mclxvn6JeLPXJOhD369Zly
ikjW2a3wXrKwXC2gOUmWuhzvEbM3C7QfTOogP9wug8+nxYR41sBOJWr+yh+2uY+m
clufFvZdIHYXansrVP4Lh/FXIxGRGNenlKp1+kPtgu4kF7jmR2rZAAXC7AOQb4aY
A5nROnfk37KjEJQjqKE6/rGh5zS7Amm0V/Q5d8xqJgUOtlM0frgYAxDs0O9/Q0vL
N3UBL8fHV9SyI1pt3CdG9BHYMzxOOczZcgC5ppIkhQt3d1tEkb/60lFZuXYarJMZ
OezEAPnItweqwlBH4PeTMXG3xIjNPP+HjwkJ92vCJZ2Isprj1+cUP+t+Sh8I2nHW
QNU07/45COVYUdS2v74U2Qde2GhE3l2EjJ5ZrFRprsttflUvwHRJS9VNyyws3hmC
7xoDnvKu0S+yEh+7rpCPvC4/mwViGr0FM1TUZSpf26dSxwrlm7eDXNbql7DNo8AB
74NVXi+XZzMTIEnJQ9UuC8xu5c6pzKbP0CdGRBx2N+19fXwG2UtcH/e94Yiuk/P3
IdOhAGMbJ/otthz6FyYPHARI96VXC+l6gkM4X2nUgSIWFA8x/FKGxWxTv1z8Opf4
ikMl95p4SrPx2nrPHVVT9VkyyI/qVnwv23e7r3DSkcehZxAOYZuhiJrW8G1mcBAl
VoI/wawF0DJBIRTqnrTUqZ0TB8g7ssAF7LtIM+08yNjdNV+LPicTjvuTTyscBayO
9dPVrEIqAmOl5FW2KqF8oo87wjWYCrD5NhDij2hdiUQbdyCJ/JHZ4ms9BU5LFMwe
OU9Dtc+FrNEexCXvCuMsuzsvpaUACBuxK1/FV4ntQMMCuD1DzpAMBhnKHbyzSDYm
o/RvKW15thPh4l6DXazAaeLJjVgssVHhAQP08D+1dneREmwz5Bj1GZcl+IvDfKLh
bB+IhyiUVVU5TvzzCJ+Yu3G2hp2Jlfnu3TD4t4ULX8glImP/qPVcj9G5dxtMgogM
tA5FOflzlONHLTeVK1eNqmVaglC3SsQoYwnA917CV1WqreFzK9A0DZJaI867y5u3
OvmLzh4q6MyFOjMXTanstKoMmDD/xUAny7HdwO341RMqEX7gxvRtDem4U4FDGsWc
PpZzsrkfR1zPQdhKY28wEZrwm+juStdJVaui2HHw+zwp0ZEn67jQTrsYCSDly7Ol
B08usQZZtBZfvaVG9uiJ6Nqkggcqku8E0kw/bGkIUIrERmPdkTuFaNU6FBFc6LXi
bGLetvOPjJsu1BcPQehL2WnoIKh7oIa77QewXc/JZXNjebGPuO5/D6pMqnFlFDGK
Qgwuhr4rZmnUWxqoKPZBjNhXoMXfPluxFxk+xxTHosasNW3sCX5cDvL/lnR5qa/Y
HqiBWe+nV3Pcwsa0ENoWxKfMefe33EITMRBYJ0YOLRIT8NyHR0EeBGw0AtCmqOtS
8Vl8J3u7/plH62Vvgs8avReF0DeE7kCinXL1TqWJcbzZ6D3jf96pjPLDdA9JWmDY
fbllvDnvCRwV+1JDmN88+u3rc8TfRPxQh1701CXXxrAmlvd7ozHUA681l2hnxu8d
ZZNFepMX9aCPYCmrYSGvBgVmZzVdUiaZ1FjD7H/9XyZqoZZXIiVqfw/35yoMHJEK
erhl0j4PnIt7uHamc5Zz3IwkW8wqvxyVnwJXMugxsKw1Jq/QfK4Zwm6iPwTdcqup
BVSvqGUITFTwFmW2J0Hr0k9e2nEt/H7zgNlZlnN1WMxIalNE10a3KaVNnvev738s
AE2bQR71y57URsrrN/VRDN1vFxeDtIrJGUutlPvRv5j7TGzKjUuV762bLKKx1i1O
psFFoToQJduafb93Osom1TYXAzKgwqEbpphHdquAgGg+UMxCBtxCg6WJespAMFt5
eD+d2cdrT5VESwRxysUmasOmJQRDyXSSb7AfU8okBb6DXBQOohzwSQROq9fWlJZC
lU98rQsu3281g6NysG0Gxs0i+PfKRswzeCrRGoZSdFWyRbmd+60eEtIOyMQ4UDYF
cyVpMg4iueJ95Txz1LbWPP2yniTlPMkDRn8COXJXvm5tbidiyT0HrsaNcqa5Fw7f
/l5FqhzzQnapeRQx/OOdhkCqgxrRxtEsUoImMFoei7Sok86WLANPJKtGaybwZqPZ
XdRoT5V78Yh3myTJ807IDXQnEopSWMXdjvLL/E9m07n9gGT5yzrAeD+YQ/NeW0R3
iRchxJRW2fgaHPbQDn3rQXOWsvJ8u/j1SR4HRVunsTxkmfu1xDoRvVlygFI1LkqG
RKP4OJuTur0q++bg9SwUBHzqaDKvoI09ZeEhZiEbzKJygse5AtQ/q7TSA/Gpxiyg
LeOYXARlrxkkPYiHsb9VzZSDwAvqlAhpvO4Rnu32HqVcYP+PkANk2rcMVr7PZXZQ
W2myOOv9Ggt2Btv1sLFTct55FkWQNZr8jGhmRrN051XjUHVBEHoEIJJFqGIY4xH3
yIT1gtHC8tA0GwtctRGlaAD9RfqXyxE0pT8NAP4p2u/uxl84UdYeDUavNok7AGAh
KWGjKS0srGolKY/rCATLJG6kxxQq+RLyMxjCLVMnhWkO6bQbWT1EXLwmQqytngV0
szRz13O5muxoxEfB97o1y+TeLBu7VEZAW1k0G4w6+ffTiAvYg1H5JKizRInH/pE9
C1Ip7nMVpCDGscsC1DULCk0ubrRTXmpGIogMvdabzBK/H0CYqvDafQW3ka2BSwwI
Z2wqHT/KxNsTG4HoZSKewHhKTHSYKyDigkpgtmAQ1T9qcZZkTYjquS2ACDDwSyAJ
dotSbPV6lgFZFvjtaOR4HJ1Mw3ESFeNuXgTmfRJ1WN7tQau08wi9Jr5c5H0hBW/+
yJSCGkdjHKDvTVCY11pycCnbay3JgEyl64Ch3ITo16A866v4rd506+bINevmbvPm
7Qi+cqf/SEer2vQXL4pCAiKcucbXakvz9Q8hldnfCQONtsm28zX+kFEfFg89sO/b
EXYcP+ENEOfq+0PFrzU5Wkvj460HOocC4pfRTsc09BVCf5by+HBMMMAdoLRa3phn
VhnmPFxbQoVYokQj4WUAgr+uO7z9WwrQxnxp3rwBj4Umu7Mg9cxhO7rHjSK5h2cp
tZxb0JhAyHKrLI4SrmSAfzyhscQTbiy9LhMbwkwJsXGkrVkVc0iKJbYP/dHTbWub
gKsAoAperLnDQAKDz++EL7kj0KJekKzmg6f86DXhU1WtaP3UCNkxfjfTFAnXijQT
ZiXThW4ULuCJIqMR5WjxtFBy5gKXdLWm72Sg/BjGLPlLrrll9wqqP2eGZoWcu8/G
Zug4aZ65DgVauv3EAsUgEjRcO9Fx7o+Cf1TxGSL3+8DvH22AMHefzVraXFUzhhwo
sfwYH3GTmUeQK7ED3TNpLSX8WzpE9Obe610G5tMXUhlZbymivvav/NXeQVydB6pO
1aHaj4Qr8rzh5W3lwhfp32GSipScPDnWSQJNwdS+wnCctK9nNofuG/Rtsb2g0ujM
fZEvT6v5e5LdwPbCF0FfE970OcDxqxJXG0dqi4/2giMOmErkrdu19XrqHhsNEmvP
V8x80mXhuwFgh0YXPdyvkxyuLZ1Aa9oF4q63Sm04BaPJ/xBXkACMtUa24W4ikx4j
Fn1+/TL56fZtcXG2C9BRiC7aHfn2LCNPBp+9sXlJH4pJvhseIKR2P2PMqmeSYNjK
Kboel173Z8jvbMsxZiH/sMcT3klrB5+TjjpcCX3Mz8G/UBFxsbVbFZJ+jE/fzA6W
m6xeNxImUC4MxdVCGzl8X6PZWKbupuH7c/CfQf3SbTxsXvU+/Dl8oKt/DB98lsjr
UBRt9TsF0Kzf7ddC2H6CaRuClGLpxnACi7iwpAtvUtKUKkjtsrHNueXAdSuMIJzD
o/ggCwPkhAvRRndeg9g/LMc6Zo7YoQj8EhWu1+ZSDS5q9FsvkeMkpqF+OQkT6n4X
mHi9gswrpAao5IoKmWHXTCgKV7T9tzaLtX4bsA2qfe8KzFMSmhh7iqDSxNQsGRSO
XBqVhdVIZ/ZqMJI57aIlfEKBqN/pr2yTPoWxCJTvVZLtQFXQuMDT4fugo9yBh4yc
pgxe5VVJCWfsRFf41uVeXcI1AiPUYDswVr/CNbfy1qy2dVo3HAnjj2XIBvIc+y7g
FQE72SfCVm+oHxzYGjzkE/PwapjxBJ1dp83SgWpkEYlyTWtYd57y1TZXyEevGrNo
RnyawiPufksrEEj03dryH76zpsPgMJ++FU5Xs0I4l7qiKDODHw+VG5qNVfztym6Z
mSsAq7dVukaK638rm34GNJt8S8OufAv4B2voCnI67vG5cpZz0MQlSA2jV3QqBk8I
2PxT1Awn9iKnhylDB3MJ5NBxFLUV/6eNTBo7yfL8p449BvdpNaPIagBNp+dgEuBL
aXvz9+u8XdT2I8TKv6FWEAqk83VZFe5qQpzJLyV8xz5pa6BvGi0XwRJkEA111fKI
Kw9+Xa9yJ0fspZosflS6XUXlSdZH9GpaKzzbo3t7xWkD3K2XMfbPPUOCbfrOJXEu
vtqlIbPUhIoG8D+0/YbQHUnjx3eEdpSkZ2E7h9nDvFIDraEUfLkPeTuQTx/35gTI
bCjc0+vdCT9C0PyCRgX4jl2qhRiZMR7JCupRTSd23YQjVUb5RTmwmj+OVDDdV41J
BYoRFeMQVtoiStAoQfvUpE6YXuVnqNJi83OwV8jGlRVhzsmK8hUGT4En4IFBdm3z
ADQ110rxKGjWYEdNGXH77bk0BTGKqb2QMjsAaUNroftK8a+HFPV2pDIEs5cAbtoA
kDq8pmhq64XO0ySeWq7Repp31OEUOLlzA2kmz0wqciRRaNp0sJKy3JBbW/KealsF
bbeJNtaVnZvT/cVHGlBwljUYZ2juHDU3L55HPFj6RwNTjziX/qbEV27AgMo46eGB
LQrsNZNGTc591hOku8uFN6avH1GaJhJRa5RkbArY7h14KNDptqvOBR0PmO1xbxF4
kqBNg7n8V/FQ8bei/aElp5owHvmaXYMToi50k3tMas70PLCiLgojYg0dM5cfmu/x
pt9ybf3YJoWQKuCrRSwoQPjqEY/8PjocjsYfU3BzabxayWjAgJ/Vf20OCR/5o2bs
8D4n3ky9R9KrEEU8UvD5GShG/xLfFe2iVWhIjIJfAFvs9awhjW7pIpUUZn1ns9Wm
k8jDUqhksdBTzGtO5kyH1gJn8E5mZuJvxTqpx/bBK47q5Z/07mFbaPblKy9FRXrW
c6lsL+N8Bc6VVG0kuMZmSzM8zHKtD6Zv4s30OGF+MfaMzZ3bniV0IW/Wh4JGDQ3f
cxq63JkKSiJAg2QE2rSrNonnLsVSXZxKD3bn/pSHU7Xw2BpuPvy/i4PUMEDBmQ5F
X3Z1m6HMnH3JutYMePm5dkDPF1ah4f3/koxbuUOy2qwK3iPSmRAg5n6kdgQ2f5lE
VacNVaWWWT4SPXU7atBkfwz9CBqnD/mYM92OQLcNr/s7VoB1lTt4bNORjB6Lfe0R
5P4d4OBdKrLebGB1EeiJjgdDVO6339v3SQyHeQ815ChlHfgu3jQa7DtiI2AhguNP
HgzimmlUvd/NOZ2oe7R4pC5ix8IjXAtndhrtJoCuB2OGfC3LZh3jz4y8zsla9brK
9kPG+YLQtufeYxfcoMiUvH2qEV9qyOv8xeWTcPsN7idA1s0anBGZ2lUuqiqqvAEA
bw5GK5xzMqZ8ShVKfoXJxoye83xZgW1UsIiKTJgvuCQTj2FlPlXgdsYRYVP6y536
OGUdnzpPhgRrC3nCirqVDuJcPu7BZesEV2oGABx0NBHk8gp0B3Za/N9lkdiOphe7
u95nDSjx6F5S+2wEGJAVG51Pfcd/r63K9DGq7vbGaGeAfcR6tVGtryw6gKBUJGNF
/8PGufhIJc9O3l93aeFIDLsUPnr6sePxQC9iOWciEKc+9jSHt+MoLdnoLb8nW6MK
/zIHgFh9t6AWOtK7enXb6ZmNTJVIB9SHlhVK5wa4lO4tDtg2Tl4zcnKTMGBzglax
a85+F1pAmL6gZIo/U95v8ytbcD/eyiUmZpMaDVxJa/CbPuTFySnGmLpjERfYdxqV
IGJ0iMwVLUljekXTcY1YU07L5GsibsdDrGftX9Eg5L1xd4msDNe4DOX6X+bJWBZB
BcMTwZkec1hUtd/InSjCaNpnC3ZrXrLQ6yNDofLa4KcWvGE3Fhpflhm+easR7DrF
P1G534ic/CUDzHfx13RWarOdALviq3dxGfkt2HxZXBEEnW0Tv8/Zx0dYoR1kYC3T
1q2gkrB4pnOheDtSYNUzgxRcYmfowhix9ESi4TF5VLhiTvPGoi2KTzZa9k85EGjQ
uNwIuTFUOJ/eFEF40G7uT/PwyBoe5HvQ+/lI8GWJM1UZkUd19kdK8NYq1ng84xt4
MuLQJBBye3WhEb00Wz+MCyNwLyNZblhTaMOuNEeuRybXGFJt8aRayWw7jUGZ5N/s
jBo2plVkg8vb8/myFt9aeZ10pwacish2R+IbxQUcYpaisc5WiG9Xh0saBs9Unz86
75fD6+/4Gg8bJpEh3jh23EY5DxQ2FgpnnVY0sxX7yjzsflT2oXzWXtchRCmzo5pa
Sgx/0Et0FOxivwuA4E42jxTMfcXYhbCjOOzP5lDk6PhF8CwYUTjsStaB2HYklajh
XWX3RuiyeN8ytbPA4pR/74Ixlj2RZI7XamIR7FtHlq9JkLwwHdHX6LqoCmHS0o0g
XKcx0+td+7tYKwf1R99iKyW/PBsrlEdD27X3/THO3ZpR5qI9I1FEhA3K4yTXilS6
yqrYq1hIdDG3TWuc0UUf3tW0ll8xv2Bc6TqyCv3m295D9nbgOVQ/fuX1fTZnx665
pKOJTQ+cb+SscH7AEZzmAD4JLW846sb6IL87EehRMsLUg028bmXhTD5rw1KOaMaq
deqNLGU7SfLnP6nbO9OJx+1Tjr+FQRV3AAXEZLqr0slrX3BFUJcqnRgYFlptVzVV
hdvZZLqbaMmH4nkshiJwBVtb2L1iARO3nOoqfLMRczMPKpY1vjH1xBbTrhNBjhtg
wIEwfaomuhYXYq90R17znvgW7DT/lJkOp3tdO84pkJFFw8NTmAg2vye+pQ65Tqf8
mOzY+kjebDyrzY2C4YNN2No8cr1OqIKGko91wKHjHrR0Nbz5uU7LuODtr0hVCmcF
QYB4HwtKf0UAGdcje7IyDB14bcSOJGkYJgj7zl1iJBzDQccZul9RB+NS/BXtmg/P
RKy11WwCpBaK0zPwv426LoaNpzkWGhAWlaFUBpFoQdap+eY88x6t3k6LPmTQeK8n
AOy9TxCcDjqSl62lOZx3GUR4ZGn+SWSoXh8x0JvlUMmmXOCcD6mGwOPUFbwQeaqX
ywZ+fzgXTnDp0nTjRKSvdFPks4HJ96CC5Ld7XFaXGFrtih1492x4e8CZiVzJRXWj
cVr6NlYJfpkT5Y5hheb92OpJnpihGzWscNIT3x0Vh3i3Xfa8VPt1pQj4gVKGr7Ik
DvB+3IaOdM59CLuUK76Bqi6bBDTjybtg6bpl0ViR1nraxdCNftk8YkOITaKrZbrp
HZl7JHcNgg8RU2lkzpZm3BePTC35mIrMeQOX4qIGrzUKeO5lHsp4yPLxK9mlPI3o
M0YdgpvtbwSA7pl4j8d6/8O2XYxcw2FoZMoN4M8KJCZhHtlX+1Xh8PdmTV8EQEE7
b5Ek1Vc0tjsumhtTqwNw1yB1BTS82ZUi8ukdK//QvuIcrKnGXY0tcSzdeA/jV1b/
J5Q1L9kYS049bmqzEV3nCG7eFGN8e09WBD7Eg49x2xHyyHG8ndxGj9nx7bHKLy32
X8GDFHBDb8QPZrw0bOrQQNj9nSV0aa4wuSFui/kbQIEEkH+cnXCn+AInlZi+XYQG
rh5VVMhmuy2oemdWej2KoslBdAh+DRRT5puZuayNrNuf98gWxrLuX6gyHRRx8twd
pJyFoRl2IfdxKOXHyN1dLxfy/fM65br/Cf7RuoZgVKx6FYJOHblvqYeTh9UucN6b
7TPd12KStpvWdPuu8Pd+3+9WkSGUC1eqzpG67zKnFCdoc2275gMNmZk4q4c700Jn
z3GtsGytAcVz/jZR1TgIxacozp4FQ2csv7yYaiAO9phsBZT6xHlfW4cUi4t3pTJV
YQadPHze4FY+vOs2RRkMPpZ3Tuc7kQ6szwhSd6i7ldq0Bz1eVawWAF+mneWGxqBJ
D4XVNOVsfwdOYfwttyHVb0WQDZyWnJz6jGjuhXAZv2EhplKHebqpejjkhN+sgBri
16A8K3I4c0CKOuhTpqNOah+tkcXo6SLqkekAGz5/QyhOoux4C6zAJIY3SQnEJsKX
Lg92rE6Lf51ZBRbrJMZdIHv3cMRfP7CwF+GAlYR9WKwVQgskGvY+Sx4PbwGsb+jS
BMiVFeGL90X9bwz2Di0/yOKD7NKy5/jHs/TUdMGhZ7FAZumNQVbwozWams37AkON
2v4zbXBpogydUyZr/NfyMpfYlifPv//K74LW42maoh5Ld9M2go4j3iUNJWoQ5bSE
vFaADOO4qiuKpLPtGBzIpeEu0+HIBrJKx6087wG2tCDqMVQYWP/mlH7/TMfE98HK
JUrF1mtpRxy2r1BfhbaZB4XuY/P6+x4+v55YIc0ZK8/wc0Ne1U74fMhKGvpyWAj/
CFfc6ppBLytUCCxFpJjtpCyG0tyYAsHcdK/xDlEfUKDQBJyIOy6TTSXws/DANi2h
eruD0wic3t9TaiiL3rzd906pyfA6e3eRWCr8ZkkzK3vn0wf0YTFESOyymKmsDfUO
InKh+r3inLnjri4K9olA+eMqkGkstXmP9z5d/iO5MnwbUEKW4mDKfRgGd48lbD8p
HoivnTAQ3uyJcUn/UnVmME62ZilZDNe9//2dML2IgWCXhkuHOWOGt3b4qZplmufp
0kDT2SFgCi/atp+VNnDKxzY5JtYAQujge2sF0Pud7FXH8JohZ3uUrtl70lBJqsdP
ndLcRoJxbjJI/C2Vrxfl+/5rhM5GI9OB7XqfrFZjVvKDKUDxeb6rWtSKIOw5++tu
6cP+K/EpIgqwbaiLMxKDyFyZKpl+Y7oWNP302eeMiyeU61Zhce/5Jit4FyDTIvOl
69kdXg+sVidD5qmjNsA3vwlPLDhVnC1uqpsBbBeK2ZP9p2QmqLUMEDr5bPE5+6tI
6s/7Z4tkMIuTfmE+OyldTCD5guCsRmO3+A5aOGNNG18//lDBgrZA5eLmUDpD78ua
Xi5i4xV+YoP0m6MKK2wYKvI3GKyrwC5TimkW7MQvAYyluigHuhdeF1k8g52NUqSp
kHUKOABbKfcYWUBxzwhy+72r7eaefvYf2JF5LOgF9NZ321+J2R4RuZf+UbnZkS6O
2Et4WjptCJ0Nk+rPzi8lTFxlkLmT1JhVkTak0wzJbuSh5cB46QgpLPwRUKV1AKM1
05ss8J1k4mKPETieZr2R3inGihXwcAKKEB+FW1ZFnCflIJ8O4qeSoy46aAWgodW3
YLaHsv18LCZplXPvbts2k/Dau6DWWIiaqDRXbzppM6Ls1DK1Vx0shbTqM3O41ILU
qgK73+EZetelqSXEfZHYOqejJHJdvsA/qZP8Nfn7cJMKFu/LchVJJcr1y3A2jfc1
Id6ELT5oH+rrDZpXG9OTFYNvapL3vcRDOPXmp3x3VQGjXprF6OJg8a71jf32alzm
d+8M+pvhHD8k98zXb9py0Soh3jVpdys5epG+onBEZm6xDN8v2BHBOWo2MEnPMm68
bPCKthBaDuKWcUpFJzwzfe/QrQy/9/q6OfsrAGprhSPFL8+E+tHxdDDuIYSuOaMg
EQebYlRUxqVJUPNTWu6LbheXj6oZVsKBAnpe894f1pMs7BHOI/xwAkQgGKP95CEc
C2sQkt/E8ZbWeUZGJ2HAdyDvicmg8u3UrDA0h6TaK+gREnywWVOTluoNTDoeoy4W
ahFSoUkOkAMULxqvJjNuBZyr1QKXw6cGhhR0vKA5/N9ya+hiWmIu29J/A944dGjN
Pl6eBXbZfSk8FvZ22i7Eegwi2NM529xOcCIEJhKWwBCtr2tWUZG4iLqnjvBH9NI1
tcaOfXEevXr0Lp2Wp1isApTICH9k99Oi+BnZOI4F6z+ogbk0O+3SYVaohRygT90I
m6S1PF+WJ1r3CT2Jop6nRz9idwMdqzpzrAZV88kTxWNW0l+DKWHxroZiW9Aq+oIk
szdPCOKKvUMuQ6dMDMqga97Sj6ZYLcAYoSo1LCOeXjMcIxIjmyAOVapAVUATthrO
I1leDH6uIO/rXWEMIZF4Zq8uguZK4mYSSvrC3kNm5opEAkTQ6T7yG4acK34a+i6Y
ctNF8ErG1zEYP7j2Tx8lBXKqpGa+fb/GtT2QTDqrPzWr6M0gVhcXF6kGRf3XjhY+
zjYoabU9+5TfSX8iPVRIB58XDD4aBcWz67FGUUqtwm8da2UtaETTKssa0rVgGsMI
B4CRIyXL2Cr7F68SjiZ2VM4ZpU+6v5Pv2pxBvjXSfK0RU5MITxC1F0FaHHEezD6b
DhFO87C/ojG5J5tFnQ99eni9sBGCQ8DDhnw1NgxoX4fYGVQXJOvO823Ro0MBitD5
wxJDT5WYmtTAH6rplsOR+g1/LpLpgqplGQJPWbvbxQfRXrozhChGOFfXqzJ9oTuP
jKvH+S8hE8ohQb4/E14G4DMBTetUJGPA+NPRJMavt9CzA10/dt7vYKYCson5zZLz
8YT5VgAO6PqjYNFCAfqdN6dKZVgMK74UI6SKuBQCDYY0VKWPVk6+PrL+bv4xqs4j
qBGvQAWY4gFB4u6cykQVMtHjENTKrcL5fAwT32z5Webr4qJMvH6PMJV7PIQRZrzM
YFwdNN+93tg1YJAUoQoAGjaKjc2UlTFe5AMYprBpLL1JKB0Qw734fQgjW61zn0a5
ojgW5moBf7y8KASrntY5+2c5VUhHjUXTXx48coK9/ucnQwcr6dafQ0SJwRcBUk72
TwbgztjHkFO/jt7fJYTk9/K70T2sZyMArbsSPaSHW0jvNK0Inp2wu30e6LDcB8To
m9vg+xqeQUwzbyjqlusbs9rxCm019ZkQJh4MjH/HaJywYdhlMO0B0Xd6+G6TO7U8
HpCYSpAI3ghA+680zpRrE3Gug8TlUsDk6mEC9aefkOtJ2rjZSDIC9m2sDX7m7pEI
9/RDVWjTW4vjmE+vaSqLHec5Cxn8J2ydJ6dicUGdtadHSZwKUZhTW10m8YOmnSXq
YUBeVP3tOJNX2ySrvHnI9IJIAVuJsAHLxl84H+57gYWa1hWbQ9xm/cvR0h3jpdbz
avPzJFrtVShUCUGGvKsdJm1Qp/ffjYsV+Qmt6Dwqu5O1fbQtsll1ZYH5anr56Hkt
NMtQIDWZkC3iw/BMt0grKyEnK+yThcDpZ9aWxkqu5I+kxEBVWWXD5HPtykspATrS
HmNyGppdNViWyIHy0ds7G82So/caOMjMsUzA0GypMwpWao7OxlsmbJNPczEJUpc5
3e6yhc3fOD4+3qBqPcId+6AK5HPgzWlOlZPB63jxlLi9n51JEl/ipGMtYDTMAtHQ
ZKUmZ9/SRNYk30x696myJEBt4clIJezTsPOidWrwHGTiEwp5SOXXwTXy1M+zOlK2
VpclekQ0h6+61MwcJ74xxTQthfCZVqHl9byhReNGI2RI6MjvbOLLEApHRLfWv6+W
R2KyMFBYWuCAnxtjmwUMw34a09kBCHki5WSUUeA7u6JLiTuLC1oFpZ5WPOvnmS8J
4sUFoRgtPsjv7vtpylPLBTl5GZZd4QE9uY15Pw2bD+yTI8/y/pLBSOkdMMjepml8
+m1k2jtVEszhL5/+gf5aENku/9aPL06RCDWatEJ/CVHTKd5Ii64reRUZMdti8fGM
RPlInl4maBjbrAJQpIUNr7gp5iC1hb4o6TBnLI2UNXS6oDHLDOXn4/Wv4kaHbZBy
xku6lXzUTzSj89Mb+3h/Xq36ldPFa6HK3UNk52pmRZ7pDFA7kDHl7mcEbCt2HSIa
UypXb2wu1ezFWO+KJrOiY/YXgEU+aN0A62gNaOEfhjdWYWfXihLF10pBNNIEx3oX
UXll4obc7649p4UDhOAGSjPFiTpNgPdRy2n4xASoqZ6m4CuBC8Swkn5Q/YIgUe86
nFRm9yt/xWI9ZuSCLYAjXIUxf0XevN5RyFQDtYsV2dZrRytDk+Vh0Hn6fLMAaabs
5SSYYBavYcjdbHRr9/HkPX6peYtVo/k9yDCA37uormuyXWcThv/Ew0tCYxhglalV
K2iLUe+AzQsiBOVWu4iFwhiGsk5VmVVRdX/gfgH9X624H7HOBmrKnvKuWbYfmwrt
rVSJDWjJseV9A9bDARFZb3erhjIkAYF7WH37aSDNaOv/8t0lxZyKPF2Rqyy9X+zA
2lCDuH7Ab3/mXYT7m8KK58wSAx0rzdND5dCYhAkfgYfxlSFJkk43jeCLLMEb7/1v
WX1j30ylMp0HC0DiQCE7Gokpw7QZS0QWbB2j1yZds2YykRddW18vYwbdOhRN2kt1
fGGr2R5J0IsX/m2snMxiR97CKUqSvBOSp/+1Bq/mbmiY0p4Dlyn5rQbUcE6agjdG
ZhFPOwQTxUr6UQLe7NFC3mFWL7/Dwk1azZ0/WZcVvrAiWy204sgl9QyJzvxATFTy
BYYYoPYwaDEp/x1JTFdBjzmt9HFRFmasEOIM3VeveZf20eDZSRhgjPHp3tigpjV+
hdhtamUJf44ZzVpN6z1mJGvbi96ECisJCEPJblV4AAknCqDNrql/oVu4pHr71yxQ
0zIY+rOPwdbnjmtXh9FEPjPVxDkewQxXrrErSnAoIH9UJasDb6osc0kdXgYDw5c/
xKF4rM4rdiDISIze1YyggsqvnMkR7Ztb+/rOSBuAviiBJzlA5CYFdQHbbsjOdIrC
TvRgBzMQOMYj0LVaLthJiuwkiVxoHDr9KSrFcFS1Yioe9xWJChQ6Kx3+GAegaG+V
VDyQqBKTk71mNLB/WzzCiam9priYhBJpqDTW5zxMSs2db/2T3vxxfmmrkJ8dZ0fK
xNeurptvFVsl0YQLX97pOZ5XQPd6F3/Zkyur5wPuRish2YuBsIg+TxC0i9egjCxa
K67g/zG+4DxjsfV1WIb/3EMaxW20Ghw/+ZMxAQWu0uEPFtOxF4kg3ONQSCkdqhuc
/iCZxsMkliFmQ/SGMC1TkTMZdVDMA2wmhnre09qLsleKLkuJzQrY6fPOYm0CJkYM
Tm/BriNjKySsbXijXeYaHtQrrWXB2fJIX6g2Q5AMeEjZics7gWQ0U85Y9i3Sad8G
HKAciKkQ3kamAJ+DK+1vT3JVnsM5FggpMvywU0Tv/HOVDzYLur1MT8DrM32gUTgc
0oxDezfMPCE1DBKHjCRtLVY4e4PaVKXGxRMRsVUvrk1k9OTTYoYtFAOEugNcQwGp
Mq6gfy3Xn2lO8+W/Ary3epp1koU4mUxm0bNh8tP0bhlt2bdVxTuIFcPZ0PQuS5DY
qD7DJWEKqnPMsklmzBaGoUZrc54zNOvDWR8BkGYYCo3LnjNQH0RJJyFsMmbvmcEc
BF+WS0HCPm9gQZTnnSxudwyPONSTDcNYWdsipHZRdRxRD8fJk9VtTZbouLo0+aPM
mabG6DdslATq2cViHAqDKydsrgW2gRV8dbpxkWz7wfTWo5oN50MyN8Vj89cIDBGC
RMvrOhR7kTly8EyP1sgmwZe50fhu/9aCBbP3brx2je4IaO/hppa4QajILU3quArf
qmqKbruiqbN1BUGoGcRKSYcyt4KOdbSS3Chs3t9G08xMvmQ67tjpWda2cEsManCO
0x5wgwNLfMIGLajYWr6m0+Whpadx3WDgCK+mGxy2kgnDNCoePASIYI22ImaWJGD7
R0OlsMCH2JPdVRT+Ji9qlu7I/3CJh6AHlqMcPqVCFIhXMEflNrV0R2IR9TP59zu0
NrceZxqV8qqcWnE3t+80RGMes+OinFyXll4leBJip0hSgOn7W7r7v0FPdUP6bUR5
Pc9fZKIBKd+/fDUx5yCBXbooZhTNBEFJD2YaGgms6Cjfzv+kaZ5w40oN8Cp+s5ZU
dblHT4dfBiSpHz6a9VqCptANACble8WLWS+F6lMxgjD5KZWZIqzzIYXOtmFauxop
IDiD9K0b22F0tJT7Xtz4jXbtGXumw4hceVGqrnDwPrkd1y6eTpQql8uYf+jSuka9
2bELXOLeDvi6vvG4BKd4PtI0FYpdFCwbL3cgALiFhZRnsVTv3pWrlTI/4hZqOpSY
/tt5ObCD4dCqVftfhgx73gtvW/B9yxLCu9+px/LyuhYWa9NtwtfJCDWfek6qLZLz
uQjuwvzsJ3RYe46RhY7wxwRjaDUieW0TnONgnMMobWX3KkJR0YgclefhupVGuVYN
dtvCRmo2l0+KfElLI05sAiMqu48a2UZrejJM39IjEHt0pfvaejZ7z+6lc9ySQ4Yw
iQ7bvkG0rd83R180mPbBvJsE2pBI4/IAGlf/sI52Ev1srzfQzp/ke/7WNtsqD+v8
ZhHMWsFT7t14Fkxx50Kudsgz0uxB3js3nptk1xrJimoQEnQkJyYTMk1edH5Lzyl5
LbS+6K9P/LwTC+deDP2BIEAAIi16+ZsCiWrCsVZBJQKL3l4QTyNSwhcIdLzS7TSe
nx+bbrzfR5DbYCClenDa1WjzhtZmWupdHpIFSWrHTpJCxQOdfCiK6KKXVYD4zrWD
/RWoATcmXubPaQX8R9WXA75XN1uy4MIyMKG5x9KBjwfwtsAWq9Fcm1lssvapbDNn
GZd6Bhq173QH7NtSrZtLF3U2Cg+ZvMUsipOqeYVbgwN4Z4PyGPjiOCCcaPHEdT5H
dUJiVMkcS6O30MXoMKGoxBC1AKgdwK7yIz+ygd4esC3hsQq+tadPO9c3ng9buItv
l07UE8RjThgvx3bJecDFYVY3oOcW7GAac6Cp8U+sgeDmzykgscv3TgNTqmCUN2Qm
AHR4r2vfw/BxBfiuHjE5DvOGzjiD+Fjl9hrqvO8hHMzEbZA8Pcf90o+Yu3S6ad1n
vQFfzqRKnVyyeue/y6NQgIaVZWlyrmoytXXSFtD3eD1ymv9UacW+7LQafeaXH08O
1jkTYM8zH0eyjtkN0Wm42SkTmSkFA0C5J19PUGc+tff8CsdNxtZ8IOV7T2+ZRs28
202ffxsIXmWx6Npi/m2okbkBCAgWS7pRbQOTdqcH6muDW4gmsfe5Se1W03HfQOIK
qBK69+AAGEaXcRuJF0du2rmTgZc/BU/x2hulJWdptgGO0YcwM54pvNNQGpbXRNC2
jkC3EFlGnowf0qjopRSDE9Ul74AH/wFz0zNvSLfmKl6E349fgMuWk04V73+Nc6CQ
WWUGzw2N3E8rPj7dKg3XWxGsG97quJxfDFpuovfgOfH967qlIMTVhTwyKLqLbG6A
6UIAsVcKtpkHpHUoOUdOC/OiDG+okK6Z92BDxl58tmJ8HTHTzr+KrZEqipT7iAZK
6B5WZvK50C7S83A8GmRtsItkf03/1GvckDNooVnJHJAPFpLd7V0hVRYyCnLGRoRv
kF4GlBSp38zizwibPnM6Fwk7nRdyLrR/LNED6ZzR47u7YCgLD+ZVEuXiuuxequSz
ODymbrDa4qdd050pp3lNO60sUeg4T63yTcmd7pPfpGR1kxk8Ifl3StEqTmQkF/o9
hx2VloK/CCzACVMKxf1OpJhJZqGb1g2fgnEJstTYDTcnumGYuFPAxQ+YTZ3P/y+S
jXxAQKf+6ey2owzuDx7MSaJ2Eidu8FLZL6g5t9e/gUfTcUtVEwK14UsWIJShbodE
fniuWRTVTbVkFpFRqRWXRiPBMRBOyxq0gVxEo/9PiTRjhEQXwzVsf7AjSkBazpPl
2R+TSsxG7uXVftGI3h/gV2L+rEtGoBxI1+YZJtBfTEAlVS5FSWOHBynQIZMKXKHz
k/x9G8sXwaL5ReAsp5Db6JjHbizVXhK6B0w70OHkvoOebNWlNMyYg9iR+RahWJG/
ojdr9U+LCWO1Nq3DPqGy8KUost6epersvR69FZoQyNqa15Hz5orH39GXUSJ0Mj9R
L+y91OKkaDVZeUFE+n2xPCS9WG2rFmOGLy+u3EJSt+krhCiXYxI5XetXXl5N50LH
FsfbN9U7LH7hwBcONKm4ocYIO5rumVmvlh/ndGpfd/V3AhvXFkZ8YJftBT+xqFfG
hDJqXhJ9LnIOw8v0ndnq3Y5DuT9FbeBKnMdoIFbHYLOi1eGvvn7TQ6O3cM/d1HMH
DE0HVd41VkYZix458vz5LSl2TnyjZYGTlyRKUY5SWAy1fauEHaT8WxV4JkjanwEr
HYV55B6mfJLeDak/MXcB5Ts4v3d6/ifPWjXCaHs/dfPpAybiqxpOKQ3lQW7AZduB
lr2e0RwUTO4sFS7zfQHVqJfPfySPnjNVb4NcLtg7L8CECWN+NTnocpIhWxI1H3Pd
4o+aMDIboS59L0kZpUVTJMfCg/WUy6fIPtMQ7MLbEFKwTKydyAdOs9q5pQIjcSE7
t6Rjx3V6vtR0WZbtv0fYOtCHPFp5REKc8odBCVxJ2rGPuTC0fGlDAe4Ggv+B4m+S
Ge+Q5DEDrpPAviC8fDqkvyQv0wxxqUlYige0lW4UmRq5R6Sy2NovlhakFJXhYFBC
tMWg9jh0fQG84lXGC0aKKjrOGa720zdTA1ke4KDekwv9MBr88cykLq2YG4pY5dJa
JgQGtow+DjVkbV2cZep0EEz4+FzevMRh9+tL7UjTQ4p8zZ82k/dvz5RbA/qXxjQ5
XlwJ95hkOd1kBIa2vJNsBOXsgOR+S27ycBbD8sTq3ukrEqtgJwFyPiLYj7KQP7R4
n4iJ28qweV64zj/MqrR1ixskUBoQmVybO/OshAw137sRZg0c+KXnIsf6TTc9CsqO
Ofd3YymFv9fyl4L2KpqPprn+hK6SZkD3aiGlW+YsprRTRLAAnu0PbbdkqSpGL3sF
m3SfLqxzqHBgaoR4Mn9CwctvV32E/4PLzDCeBcWbd+mPSyTTsooQkhblf80OQHLH
WO+feoNIILsEkeMrHMYr4ZVq5wzPixTMukTb0+UE+SzyMFEJAnw2ixwi0+eiESWh
tRNdRAxGzufhYi08XupvUka4SbpsLn+xs9lplgs0K0QgDJkA/SEZU6fkxXjpwKTQ
2XjKCP5E5AuS4MT28/NfFByvZTTQDatvQCrdGd1TIlxb96umWJ40wD2I1O5bh4cb
qrpWApFR++srbsyjPJ4LSU3RMX+8j3bcoAiWHvnNIyIlqJlCoWVXjj94mzMR8wxX
EN+eVRyy5Al29pFt875L7ulLHX4A1yFA4Yhof9td7zszt6y0ojE4xgy0nFG16FsV
Cwr1dj2xYzdulk67FX2NoIvGaom4PO7ldQ9Mh+mBWDcAb/HvauijRpGsi00lOG/G
3FcP9cq/ZY5bUo75y7myI8e1P79wU5TQCLiK7yhD3i1Pe9pxQfhtQ2MJeF/mQrmx
GS+ojcZx5Xh/L0RHXzsikjispbAVnJo79PEpVoiNg3GyKhgByuRWfwJz6CwFmS53
/68MYYMvlTS8M6cy06toFUzuxpk0wSLAglkmMSaeD9WLdp08+7WaaSKXHHR1w3Nl
TptLN70/UdWffCkGAoBNACZMqdayHQ5rG1eNrf0TLfzKorukWgdL3WjLKMd3ud95
xMzyAITeDS7MTr7uvyzViPmZ5tCywcfRKQhJbCjJJ5Yds63A6QtLUtqXZlqKk7Tm
WedCBdta1F18X270dgJb8pGbQbRtK71PkXljo7SmdAr7HUFGc0ZmCBYk+yOluLS+
oIQsEz3d/vBemHhfgsS2oC+WzD5xXOxMpA4tgzhiImqwI6eK8YX027AjKXSEC8iH
xZZ0MQ4YnkfbgwjQvariQgBXOiDqsVklECGMuyqfvBk3pxb5DKBevpKbjLL2xZ05
/ySoY9WQW7h5Uc0+ibd6bZDQMPkNeMmBqmyWQR3mVPuiPH/OttFVxd1CcufVLmsg
V92U653tJL+6q1I3380TYr7L7J5qQn78tSBmLvMpoQUp96O6vrjdcSaCycoboFpV
vWiSx1fvGEhRucwI9i0wMRMTd3fY9Grf02gWHi1r+JQdw3Y1rcRpdu69NwEW2CdZ
HujTthqDdwLmPrbNzga2QHs73bkcuvauVJP7Q7F4wgygyO3HIvtyLOMKgk8+ulh8
5FdUcYbF8dK/WmvY4dpmk9F6uEei6G3QqcSQGmQKoXWlHRc/o3pu0VdrUZ7WYMsh
aeujznFmMJtJbXltMyvpYKbPvZ7bBtoTIz1T/NhwP4bLlFfp0e7kMvkMUF/nKEKX
m50O456sACkzp1sFd/GPo2K0bLuEi/VTfM+3IIgDjDycrPPiICNlKOIixBtHKcXg
OCQv9mnML/UNXPbH64ICKRAix4phipAftesVB5HIoCvRZ6QZb3O9JG6xqJfQv6LU
Uhn8d+jCAsp+rcMi1JZIt2gdjNnKFJu4wRi1TTvMbE64gafRevz2OtI2Z9kDYhpw
KitTR7Old5ddTNtRJ0TRD56pxsxPzNaAp6Q7iTAFRLQcHX7DVEazZ0x5TfUa/9cL
j1A7tN3w9HBNZvOZ7z/UHXdYOAfOKTW3HkxZUrlTVvoDx1Ub0WQSvKyeU4dP6mHr
QrZ7ujdGqPwigzT3v2Af1/T2L6Cw9s1WEjepkVGYZAW4votAuXQn9InJj71YvWrx
3khMemNrRVz+EKXFjLEkNMYRH83Wuhv9dOu3GG7RNCGpGz1nFpH9pODuzL+ChQkg
jdBXbH//Y9Sv2XGqYKhDRhmbaIXMRteB6OrMCBShNqT4t54iU3eGT41TIC/YdgHd
9Axx/1c1GBkg5p+vcYD0RYwYz1zRM7PmUSqNVWUXORz/O2G2g8JAu+1dKVTqZi44
4GRkp/Vs5IhUGhdZpM0EYr4YqFSwT8J/zJm0RZ9vZtQCHiAvIDmTu6lnfiJ6ueBM
GfgEiTSGHS7/zHpecklc2ZSBhhZfmKskVT/IodOzASwBQgcRBW2wmpCbscXf/8M3
cSqViWGBcwXTJEo4u6srtDkbQ+rxiCvHWbN5ye6VQJp6ewZz7r0tCJGSQSj1MxE+
KnisoZrYX6wLCuvIW0nJ40X40grU7NrTbTIY2mXmjessAetxhsqVP/wb4HSgSMAo
d0D4cUN1JO/+cA8hHucHmIA76aoyMH8lZinK3IBY88rFWqQy2ikNWUtuHiPT3Hk/
LCGkXCvgGTUX+EJT+eGlKv7oroSaMIejAU1xBW++biAieMHuONccJWWVoWjuLqKA
ejorokWPzj4jwE9YQJzTGeDyEKvvvzfbZJA/FUngfpuTiW07LtcrPgsKVnFKLxVI
2XntBU78/W2NZxJHBe180Eiaf95hznHlMXX4JIC1LwU/edkeCQbbW1F+3M8sucmh
XJ7kdyCkXH2Okp/1wDJTPiRx9Hc9ta1kZJqTtyqOG9teEEyMPD0HmlbQ1yHZgJSg
DH1N0+A7EjtAFkB8vP2bX39ACGikXlEWWDlQFmp1UIWfZEEpWJwscIHkP1lESAek
Ib0bFoI3TTsccCsYIG5ju91F/AaIzMroC57bbUUH1ktXGqQlF9m14OW4S0sSp7r+
xNN5wkJJ02qKp5FzfPbXfFCCSe4JqA+AUcVZn40w3JTosSHWs1o/9zOowySMh5nh
b+IL8ZKDAVvZ4tU9hK+LjYfj2BtqcuIMWjbgD3uQcVjjbeXTqW1uG6koGy29MGqP
jpaKFlqA6XaoAmcMXmKA045VFyoC0Ba3tZCV0GleRnT9DTwjyoUnq+gXnPyf4G7e
xFh+RSJbg9zAKsEe/uh13vKVz1eEddrAhgRdfSw+hAD4FeupqCkNbOL3pMdLsbzc
expAT7NHQoSrp3UAEgKCpbNiccti7iB/g64C8YkgZPUHmj6S4vd87bzIOwXV6qjZ
woM3cZ0Fq+skYYMtBCj+QY/gSiCBRoyO1qzN1minqnqp4+UaMjWkULD7ixuZ9TGH
VxEGuGhV/01eAad3SqDA1lKTpUfm8bSwkoO4Gq1EmHk1ze8S9gto4m7SGU8wOqRq
Z2XdBVN6HN353jR/MQLPGUyZttaNgTTF6Y4fw3UWtwObx5PYju9rL8wAsVuR/WLL
HFEwp5OuVq0fgIS+cr/M8E4sgdh3SQP/ob51ASfxVnY60C08xu1IPMFrUdbdUv27
GRVu9JGe7ENjVG6DI3h0AAXp2CQHXpFCt+EJLltU600MPZCbF2tQdLdGVNEV43kw
QFSa7JwwPRrpyDKDwqnHzOztMyFAsJH+1Wq00b9PCMPDfStNLeUma4YKqrCbRWXO
2Uvkw9sOMCTmvmNySz+HoVVDRm0liUm1Ryq7gQhAVScQZl3g5JES1m0R3EPiR2lL
cEJmkhsJhbKDMR1fMXTe3964z/DK5jWqR+pKe5+xiyj7yxQ/b8imj626ScsggQdb
A6XG4Gff++dGqmmCfL1vPFv9u5y6NMAZrkUjF+APHYXnW73DfiJ6xXuznH8YXJbR
X0VV1hjyJ4nrP6nxD8WTHOaZ2KmWgxIWYmLo3EzF4rQh6jzh/ixSFHWGG5cQsH8f
Qc4DXXAuB6AdasJMt4yozubZUwDXBh5DA/vt+5m/GCtRVbgfHPHa4p2gsQu4NUXk
7aaFYnBqnt1Q5x+6JHNMBKF+TeoUUyranYE35jMaDqQxYTNU+0WSzG9Q7pcIm9lK
f14RqgNgHO5c2w3LpIOSJDO4Axnz2xa5/ju+N69EnDFeLlVsBISoYjhsTaZph67H
PEPncTTNLHKAEB7+ISjjNd/2cgthFHl7AjUbDL7gIYVQVrI6ze0dlXyGBkwDRUxY
PiRiol4vWidhRR+qQXBZuNt4BSaA4QTP+CZ1bnjT9OfOkAe2onzaxgL3PKFvp3Ap
pQfDBs5LhEEXpt5G3UYhRMj1TcRSZuxHg3HHoSrhkQbVqNxsNsZC9Q8/7iky7y2u
8ZIVa3z3RLp2u9mGtQvRDDFKHa/yAR4+DdhS5WYX52ZGYycsmwdbAOwqCL9JdUKp
5Fr3q0U56eivYoe2X9FFSMJPSKdEI+4ZCxLjWq3AM7cxTo/uAzi7khVYEkgEFtCa
RJ3ylYrpxmu9XCVvVHEza3hrGYVQyApHzI59LJv0Cgw1Hbankl2r7rt9zTP96W7y
4ox1qiPI0wcl3U85pQNmOoXr03Mj5T07xO2fTJRmBJtyLa1nVP1wm1fsYjlqibYP
cI5T/zpjXtzxBPX0O+jpHmKYpRHCYhBmEq16lkdN2NS5K3B+y16NxOsgUL3YajJj
q76N0WTGdnir4Yl9wcepYH07yU8otTT+MEWf7nTdVki3BcxcRC/po/ZQZp2dvv6a
kAi+tnjI3nSY5mNNQ6GDSBUHN1t2lfzFl2dEgd9UiQlFHFhhRpXWDCorSbMBjtrP
zp0EdujGBdM5YUUyKU8OP9ouPVtixiWR2pWj2CqIkuncXNxszBylviGGQy+HFlZC
xnZGp0DVU9+QtMun3e3YnWNe9d0O6G90gSHst0S4yJCIrr0rQGniNkdzMsCWOxQm
oZQ1CxoCUck/7f0wlfVkLnYA531KSeQE3YGRTQWWi1rjBZEZJAWt56cgvlIx3uDc
KxulBG+doWj1dEHml0bS8pfi3vLOD8sKVN4BCcqhELczbewxhwDmxFcEE841IRfa
qEktNRiLPdKad63RkqI5OjPl1NGyDZNw61INNmV9OXfytmbUhXDko252ivy6Of+d
v0kD2g7uBbqJDHUmQOXhwvmAAI2/npPxeOQyS+slgUyjNyYhNz4gz9ikRBhBVlCO
pDRuSYK5Ra+5F/RsSgHfVQBp68VqDCyV6gz+B5AIZx3p4Og4WJ19sTiHoMGFDBLr
Wn3UD8ckvI3pVTGo5NsbYK4wTA/hvJMek+D55mtjFdpg4Du8STZjGt0CvREQv03T
19CRFK2poMZstYkuaCAUlUUNH7kiGTGl1WQQAJDR3LWV2q1fs+/m2usKACYn0Vvl
CkvC45/743KYI21wFob7J6hQDoecGcrmQr60pn0vjVEx52JkE5lHUlNECQMjGRsr
vJznCRKezdlnJskTL4g4FIGaJnd7GJzYbXsl8w/Vu1KWJtC/qc1LMWvokhmU+HbB
50dEqwJfziZIF6SHNChgQRe83JZ/XCHP5qUSQuuUa0U3d5QEvHNIQeDXIVeGsoAt
K8wZi4GnS4Lp/vGxk1U61GRfTmVNFD2gdYyTnlgEe4bFignDj2eZJZgqyA6SHqKJ
N5LGoy87zR2+YqiIi1SQkuykcA+AYvhQrIBVEFV5n/NyD02Dnx0CELztEgkTzcX0
Jvk8nKbyjGo2PWoJGdLiAFwZNYYuX0ybCEE67tMyO0obIzpacBu8D1TzoKcvXviu
5Jc8TTEOg1UWLzpeIQ//c3M26arl86SmTOOLhL+Nvs4Wtmdc/IdjzDOd8IARARZm
lSJ02ll13TozJG7cNsDIsEg3tH819AljCbKZCaC/CbI5sRtfJ6aLxOHVnRJNbS/d
YamSDtCT3+PxQqm0oI/8roHORNTWYp4qEz8NWkSMClQmf9OLxSPX4RN7SostarLA
eTUNscnYMDV2CMGDm9ch3neso+fMVZnYU0+cFByh2+tPFubysE/xBr3onDKyGAxO
J2VlSBd8IJeIaphq5wDLadgcnBVZpOVCqyb3oVe/xG5i84BujxyS8+Vzyxmd8NUv
lfdqo5298a7y/ASA6+BhB2DCn261itCgsJ+2xsJLLfBwJf4MzX3g7nvzIpbIQGS+
S032jukxQOHeczt7KsNb2gmhDxVGilHvYFIwkXgbFYwjjQmfdgK2ObsnOKopGLEP
ehQ4ehzlwSYfNekHCGY0gF9oSaqkTzVcndmt41PBe5yJyNqWaIx/HEs63w5myBYO
iXRq4lMxbe9iU1Uhva21UL5MS9k5YEpUQP6XqTvs2AcKQ7sf+k87UXAdn00BLHRi
XvFMM+cxA+nl77HIdA04ZzxCU6qKX93E1Gocrcm1W1jh7ulA7QtomCOJPxNTtApf
ByYxkIIqwDFGaGlVeMqc8wHnzffujapzHDGuElZE2/vjMMb7BXk9era2bJ5NM5ez
ObKYQO8jwhvjiI49/GYtXlSEBIHAOc0v9f6ipDS/QjAI3nrS2baoujuoK4Vy3fcM
PUmnJmh0xmtLcVjyKeZOZux/s2Q4YWI6x5NeMF3uyAK2IoGFRyib8cx/kI9+efiV
9zH2QxxyMudK0hvQlv9Z2jdJ0Sq6XEesP2F1J+rpd8G2xpAMsPx6NS4PR5MWgsFy
rZ7a/BftNgTmzQLZm9YAmwz7lYkGR11AXvEqvtfSlvKF8cXOdFBjCsGeTBkFZvrE
nVNiMAxS9Nl3R4UzjviA7nrxNYdLA9d5w0C1/b21f8gBHXTc3Ctcsun5urzSjsQ0
jV2S6SmJCKicw/ecV0KCAEMNX9z4bK5ZNVBCZ1jgiYz7ccVv8SCf274BpHS0r87S
8/ylOyIJCp0n4w64h4vNeITiOrddZO8kCJovPH5A1XeJ4ffF25mC9fh8AdHC9Mev
37oxnEQ6R1aa9d49OgXyOmnyv2otPz0IzsUEfLdyzsH+8pbYhtrnaybwbIlBe/S3
H0wBFNn8Ae4N1clgpTF/MrubgzFr4m+0NjbvExaCSDBsQ8xJdPNGzvkQ9a8v1yN4
Lm3nsJMUD49Nh7gnLs9cvkqeuqGeNwGxkO4mhGygdKAs6pKoGs/rZc8RxDo958vX
EQy944ANhBKOIBVuPpBZpj+84mf5wKe0o/oR/BiCOvlwIRt6sSgKjuLEBNkkbzrA
UVSpjrWrQut2BC/qSxdPcO8Vz0CJunhVY0GT+zagseq9oCC3sQ3Agjc/tyVvw1jM
6aXmj9Z7X8pdOOHaNUx2dZuIrzgKCn1cWARFJR86rkpiIHD0qdiEQQYAoUhStpEu
si+5HbMBJeBJV9ip5uOhMmhMnvGm0tB+fWBNgMTs26RM2is1PKdtOFaDH8TYgLtG
PVUEH4/EDIa3LecPlg5dI9LajboVebV3aDlxEkU1/jP3iWLaXKZRW3tHSVlX9mP4
qLVc17EVM0e41oTU3PBhaSYVb8/5mev0eyInUkHPEG8oKIMNuAj11zE73eCmivoU
bE21hpLNnf9E7uWZc3r5f6CtTALPVQH77e4s4lqhpxnjObN2x10vMACG2ShE3dtq
z0+hav+vqin4KMJbevpvgbDohIOJ0kX5xxNmmnUyyg9adGwZ5dNLo1BApQ9C4Jre
pSFBs7Sqs/OLSydH/OW5agdET8hj5hGUQTUfZXkM9076gl7S5RVcvbufGnJb6sLm
ewBj7oujTLPsZogZWRu5G45nAX/11SYuNuxyND3Tvm0whXawG20XmkNx6PHACFdx
/9mXKbU9RzrNYf0J7n4L3POUWluuoO7hVy/7NNYLOlYkUsSqOzw1SZXjL0fyMebc
/L5+OF6muG5gJJDpY0P6eQiOBTVUq8SIu8KqKo0U2fbaM1n44X2drx6Sn1gCaJgy
b5iew6h/CrZUcyLh+0U1YiiHfaHT6SrmvCLZILbY7KKFO5ucKNRdxTEbLH8cjt5w
7BCw/8G9rakvYlmFO4eE/+2iJaDCuw0uSUeO4xZafVpimCyLqwf7H6yBt9kwV+0A
W7ZWP5oaeqZlH8bS6W83TeHi1LZ+70OMZg+y3DxsNarfYIA2uPg0Is5bhArX1VxR
dImXgiXWBZN16zUgKi3O9WHQqe1lLHbgnUCg/m9trSoTOK0eH4UZmSchebDJvj49
SKMFgJcxFEixOH5wQOMDjl7zJm/dg9F1FmpxhD/PDwJ4vWZdfW+2NQZHwYhMZULX
Z4Obdq1IvbhxC/mFG5vOPLv8X9hJ67X9wY6fXpST+Cm/KfpqYVZGf0mU+xLCfxPd
0ZdL6Qh+njbvVS+iSFIClC2vJySR8hiOin0JAZWvcp11FKoLgVB6iPM85HnczbGh
l8GEzTT04eU9q4tlQ91yEJ+gGSg1pMiXJJmLeaJKDwFWeb78dVfvpjQGErzMn8Zx
e0h0dpf+/zuen76PuB5ahCpSwpcpb4pK2e9L7/olFt4Sea0CjjJjGKdKCxEj9pzn
mceRUVAuyYD+CftjCdpoD+Pkml20oEn+YRD+vaN4bTDt0yiAIFseSNECfQcHUc6J
qQOvFtHL5NTBVfxeAr4EGRITNL58mtYMIboShLNEkIfEwcO5sj7fBFQzHf4Gkv4k
xoJpywas6kWGcaxWrIzg/pdtzsUEms6s0+dbdf94JNotxGX6pQiMoWujM5JChxux
OsFBXSXHG2YIO0bmgQQC7K5sGt4zDiqnF2uEb8qoAw0UoFUmgYV9OHNLVmCNZEfZ
gjP5Qanz91TYA8sqeGpntmsNUiIfxi17E4meb6E+b4q4Bj1T/EnCBClTHkrH7n18
XOhxSfU5IWbx3AOYpWQbTsJrO4bBTjbeZap3n481lntJphDpjZ1xDFL4WTlXIRFg
Ve8DIVD3yE/bbpt8/jBq3tHS3QpKZSO/1o8pI6z8Y3TG+CfUB7kpFxWOf6DKEO48
Mg/VSMUQzrN/anEtnY/FVEh+YvRt3I3rFqdbdcCYLxNiAUSghwo92a/Yj13BUauS
omfFS3v0u37zqck0OT8DIlx/EcHp7D8rw7rMxeEBibopjIoGpJmuApu2eSMRjyDi
j4aT0X3uVvvQMrDHXMkgOoH6OL3Mxd7qKIDUYL6sZkgG3PPICD5USp+JsFvzKdGt
0P/iTcF6Rj8hkbNImI2MLTZ2L8K69hvwwcZRBfww0FUdqbnEBqJVlkDqVVy8oCld
w7Nl0c7oj4QUXFDxhw1lW8U8bZOeF9ZCQPRQSHOga7ieKyyfBDsFeTvcepe0TxtI
1DX+GRwWmYXKnJqn+TvQQWqOTFq7XSe9j4HmYYXJm9gR2w9rTipQBPgag5/WYsoG
KTkI8iFR7TeKLdja8SQUVBXcAMPviQMqhZT32rTxlLCo+rblWY708YZrCViIlENm
Sxkl4xUEAo7oJgYp+SNxQ111oXeDQk5Jd8r5kByKh4NTquFXgjt8CEoAEpzjQkgm
PGZ3ypccwGB5cXcKLbLRaKD9PVFArs+ks1mBmf0CwYjdvZzYLcaEJxDQ/SailObO
edTglN4SNb/5x4ZAktOfJlvYON3jjJhbP6HbSwUQJz19y/p0XD/DkYpvaElOMkXm
ZVNMdDm+DVlTY2a06l/+V9ya6SKvZGbY2OG3ozuku4LBnONKMtYn4FQ9ut0Td//O
374hkfTYnaAfTYeDZPqs+0S4krn3YUXntZQody5Gz+3U+i+WpSr19LXrne7gel5m
yzE9BEUQMkLybkmUk5TmxKmSaAAEJTBEXiYnSNpJ/qDoCkvF4sZUENUfNh0CY8t+
rhYVMGMLbLuJRpVpykIVKswh7h4hIMXOQnJj+/58LmyLY8Ane1Gb5Z2RKMscnz7p
7tHvkTTyhDE1eDby7wEQ3vN6ABzklXhahlB3d2StQJsAyPohEAo/V6PJX3eRACcR
uFkyEv14iIC3jGXHKATzBB9Mzwn34xOKRxBbtvhukgDj2cAag94WGQGhmR+oH2XY
xULdEa5JzjniBwW7EQDNb+6M3artJvS+oU3pT6kOdJlx1N0jN40Ohpq6f5w+WK3+
AOGbzvL8WhkAXy5J0l7G6HJxUJ/mi40p9j72NTQUo3BiRSNjpwTMgrE6PDU3jK+8
hIbA5yuHNA+cqg+hoK7pVl3aOXFCy8r6LK8574a8nOYFKUdAyW2Zd03pmT+RlR2N
hg2G4J0rnha1g7sOm7GSjxEmUhfJPFk7vx0JrGazksOKo10epWzArOiYb5aq0i/x
qUTMewuOkmKHQmfWe7dUoFyyrhgQlmOtRlQhAqjzUorlrJiXJypA22BqeFo6QG+c
KoDIoo5LetVNlc4hmMP9DIsrW5ilVGpGoyk0a/abma0FH+Hy+7NWnAS0WrDZ2eYa
ZSXr2LVGRhy6ZyEeyrkcdmMoTiIrHyluoubW7epLfs599RRFYy1m+QCwzXVOzDMy
uYpv8mXksnQpNL3H+oJx/k/qrG/By9H3NZECfJyp3GiiOTR9IzR5/PmOrU0UndS4
Ihk8INII0S2gayKaZIpUdoiizKeP7PQER6XBQ851ZIIYMk/J0m4jAHzmqeQiUM3/
Whl0c17q0i+BNCHDA2m4QdOK1yRDpX0NvexBzRsLzzgTIbg846uks2hjwU3Spnr8
w22LrEY31jl9EFbz12zIYrF40l/9ID/QYeBkuXDtIPaRCGJHc5JO4ds4xNU4p9P5
arWO+SETnbldYViSYVq4UFpAlZfP+HaQl6sRYR6qCtYaUPGPdkZwIHffC8Dl2mnw
nMr7shCVNvQ/o4VknyaYSKhF31TncrCjKNJo39am2SrjwT0wcnysSB2lkD9PNSts
k7hTqXT8VHzQ24bOHn58rODau7/Y+RJjXILNyWrmw6DDYkkLXbzo0e+UZxo20gMK
F5v2NVfwQ1soVa6U16LATcXPv3ZgL8AfouQnFVjF98EE78xE3RAlrLMRSy4DJERY
oZeU2vfI6XJ7HyqvjJ7KK8hYvXgmENYzZvs8gtZlQvPAeD8ri/3MkqYLkwjVoKnS
sCGOhwYUhNRthwPj0s2VOFcHn9Y2lDUQq0THx84TVuIDSvbPKLSDRkx15UKypq/w
RrVENxpDkS/ErNFcaZNWdJdoKxEkFtD3etlTITKB+SVpRwVM5D2PFjE1+tXZSgyF
J8Xd4SoOXt3HvLgACiUhMBh88gVzuTuicUccoWZ0DdUwIGsPw+6GQdfwzVkiSB4+
hbLGXwgxeJHeqmoW9/uuNIakp4UpZLAEc4mOoY92oHeuDUf5op17y11hB1n2SXcW
o+MpmD0SvJsW/qY8+w4++kuYdgIUoqy7tUR/0H/bCz8DrPN1p1ErWfL4eMe+Ilc4
4hrEwCIaQ2DWo0ppr33nZmZ1STmF0nO7L7XfONNV96qKxp+to0U8t0XjPDii2Mn4
VK+k51OcOm5KzNXnKPlX02/wbWtX4zBcwsV/QSMs2n8zRjXfLsHG94laljjU8AZu
xs8gppUtjRRWiKuu859L4OM4lwdHssPmEFWhjWD9p7XaMBrj3kDdDadVe5o7p6Nv
8Wqpg+eDIQJUBXWxz1xcHWrFXeUk22OOSG69fVRw6yOyfRHdlh8AhLq/XRahoUzb
jzI+MX2zZFcEubHB2t+KfrxoHSqfwAlrU24QQaNfStXxcHkVjGWQvufpAFDnkceZ
P4vBI3Clsmwo2bwyK1+0mWMVw64CEXEXXRgsVAlXZxzyNGCnjNBkA160VTEIUE4E
MnWZHpJwY4ygrIq7XixjUej9Oqnacy7MggjlOoxyszkT+VkqqGBvTwb/iC+Usx48
xIN0YPevxCGpduQsSLBvui+6s5nj6qVOU8UnEV/b0v2guR9MTIU83p1G7W0TtTwg
5bIyEOzjTytRE/sJjMbQCjYg14mSmjx8dMGTvtNmc84RTVhhYyuddZlpV+FFHmYJ
0AuFEfvkChvCshWsH62U1QwT4GV2QfDHjfXys4pF2UcW3cUNcX/FLSH4Mi399Q72
cDvNwUu10mOdN+tI0Y+A2bpAdX4xERh120JTeUyKqA2Y7cD9Gq3F96T0Qqp3wbuI
uNfd0hisqbrgBeQsB40ywVT6elbhh0lTqWUESntAnDlzbeMljWwASlf4ZVr7NKyN
CakE3xkOiy2MzYfg0ZN5Tu+c7QsO3NXt9z81Tj1NQGOcgMKl+FFmAkZrBBl12p/+
GQ4gwSyp60ywmqLMqPIPUMVFsdzj9mtxMXb53O6LRmHJQNbp/2RVv6/CagVyKjq5
5my5zCBnc9D/vkdMMHEzkNYaoSTYQfFh7CNTWfAPyDZ12ln6xg45FXmp8qHdKl7j
4fPi21u30amAM8zWzuhkEKBgCmkE0HkW26kudeRypoqaFXuXcssCtxClm1VqNLWN
vg2kBZYOpRGOdpbzJ51KReC4m3N+qyUauYrptGFe46NXpPRLFdOEASKmbFiB1+wN
REBVqvVPi3uZtHC/OcNlW7OY9u4+dxYwD3xiwmnLxKjN3a6O08X7tA3TNtFhN5fq
YCTJYAt5L5YDI3eqPWVR/2rt/02BDt8AqEhWOsQrYt+46+hKGYrdoWJNbJFXTju6
FFR8ExP0d08tSVUjasoM8DVdJW7SJyEQQCBz3sUN1SZA/vOrLegMPydipqNUP1Lg
BiBAAMBm2W0YA1yLzC+J57T+uGRh9YZenxwZkxMm2kX2dFoQZupuKKKou8+mMP3H
6OjwbKfygV8Bpajj/uiSPMywjwdbTiP034dLTWkVr9WaUhSjP87ucGtJKvUrZo8W
x3RE+oIj/kr9HTYPjPKaHwcleCuManQNJVsKZiYVQCVrzGe95aMB5JPEg1vvA6sy
zr/SCuK23zH2OlsQZqJyJc2PpeRq5Ald2k/gFEIIKLGcTfrdYT7Lcu63KWmy+XzI
BkNUNBhBxNQ+BTjfGxuBzmE+lEWW6McvbS3ISrPa1mlOeSNuIIpT8NyFr61frQyZ
BiT4yAvxB7UMECLqtNl2HW8AgFRGgaFxNZbkY2pnCRNDWSXSnj+N+Dq6m667htwA
DTQrWcKkeZdvhUMIkA0i4Fe5OUbkKogKMwqjD3xBtxSXkY8sNeVntIgK4BA8KH3z
GE8ovVv+kYBXbO6/kOsqtXdOZwVFUgQIKgWxHgOKzZdeM++9VkcayQJh4uQ6cRl6
4DRTXYk3imb2pRjJqVy0Vf6NiOo0sV/RSOFJMp9WbpW8TN8adxH4DZQTgBp0szRG
ESxVOxDv3EjfF356SXdVoe4ZdyQ8GpDeyqdYtFwPkCUgYJOMB+sLEYqFXHV2lMCp
t06GKsJCJ8EBdPpCRnM9eLLPH7R4CRD4/ZZA41VC3ZQEPjFXv3vMs1jBFwa5ND8w
+2bHcrojowGHSMUIVT9HQnJNaxq0hah/1+dHxecZEEhWEAdi+Xnu/2Lm6k8YQ1Tk
p3nE9lnTlSwUo2Fj2indaqC21qZRfV8MAM3/tS626Vidu0FjlMwuN7Tf6+YnJvc0
NiARPy9F2YREieCps2pZGa4VapiG/F2TUQJdGbFUOzESShdYd/ZSavvkUPRtmUVU
b43B4TiDINJYaE98+d3pYBQtNCyR8rw8roaPm2u7JMF2PnLeB6W0vBfMA+mdor/9
hKccH58cT85NIMZU7fMJCU8OZrl0rWKbS9BppelE6fNskCIaUfJihIaSB5r/JLEy
TQhxFITsuCyge1j9LrhAiqv0Gvng+OQVaLG84OOi3XKVXft/T+dXe5vt4mKHyNBD
yzQIgdyYH4WQQDAYgmFJaLlB1F9nlPiA2IQ741LColxw7lUhWhRKZKMC+H50ENUV
z/S1WdGk1CEQapkPV0rrm5KSovxNrkUfkyjG8hGg+fE8ALXMBVraJdvhr6XxLcZ5
JW/Igfi3lDBz2J0z1l3HfXzKYQv7X8uyp+mmkp3Ku1FOVRJ0PqJbGtxIlbrkqZFT
WGj65//y2btNiDClHdTlBsYpGkFD9HsAF+RB0QhrOm8rpMZtrT8VUJiLLUE7HAvw
j/ufajoySAvMaTUEMgI3q6oS3qiHIvpjsopFm64gZCP9RNKp8k1R4nnPkvi7bJci
lgpz5kiOmw99BziftkmRopTSj8HqHzCgpS2KAhvmcXfA4pg8wJ6kaHAq/cz84yHp
3xqxY3UrKm7KVRckcfU+yjYGGZXSw11KJQLUQylRGxRPZxPV+eQun9qyxprkUPHl
OMjYP4bRvlbLhM+VYMInt5e385+aliFzO+/9UM3RVJyqyr+9CWjjpy3Er9/ixb8v
TXOJUY8Z+fPdZj+9M6jP06Jn/NiPiGOTf0SZVW9EDcwmpSGTveKVcf74zM1TDIpw
RuRvgx9OhAhbnpGMLspWh/wb7d9fat1ogCOpoGGZgF5NVQBOQVHNuQmIJDLI7sCA
GDdzsF8PGBJqeuWqGUJzH0hpEsE/6+ceB2OGlabjnRX42NIHUzzuOyKCBD1Mnxwa
XAV17KupourrHGrpvLvVVudroXLodwKKfXlHrcnlD9fIApuRlG5PjgLa3xD5bXAf
X/6+xb+JHgdFJfMsaz2HuOWSegYRYpC0bAwK8z1qYo2kAcCU79gjJq3+AYh697xk
B4LQB5ExpOCO1chn60YX0jAhmvRNYxzvFheYpCqjP3qx7/yJhwGAZGVaRH2DuW8I
1iloA6GebC+mqHnzj980HBeVk2KV1Tjhb/9dW6zUMPk3Ch8Kxl/OREaqlzevERJB
9WRDtFRWU7iFWZH+mSGIfGyJzoy6uHF1jSaPQgvXsQxItS9N2GuTuPccKTN08BOC
xocjcXgbyiedD2tLMEkMFf7RULNayzuv0c/Xvv0UbOysyNLInQbWDqXXOFaPPEZJ
bDfN/Pb4HDXM10Fg8scHEd862fjHmv6p1RrUIgucfeUHJPf036hYz6NzCnbOj57X
P/B9cPp1bFBTERj3NeQEblKQH70ROtGUh8swGdieGmSktoBWdFUtPAiYSLpQ95q8
gfTp1U9eBZs7Be57xlI+KDhoMahSOjpqYXZwP85hpWKU8/JMEgaKlnBrsq2sCGJh
T2fBX4R+8YHWxnwgA62/3ywhUEUHYyLcgiuWlohzM8Hl7zdycSBouLBDQCYIps4M
WOwnPhyabWjdguMROizmIVw6sbabgyJdLyBXOar7Ky3aI+2Bdy4xEnJI4Q9NhpH/
KxCzYtPf2O2yBS4+/jxRWaRRAONXQpvNTDlRUrlqQhG5HJfuSa0fSMvT6nx0MyOP
lie/L82yX6ZL9Keo0BgQbeqKIhyF5fE45302hRs4cOxttYYM9jx7S/WrLdbm6gfv
PBBPoDzO7lzeRTv2FEmF5Gb25r+ReCd7fAbtN41wArbwkTa8NrdwL51m1hVOYyoD
PRt0G2kiOBCvQ6oce5gYqUHM5JuBnaeK93M3rViyeOtnOTRzgb3Z/1bp1PYxx4fs
GzaVuWJ/4DP/fUXAgVzG5mYWb2LDNX9F7NLM/3rOArQtfAemBuiJuXrTWLH7amvb
ADjJUR7f4SK4ee3cFnZRrfX8k6qs0ucZFyws+9FJnCy36wyUOdujWIdoHtRWFkR8
tIPSmJig1EVMZqMaamFTxr5tLdW2ihS3CkgmrP9XcislmpR1Bsujvp2GzSxb6MMv
yf0tTgqDL/IvNmxZvjG12PBSBWjI3LQI0zva/gCdTM3osuGD02l9SGZkDYIHlNUA
bQlnGQZ7+0Tf1oAbEb2SXqZ8Xfll2FYIqqxcv3uL5bbhwb36wgUNlvq0ScillCrj
dXicSeH8HG57uGaU8XfvWVPjjcSvNshPiPOdqv+0R2z+M9nveYwjWs+EDLetw1J1
2a30uc2UVwGPFEmRd7cmcHmyjp6iEVwQt7JsRnqhFQbDRD7ZwwfPvXO1SEKFTHjh
OX+AZMAxf9fffHPU26YJkdtkUVR4r92/qgLE2TCqqtcB4ngbt6ZmaxoiU1d6LhX4
t/v5DJBCbDi+DN2LoC+oOfFFuRa2g4lvfo3hOtag9YNBytKXjORa4oYOu3KczpHD
fVyCoqElgQlG98gWfJoVvb5r48Ph8N6sjIlppzCmMqNjSDjj3Bfo/yizXZDM0V/q
jEnmGkSrnGIjOPOKrZV8ZkK9AiCObAY0BTch6VCeQW2SaR1SdN+w5U1E8Mh9u1jR
ap2dMii+c0bVRWpVDndEblzu/18PcTlvkDTNh0GEpN9arUYH0+QnXhoIl2e1At7T
mchNfYsTmgoI09Of/umovQNS7eS+TwtLdh/I8pWzA9mBW0gVuRbzW8WoJCtDHLmx
D8S39L5shVQRpRBHHPwvg/rh5Fis2FvL04wJi/e/v9VsraVmebMX/PzHGjJoC9UQ
3aeYdUIGmqmIpyYgwgLtrj56JCxU4iAD2IujBrKsi4ZcHh4fUyFC8P8s5x9npYv0
ElWIvc/6TTE66x6wiTEIUzzR56MI6AEJpdoFhMGRxRgB1BR5RVBPWE6oPMYzxx9O
KoHaNaDbfKGvNSLUHGTnMhO47ZAYY2GK3D54UZS1JS36Tap/bDUsJz6jD09HzOfD
NdWDRYGMqDLBKRIY+c+gjgkBqsOBIlyOXATBu2tP2P9NtY2BbGC/3/ckz7oXhS3P
0HqPQ9r8wrZpzWY4fklhDONXmRkS7YOc0Og7A6maghxDrNZcSf+pWToCAnJaJZtM
+fXOIlpRzVsGfBMOsjTLuoBiJsjcWc2UBIp2zb1+OJkxtMth7IybDI9JgaD12HKL
3EKob/AkJr1O/VTEFWaYBeqoRWpeRxQGtC0Oj5xLUKozYuTdiRtHXlgUGauLFQVR
YPdMrqFjoXSlwymUPxYEUxCVrV7/tUM5CY/KpPLyIV1PUF/dIKzeoocZKHYULng2
XxgfDeiYZiqwGWakLlrmdc60bPpQ6lca8I5EvySBIjwNBHZ3ufAqIduje3juQ51k
sTlDemMBlRYdnduIHvRwexWl/h1Kk/N23uhlHshbAhySiHyAffbCzktW4D47JMSI
eag3f7IOkh0ffRo4M8hR1sZuDmZj7OWhQkR2A82h5eDy9rc42s1iN2F6li5ZfHxe
77g8OFCLOsHFYJ8XUfqTSznh/BfhutUc6srgNpMA1xTIJrEvOlOUYutAO7vW7bs7
5rnLDKoirJ1Y6vwuaDVOqORyZ7eG0Rk62PFhlN1Mp7ng7d/L84BwWrxPVN6qVQhZ
zSyYTNN3IErtjtza+LeHwdL83YFphI4xosMQUN2zGD5dYa3RR5QlIBxMqh1L+oMj
YZ3N3FooU5Kokp7DGUyjGDYtZLKGyN593NEAauoFICPqn7eJhBQfKOmYD9wEUhIM
F1iV7MXP2lhR8uA1uYZHqAFpb6YWarXm4bbctVAQXYX3E8EqiEsLYM7lRy/Bb9fl
+3UMiTuOR55SH1EO8FuqSUxOaX3riqInlaFSDp/8wwJ1e/F9Jh/leyN6bhOh0N92
9wMYqHnUZSVZeO4eZ+ohKX1W304mKwNkhf+Z7qvRksED7E13cwX5TgPDhCl9E6hj
m5lkzcNr2hURqjPYjb8eDojr2O/bQQItF/V7hEEspgBiZfUN1OfRsn8H2NL+Eqv+
9TgN51AGwa6t9BWdQvyTA/c+KLIqXGKA6E+ksZyA7/PEtxig4e414UKuUTgFcOTD
dLvyOWQKtLY7Gy0gCOGidmHoI1+0V+tyrjUXAK98HWzIwhg39OspySnlN4Mw63fk
N+bbq+hoG61ajt+30Z4enoIMSQB4wlyeNldUiOY3kwiTQnPYFXcslPnIbw17aWhu
fl7MHnj0bcZoUsLtLrldX2b5t3yNdsSWTGeY4e10ePlGrnGlNjfsQLXUfTA1+TdF
BtxTTsG+LnWhHR4Di8NWW1iMNjPuUf/K62S0drcGyRdlX4Q7FSkBuHCJ/YiGMb1d
yCEzpU1Yiftb17H6d8nik8uW0EK3am9AbOAqQfwpmIa46ZYDVqQoblM1w2R5vHFp
H2RV1hN3eHs0hmsaIeE5FZZ61xOYTLlYSGZGrk64CJmI1+tLxs6SIXLD2J9L96wZ
8EpLLayPXiH06QtSSPI0rrALa2f+cSEcKLMMueQUIZUBtgtCcLfAB6a5GKMqwqPj
lu55o8Ph7Xy1RwBXFULtUzoFlDfdw/QWR9L5RqcVGnGKM9g5rcBDrc+Y4e1yJ6OW
Q6/PyWGUfhBCbZGli0mYx1knlZiRBahJkMzdM3a+X3YTwkwxzWU5uYf6UEkGIoe8
Fse8IckU0zF+qGboqW7i9rvEvfBaL1LR9sUwbxrzD+bnX/CmFfTTBkQXWE0x4ACe
2W17mQuRRbnqhjsYhnEPNoukAD8zIKYH/0elyVqYcmaH1UixS9WLJoCAPWrsLUZ9
54uFVwd/LbWmgPGBfCoNqb/JE/7zG7Jn57Sfdu6ouBuGIgvXnHmG7+kfuU95fHDM
iiU88+6/59Zv7RLDM9pxOUbk4tV6/8qoZYZpL+VIQ2qZQYrDN8bSmWl6I7gdKgfS
QSiwkqPeTL5HqTwM4mvIjequPwHUBkjgTklBauuTscwT66vhaTckKOqvDkfqFd9t
tx/hmwvWIZBXDQsuKkZwr9/hJNiqHd05SWHJ8j5sCxguAEFT5a3XeD7rJEdzzI91
kPuLeosbQc2yo7h6564sGcVjx0wxlx58ptRLnojnTCb0cx283wEc3m1hDyqdctEQ
fZZyGCt2IaCB5XsC6CFcaoBWK6gPeNoOKwVZ5DhubHtH8bjTO5nNuFhuUINihGOn
Z8Cu2NPceGUSi310JINIiLIXARHf4zoHpFFbDR4M7YiNeAPNet30vHM8cTv9zwRs
Zrc7tqJ8/IuqsFtLSS2y02bWphEiPyCCPo9o9z/R65kPXnAAIBfuQm+P5zfKB1CV
sDTIUp9eOc949iLPNYZcPvO2S/Pi2lvjSteGxzZXa5kJUahuLfyDMjc3BQFjJ2gm
GfhoOI4g4g6W8IxDNPryeHsMtMls4X+GMMHBgoKJf8qoEY0V+sKJkXwsiihqpWmb
SJ+8X8bpXKxK7+mBklVYjisHGNTuJ/2K1n4xl6Uo35OFwx+R4WbrWeOtJO1IVsT6
wEMCuGUDivFgWUJic2fAEyX0lScPa8+t4Dq+NmqoEvJu8Q+zMBNrZTJmxgRAOt95
yV9yrHICCWb6yBd0u7u0r6WM5/8twVJxF18i97545a9DDjZNrFfoPze4TEANfQqB
/CM0HhipjhgJaaNIULZesncwQAPNAXUEMcSuUC6Jct5x2bY6qgANxU+Kh4SUqjn9
3kjwCi/7glcLxUd5Ewl1S/R7pGm/qPdHcR7NzVt4vhijHwbsRk4CBkGeAFPe6qei
3f2QMo0YnMSdWiwmAIS//ISDZfUb3DTObOvY9geva1XDbeiDnlaMlOabcuXOweFB
NuOkV9sgBJgnKJEwKRWGc4KzsdnvZ+lX0KrqHCdCbhCGJnEhDzXh9vKz6y6rIoMJ
amipVrsPd8EbPoGdgibfXgjk/+MakoUqMVyNUYMRa8mMqUQveEs/ddYRH/MZlAUp
8d/xVVAL01YrSLLNhlwGY4jobJIvMxT+1qE51Y98blM2xUHy+bwR8p3G9ndICB43
oYqcS+7t1ZLrS4/PTT5F84JBPP6qWbOr0jiRYfs43L23oJF7q19qPSJypAu+YNgt
CiE2FF94bcEa65csUl0+hgw6jHA81ZVoCfDd2wZ6YwdWQXe542WM8bjKIjAsN6KX
G1XFCZi5XYXLaD5snIZAtnNREdvxXBghdqv3uYT6sBEx0Ij0ti2DdOHwyL3vrY5b
usafmsaFBBHdWMbYoaZCSIcCUQdl/WntINYEX+dK2L+lFew58OF99q8DcR8vse2S
TtpLjRJWFzp20tVwGw1VPp6IHt8u4H82ypTglk9qvcGz8oDKO8gAaiTCUf2NxQRw
Zh8lDsmdpDeNgsxSfOy3tmPJCcQopR5l8xancKp0Zb4pleSwtwSa3KNkc8irc0x1
w5znm00iM0Xdoojbxihmj23Sat73yk6P5SHBNWQF2tNq27uldsFLlR/SxpQ9NSbJ
fVwuJ7l9oGGKAeeB9WRRFxQqBsK0JdOzIqh6ozIMQwBZzhIJb9HGYJg2xj7wuSkp
sX/CeAJjki9eA7os/wrIPpt9v+1mjbXxiBrAvtXQy2XnKUhZifdWIvohOUWpT3Lo
2wzGFqyzCe4vyG6I/QcWZJOykvmLL3FAV2i5nMf82XsrnHwHnhp3CRrjy1A3xICH
s0/dG9S+th+003+pNwpNsM9McA0d38F1b6sslrQwXgaYgL7FATEu8sjlqTt0BB2F
aC/l9HV0MR289gZDs1ZIEdx42rgSuRkzdTpesI16iWtvwL4S89bVz2Hyza4XCgnl
eCYVnG4xxxli3X7M4cRSb7TTDprh8BdP3b2PjS4/3XTsbsUw3cJii+/yJIKa6AOK
Wmn9c1O/YJHgkGzhHRR1dkxq4hnM9JQnVBddVojPERLrmZ/hYrjN5KQvYTuHluVz
u1uc28KBvXJVubNOtisf4UM+BfXrThwaCo/rmrEU2JFUa9/MopW24yF0sAo5X1m0
54QTDgO4WALaPXIbj117hY32xoDWqeRkayfiKbyez41VLvClntVKQZfo0i9VC2S1
7xb22JUZNZBfx8M/jr6Sa83OcL0eDZSqMFRgMoBYKUwEoSIZNTvWFsLuDXrjMlCI
MVHRdt/VeCAkLFv0qYBp6X//etL8gaJZkhsd5cgxd1nX0WYaoQFopMWd+etT3NKl
qGAcv6c7YEFsopV0IGlzWk6EYirxNkZIcbMoYKfWKZkhQEsmuCQO967IATiT742a
qJK2d3YEDhD1bvqdLY+BOBqtpMfvlVKJHKNDKYI5C3w6e9c3/IUGgfi7ShJrLT4r
HQevmNQ8vzggF6xDYq4D08ti3Yq1m49U6O4QIH5lmWWssEdhbAU/Q4mSkoDm6zXx
vsxQGXxMeMh7jqOcDP7WD/jZgdgKTXalHL/g0Hvv1brLoX7lYMB3xiGkv6pqOZkA
UQLT5LqNXWz+mFfaiZuAjEPumMYVFAyiTZZ9xBH32O++vADHWFP7zHp4iXrIDWP8
RNxQvntAfF5sPz4EDtbdyRr7Gkml1Okd1ndNFUmZEkCxDO0lOvBE537zjhZf9I51
0+HfSPxXawQO2xtm0lao4rTPawnGprvr4aTUvP7mUaWMkhMsHyxi6i/lZLuJBYFL
LRPZQUbbx0Kn+yVVsXcf9FayqT6MZxSIvRmBhffq8RC0NLpEW4gZojwTS7WVh9lt
m+JfqTtgrs502azf5bTPQk8pRK+LIfMpe6+URkPTaEHh7ecnxYtCjHhnFoAYm2NM
5vvhTEhj7CewR0WOWn0nE6OJLAl3h0Pa2agDexSQ3sTkX9pKDJu2weXmui7xBJon
lSVvP5DEson6GQb43HmAyVwxpjIgtXPLrcPdUJo/daLBXz1MDYZQDx/1Jl2QQIEy
G7ud4DR7WodA6oiEidxag9UwGmNUtTAlfh5kbkbFKaW8jALuICtOVNmbCa5cUmyu
OSLHh4WjihLgMeWus5eQz825kS5pjVxPx2kQ7P3HQOpekFPu84vhK1LCMqhXljxA
UQzftIiFbpjlJHUNxvqsH4+TZiSJIobpztBrHwTr50VYaRujBpBJtfV8a77CYtJX
cI3RJ86wxPMBWNq6P88r0atC1Y+/SZxd3EOz6L5VIpDue8iLLCyfg8ZQ4Y4+DNOM
RlIlUdNfr/tjOb8sdkZDneuivIOnu7xG0dQphxsWx5KLIMpvnDYF4dh5lhtusaav
OCthjWov7awY6FpghivVAP2GqCHnJqYZp9ql4ptyHbm5V6pLLM/vhDpIsEl/DLcs
7OqdU/TEHAZOx73m+PFnfqMV5tmi8ER9eGdPD1ZSzZuQhlVjxv3tNNyBweiJJzhi
yLF30EOhOqtsoJGLT95uO3fvpV+tkXpPB3k13tlIYnNYhWS3SqCf2STWDULH1Mqr
7Y880BdYyYHs6OnO/lIXR5URTGiBFsMX/7kwRJhVm5BCbFh9IfSmp2Jlo59Ic8vW
Pp1pbhmiuY9y0FWYOCqMWOrmL2JhmW0adzToiRGuQvaK5M8wCJ/ybRw/9p1FECwZ
twH0alvGRHZlZbl1vAZee4PrMhUfk2fVS82qdCJ+GqALL2ZD6AYic1EqiBKNWMvc
EYrigaPRTXyZSqDGA/W6cVfctozvTho6PyBKFbdxlE/HXmT5DDHTXNdm9ZOvpOQ2
goHP8AZveBZsPcCj8z5RRd/HeBTGbtWA6Lway8ktWH3PNtwfFCo6YuKQN9CdN+0V
+CoIIxN4Kdw1hJhAHR2FPDIp7WCGLEKxpwGIMz5Ta67H2CzSYi0uKyOkTIL4BImO
C8+ZMZcrTwAUbYbzknz2Wvwum4MOGBqqws1qGD05ZnUcwEsV067tMkc2Hr9hPxZQ
W/lF0bWwg3aXT7vzu2pB4tBrBOYYMwUNL0l6Lhe7IAPT/DJfWW4PzwW6mo8Qldi6
fBX8qX/38/diYcn56l1fJlT0w+z/LBxefSbdsGvYmScfsYRslazjzr9EFmo5qH3v
bFB2dnhVcsVqLgUfECdSFfOm3NawqpQ7Jr06xkBmd29mPM1MUgGX+hcaFGkNVpU9
Eb5NqVaCXT0ecVV5FVBlJy86OvSYUs58R6vlNaqkzLxVO+ZLCa5eD/8t5cs6QMnn
1LoIvqWIjRYZmgxEjsYE7HHcdFDlNC8DZqNOsO4Yj7iehpE94WSyyLgPYniJINOn
FZxdRQjLc1syMCueFyLc+vFZOhIhw3QqTWW6ILtoT/WdV2HDrE6+ky3uM2YT+gzF
om08oSZPpc+cyLZYIG2qaRkHx46N2Kvv9HH9LPPY3ose1zxb7svSQQqN5p0+PgLg
UJ2iMMuiXFJJHT5JnWwyQlo46I3S4v1BgxN0z9XqTJZIH6fK+8XxaH9zulvl8JwH
K22JdoqzTbw0gzQO+MUrhGQWPHxVHgsbOae0eKmO50/gI+pr1cRvTPP6RoVucemn
Jxzz47e8d34LQ1imIAZFUHnw573yr18osj10Z6TSb08176+TU1IO0nyPg3uAz0ag
xtLY6DuHhe0oBipdEu2o9UgFbZpzzb5uaIcr6mCGuDRf+up79F3R2Orp0iqB2xgX
t3HHTIlKQCSRNco4G+wRygf5YS/4zDt6LrSSVpazRQJfhKUmgIO/7LdH8s2wfFHw
QbeDrC+qcYnPyNymPMTooTla6vSA9G13/b1/rMjEGfL935lil2rGg+jgGr7Nzk86
cEjlsWwSFrKcTE9rrQ6QfDXVWaIVrkOaMUU7Kj61FCfYw9hFMnPXnYHFL+I22aud
38y/6TXbS3eH3LBd2bWBDRg7GzxDoafvymzeNONK7fsYtZ3FOVWUs3LmYHk+iYZP
xewn5nDzi2QltEBqPrVq7Iso1Keo0tnvfJLVoXhgKNbQdwxqrp3MEFx+j3tgL+yi
JfCE5J5Ya1EFcXPoymxuOOT/WjnUwFxh4zhOXZCy7h54zMDw07M6nOqWtZTGvFEI
Tb2oggsIpE8cn9nxLUsU0bKn+r2NnWilNqXI8cN0NU2kfiDEGTSvGAgQAy1yGEHW
TgCetjqV/TrtFYlt1fwgpuxoLwZb2L7tUJGQ1M5jx19oNxxlaz0dWqnpGuh1ZcdE
3EHjj96CJ6UAmNZLYHPMrYN6BnQN8GKJix9qOT13wGEKCLWJdG1ykdy7O5vSnrpB
/ctMb4/LJPMOGR/tmvoekaj17+a7vYMyZbcTceQK+MILRJThgPfa2tUUgkJ2+h3J
/XMfFzTDayLsYonpPMVrUGxms0gwZAMUAvRr4q/DVx3uEtli1iNIxdn1pE5DvXMc
mZ6cmqa0uc8rjAeczuQurvXdehw3hJphLgb55yoT+mDtu0Heq6MXp1DOu2wS52ai
nY4IAdWTlGvUlIpgquJjmcP6x77TwoqYGhjXXkhz2/ZQBqanS2zhoQ4iyv+J+y41
fYxCbaBrZKGEpsoNOT9DH3casmvX4HkuItQneKMoEN73jysab9FAD5d21BN9nB4J
6P38gF4TEzXUtsuejJUWUX3kJcevqCeMrrliO5T+68QSefKiv5Aza5V+ACZN3CUW
/TAeiFyuHQBalXlV3vukup66NY85AdZ8NayZMhRsX650y4HzR2pnED8gx7Bmu112
a6NovGmKk9m9qfSbkdnatKofsCD37M4D+h0gYDkTFvsE3REShscBsSFMKItJ8rE1
L+iq9ZXPIyHmDypQU2b+3K2p3jDELV5GuCZa6yHAmMywebw3AV2BPEhBRpXVssJh
I7UUgJtC+spy4LjTZNOOp9nLERDFXxNfQsNtdL2dGHH2dJnLMWQ1h+6rUDCB6waq
l2nxsObyjFR0aSsTYiF88FonlrjQTgSDO1ZTpbJEgSsJrPVXcHmpmsGhtXF+sTzx
tHw1d+b76r2I/GtmRokh5OeN8E2KPNi7azCDp63PLK+JdVOa9B5Fv6HyaUUcpusC
PvdmeCu40XVQG4lKxbkKTY6Mlu3T8GXciJWq09KIFZ3n9Z/weAJx8zeeuNyIxzcH
wMqL15nDtcGDGKy6JtYLPfs+g20jChyaehkTASAcVc+3o9zDObwLj7Qwz3CfDh2N
mTeScV56gk/k64dg04ItmxNnUtkRDTkMYqYQNk2wU2rrp8/cN14lhcTkqca2TGgW
JkPHbNR+NRj4pQCF/zYaTJQiwaDmn2cG3oUC8RX+9A7oXeevH+DxUGSryCQKn+x0
1fzli3NqlDmq1x/j6DhZnYRrtWNULHOaQQ4WZxPxZdRBy1NefBlwT6FFxmo9i9iX
OFAV8kQ7gYPd89EJPUIguVYXUOpBBETiYdzY0uQRm3R2yjeXkTiQt9BPVMMrEnoy
uRJoAhMV+6MrSKcQqfoNf7Ap6298iMcEa8+xTGvf2n1Vqpo8SL2D6PvJQkBW3j6k
RwKb0DQmwe6uOOCOzUg+99V8OdKZKSkyi5Rpt55jaUph348DOqpbH0G58EvYrg2j
X72tVHgeKyhuYcEb+eevYaeo1/oTWGCjJp68UspYsSCWuIfKgCAwvlEU2vOQRN9M
tcFPHuIwv+yXKlxfIqG+gsqd3E18imp9jwNBZumuI7C7AgPIg6flzYWE0LZ+3XZ2
flPwulqDeHAUG8tSIl5Ox2eRAlJJzadm5kViYGBXxrg/SzPNeihuqhutHSz0u4FH
PgZ0gWrcqodfEDZ4/6Ppf2B9xdGbYutXrDGrRsCtxewHl3fmbyWHqcuKgOYS5zTX
NdDXc1bqM1fanZF8A9QpXgJ/4L+xiy+Iggf27ym20qHERpc3NUE7MZmbMtj/Gaao
fJXxuxoo+Fh4sVCjwDcNAUGWjWhEinDNMJJMi0cCOx5tUuk0SCzfIha7QGsWCa4e
6MUxqaT9B1yfmlKj0hB34Yl+AO7LGtTHqaqaArwPfHNKPOwOPWTIf6sl8oWW3QHa
qCQLWYBUiXhGWF+52i8QJKz4lcEugjv4et0SL+VtCaYiLLPz5xB42j7j+9rdm/8h
5+BRNTc+SUeSPUsAzvoGTyBZ11k+cE8SBiOaBNExgh63b6BKauTqX6kFnxoHvGFW
uVNqptv5dXUQYjHp5rQo5xTl77VdbqgwF1y5o86UAfdRnApdrE8wiC3wOIVL1e+O
hs8Pfs8U6H4Erz8q71wKl6zm5iE04Op09rLVTS2+wDtwImBzy0NyQd1if92y6aoZ
RVHOOL+Ll0r/LVJ6v6Gqpyd8C2uy3C1cK1pyw5k3X22tW5U8LQhvsFgxWDUwaUJv
GlF/RKuk66qBPQnU4DxX7f6qro9uWgDiq+zc1Nxog0nfcPjMyAjQp7qaErRGG1Qr
jOrN4jD7uCoKDq2ggk+UTK45c1qctzP7fjm3ZCbAYyTLYZIrso6/KtxmNe2tfQeL
pKJPIDF6Co0m5bWv6/XgIKAXLj/9sQ1hhH0fp5qc7iRk2+5Bw1qfld5MRim+MuIF
Nw9+ILKAxQ8qzPO71FNHoeW1CY6Tn6RxC6Cx1Rnk5hI1f+m272sDB4buEd/q8izG
1M8IWwVe1J1MTLpDBGVOSSWZ5Sy5gg4kanOayKuTdc5FwbpgTc+tTXCOCq5JboV6
jJfLPomMGAL0GbVijM227h4oAFiTvnDbIc6Nwc0iuYstpNWiR6kgwdSQaVgsjP8J
KHdrHZi0Dvz+sjIoMkejwRv/YazOn4IYnRGKcTloYkeQukhXBhU3NF3ZWEdRYVHz
fhcD0815FrMOS0F81TOt6vHkftnkZgXYeIwrzegE4UXf3gUrgtNxe45MHiZWS6nB
Nxp5PeWALU498I1Uf73VyvDNWvBrOq+f0ugohejM0Y2GYfDrtIWvrRP3FdYcWDAj
yhBFsl1WAMS6IotCJ3NZTAV8foo8+NU+3zjhDknujXXtXZj+Fwmb3GpRz8htHQoN
2Vq7B8Z2YwDYsMbo2vWNJ24Crkak4+rw+snMGQvkkKrLpJMvzRFn/llm1t2j3Qqn
ojCG6BlfTN2sxHCvnR/UQb+5tI+bOVtmy+kGOdx+ZmiDbz7lH8bQbHwZ+2iQbmw+
WT9CNJnn3ZctvoLZeUxrhCwfx2mRT41P6US5cLxcAaFsn2GN5yAePXPDNOrjZ1q2
pncbIJ5wpiNTXGRSSNhl25bLt7G3N0hxqv22pPnbkBRQCpwxCChG5gE/aMhBI07s
4um2/6B6nQ2I0XO8M+HKITMpnn5Y0AoO4/4YWA03ttLY9ahGxvmPRiPIUGMQBfKo
bSgy86w7n08e+FfDFtu0Zssadcm6vp+n91lD1lJB+cZCr2/tdpgqJ4ob7QjQ3XY9
4BWHr5tQstDGaRJoFeiSurka2comKloNWX76m5/EB/AuHe5oH62sUSQmJIFKAYed
D46+DXM37u+J531AlWMU9bUZOfZeL/2azGRgjGfVRoXj6b2XGiGp81h0nsX/CIBV
XU+xd/7YXJPnvQX1IG2YdpUDS38MqtCYkAS8gGnKTBIH9b7v4o5GRpeR5N/bB5z0
KTGhYjOy/XxiFaUN1nLoqof8Ii8ivVHY/Uu6MEm7Kts3HQnYjCNGNRnYlWdmoewH
wW6DkBjCawIsvPfIShVtAKphUVgPhnyAY0Wxx59znS3UEJ8sMnc/N3QTGJvsd4Rz
o0hIdHhyr4narte3t9D2iqLLCFY+SPmWVe/yWouKveizeSHq2jYXhtmrTr5tmRIP
UKZXj5FmVHPWbc+xytwezecmiTg7WAm0vskO80ieJf6HNriRDIxxjFWW1+WOUme0
aRC/thbiD225tvzj+8uHXNpRGRR5nPHDgxqegNb3zXXqaamT5qsxYWHHqtU/wz/F
9FTN/MQQYErnLWHUTA0Ls8KulcxiIWtHU8rdJ5B5NEjtSVhrXVSsCODMkQSELALv
QLSmAHtqG94JGNqzT+Fcqx9X/uTZcqCNijyJIZ6TyaHqwZDYSnQnPxAR6G8wAFvL
QiAlz3UqIPhX4aK6Z/jp3P8QOqJJG4vgw5AsNA9Uo7j+IEjXM9crPpcSvmUFDoGs
LyWFpLpqrJIfQkEheHn0X0LCumVlQEw43JP90q/2HdgEh3khQoEnpEp/LB6IoINb
nN1H877ud9egBw15/4zGIYJFJxveGUj3CL10xj9DlCvQgf0wujsx4jfo0F0A40fv
SDdBR+3XvJPjHLS72Ug6+LvVTFpPaEKJuxPLsr8dqeGFNjbBKBe1oD5OwBqCc9DF
iPbZNaWCLTHmZ852p6yZQBWCuJAhJS9w415sR4BoGLF/WsSAzh+t71UDwTszro7O
XkewP/sU+CZAjdE6Lg9ok6QIBn8sESALI1hoVm5pGVx3LFszOQyXouz6C/ISqa8r
ITjyQTmlOV8Ea6ItlH46TMgnKjooVgx0eS4+OlAbhRUhWyJ2I8euOsfGcuc73Q2V
x1nodILx7w7HyY3/W/6qnteCT8QxFjlt5XcI+zxKV0Fk/VEV3Xr/H3tZ9TGGP7WZ
IfApDDCiUojzYo8IxxwLQ9kJTxrxfxLWQFo+TQqU3NTyLxsKJSSeUUTN3x7RV4D3
nGAbXlTxqIYirtk8rfsBS10x9SJStljU9NooInhyqBoQzhu1BGcjcOHdRDeRrZDo
7hcFCzvjAefK8jrbrmnJnODAu2UIBgS1lUHKlcxSpEFsxbFDbVG+bIMENAqsUK0M
CtnBFJmMFOE2G12x6VIIcun+7l+FPb7IL2dNBartsaI31G4K2SGiq4niQZ47/K+a
BooC3H9E0xzUPmk3ajlcKMfdPwCatIOzq+gErgQBw7kOujTyv/RyE/wRfVGY/MV/
jKf+qUwD1jf2G8guB8afZF4dEdiLNCg1P/3Vtlo+PRZfEOWk+huY9hpROUGpfk6T
w3oEr8uqlBsqrHspEMNkG6FtHc2KPAhygEoBnCEPQOjxJD2WHuPpPuhnY4+TEbOd
0yX1BBhOc3mFGcc3MUv42Dhmk8hbccMt3FKV5xqcj0fEv4xfPWVa/iuxjb6xT2ee
gNdEY7QdiF51djS43E0mMMq5KzYUSmKiWGHWXb9iKafPMFVwhc+rGPdjU+XdV9s+
F7jMdneuVLHQBnwa2n8BgL8sv/mwqgUwMP3u3v0L/EOKC3xogaT4/wsbrpmFyG5W
Zg1OtdYBlVnGqAnprYUSQ2fIyOhu0JtLnNg7f30+XjNRii07s/zdIh0f15llOB4X
KBORmxWQafFD8TLo9ppajMcrBUUtGS6wgkZZyWH5xfg0u6Xc/kcb7IeWOcQjmFNN
B4MChVWIERuVCoLgVRXqe9fAtGPVAPEQNQJ/xBLw40NxSgCCCrGscPLdfq31aZR1
Inrtp/g3yeNEs6MlqnulufRbXQ5hEcuL6lbMG2HoXqJQPHYAIt0jh/QfD3KrW5Ye
9H1bXYwfbnS/9ij4KFcV7lA+nCVht/x7+4e9OpCvI9EjRtGllLVrZaAvA+8pAMcm
7R4K8m/B1/l65rlaaG4QVwfZ7soga1exto/Ur1LoR7nl/XgmrSRFYW8ybt/D2gKr
W3futt3+kLQTLC07KUhQ0NBBOm4pUJwWDgq55/WuYrUwOYDsjYC5TNjofvRNdzHn
lxzU3BzUGYWYteZeKKi8/lSWdm15PSrRf2vzk18RDWh4PmK9qh8F1zOVHENET7HH
HMmllhI6MumqC3y1jjEWkv+Cvp/cKXzpDG47D3YN5uKqvkm6VkqPumR4wJqWoPZL
1sa8CqoVtP+1qkJbbqmAvivAY9BaLM/lnOgpuJ5gHFoHjtszqaxLvZiJObBHigqy
rOl59xApvPgQQnNBwo8IJ9E8g1kXF+2xfV3BDmFGdoN2FTWmrrk2LrSgyYPvF4hm
LylNgDAIvv9O1oRKxOlVB/Zfuo+qunxr0Ac8h9wDlurxKw7emoxYwD87JJmuzCBj
gD55V2HG7X5xBYHRAamQWEf7WahRWHYQtmomZnx/1HTbRH6b8JNm+rg+y32bwcdk
x2gwF5JC4oQvQHAXHJm7UdOuhx1Tj43tRnG/JKlOILbxRwYcUl8rV1gS1Cl3FnZJ
x3AEXyF+FqT6d2kECe8zeZnHtDMr7ipFFrlBP6b3bYOC5ynVIQqCy93Q0vOZoUdZ
vk5RAY+OVccGBwEzEeqGUwbmBHzJ8GmiMk6HxXE6lQRNicchE3mZTL6BKO74n57m
os+aej1LGa7aM93htm3zCF8b+TFddvq5Q28fL3Q2ABI4/SC4ZCqSsQF8zUPkQXOX
x6oIecoSgwc7Hy4EoV7rmlMz0Js0PMQN13fXyqcd0hNkBnI4/Y6hqNc4UaDspN58
zxzqQWaccRSDGLgDnbmHsAPpcSt0Ekxj8j0InO0oNk0KOgHguZUXKQFdK2Kv+3jl
0G7p3YVmn1PkAq5icG5E4rLCTKzd98zif/FrdXdEy8y9w3FA6rAwjwizLDjG94w7
aMZxy7NTVCfkHrKJZ9bI6jR8GGiRYbx9X68pZmnfH3mayJa9N3w6xNqU9MbXuXpU
8V3xUvfcrQfpK++9ZPs9VoDdQMacSTiGkvgvRVe8uYtMpHgN50RozpqDe7uu3emU
NSnvq3GvHKCh1G19Kuc4HuB9aK0Y1l6Wu9oi0A1QqUyFyZ4AtTbgytEmEuJ76HRW
0enVh/xLdoyQZUkNjyaNIOtmR9LENbjeWVlfaxN7w9VYVan+W0UkRlpJkbVXVK3S
HrX0M1HOVDLvOL/BVWmp18+VYYzNkh0/qHTKaH8jaiacrONSuEZFOsrwwSuatvgt
hAWfsQcmPJWvATMJbxkuWt0KBObgn8Ob59iTnTkFiNy3+TJKH6SeINb4fd2VcBhi
opaSmkADWeVsLqH6Bdum77DDlc+R8cVutfbNEwJw6qwFTwxMKb6f/Pof66R/CPmF
A9NfPllLIsBSNKq+Mfj33kWme0Sw2CvD3YsA/SCSDINMxEK3CQ5+F4V+KmuN8rNk
VkQsQH3p8VLVYDgoOur7bNhcwlYn0SWwDWPYF+SZdLxTgYX3ldVrJ2iGskY/TfeZ
VKi1MkFCiSakkArsUJoI+GnXSMlS97F1McdsXPDLSuQHyRKVNRMbkONoTW3yvdMj
2Wo9zoYoNrz+kYffdqoNxpaMZZRPl0qHo2QAD2vQoYwiYToCe74Zk7KFoAqiwEkF
InjUtFwPkYXuNU2x93iunJ1ypWcBVIBDmP33Adj+ra4QilZbR/WnJgkhbJGM4XRi
4q0UllE7bYZXVrAhUbVTlwtfZzJmRA/igPHEOljlkI63s4VOJj7LQlaYxfwMvwYt
Sn4E+Kec1ls/OZFw904ciJjdnBOKdadaEvJztf3N2QBesYxdCXhftj+DUAhITuPI
vY9AxkrtdY/5IvNcWMvV+Er75waul8MW2AF5V847BrcwhdVcLKhsNZwcood474wf
2vlLG5QwgRmAC8P2BD9jZa5RyCemPvd/b5yHovPyG532RndfP2JAmStmHiZMgrJw
m6bueD82lmWAGvmnJXXl6+MeDHr9DZ+KaaGC8g87Oby61S3jZiinQRhom/vt+8QB
K5N1I+mqAgTRlf5bqqYGhu64NnJm3YG4/GF1ljRH9Hs73yEWZpBb8V6tlWw/p2hY
aa4fNIJBQY+yNo0DGQlqBoD8whOOf887dc9hE7dK8CMMZLhwcczyww88OkL/y205
1iPNPqXpKWtnTs3P+lwVgXFLtQ0xkfI+2B80TYln2C3I3oA+KB8APIijV6p2tNju
XJeV/FyEj7YL0cCd5CvXiE7P/xm7t1ZxiHyoMWA0o7xbFR6E1WWNzsIZU3umNpPU
+P9U8EBbPlNv1K4lMQhnhAqH1arbFWsFCTyZYxhvGVN1dCENed3b6oSC3vhBFbKC
fXhyquBp4V8oj+6QV3nY6kx5ybITwxNh11mN94E1e8OcaIWkmwLlNRDCILfxyugy
XQCXWrus50WyQDsEyE4FMot3X4VeTZbCB8HTukaKCHrNf9gE1w2a1e4nqg/Jzeg3
ebWH+T0A1Ovx4jsk/LonGb9VruHsEPliFInGwJsutYzsZIHlDhDYC9hzC5DLZBGf
KI3kmTS7CaCMW7WFzeSE4RqJEZKehxObaB2DKEqIhNB4VoLLQ8gvtNc45v4UWEAE
5jCq3zsB2kYOB3lI6wk8jxmzhIJ2Bt6Vyr0QNfv71e5cJ8s23C2h5kcs4LZGQs32
wFufZgnlFWhiOUqCTBsCoNvs/sf3HbbJIJl/ppzHUfILlXDBfYyCLhrmWt0n8WwK
DVJ8q9NqKZ9VVogfkjqhxIT34AEw1dhIRgvhdbnqVUo0KFMU19MtLGNx9+yKRMpO
3B/rBqEBOb4s51da6G/CpSzink/SWVBhaGrfjsYJcy2i0GAUdMIKiviXDwY3T0t8
6yRWwo8x3SOB99kIa9iWBDsrC9y6lO6g+EpnXChX9rqL1ictd5dhUnhj0eGQywry
wB884dt3yL9JyS8F5ktfZkJPXfgGozdmN3/1oaCU3Q7DaZ1n7xcoJRWzJtg2bukZ
R6YNd64GjwFsY5C34MOXjuXMkU/a3ESIYVQGjeWUi/XtONp/HgHgEo38YrBvpFFi
m1Gp5Po1Bsi3tt1dsqZwiZIXr6vRxSiY1CZTvNSjOJi52tKU3trO/3dU5NE6dCeM
kLcT40akp7n2Yfjb02TiVDaAXYjziVYmekhyH3LG9TGG5UuaIRfT7NxcJPa8Au/Y
mldjvczmWGFcZ3VbqUynj44GOyMhR8L03Z8yFLfRCS8bzsmc+ubBAylUJFtuQhm/
02VcqMkYzoPyRDA1wSvO4objpIpxytLFtIxD3FPf8dfWR86u8rlOL/CJwShmRfb3
18ZerrwNnsU5QdBe5DIFJG2yLap77sVH8YhqyIyswuuwgeyeewRCF2m67imZKxVA
3l8+rK1mpKZcnPfnJIxNo6xhUmfCtFhpsYDOwiawIJG1KjQKln94R85MLJvIJD4K
UmaUcFcTgu7W6xEa5z8SB3lj+1PCWSGTUk/jroBPmDkC3B9ExHSIHwOU/VZ8SrbN
9yuNTVYpD9CdT5wVdouTOQ3opizAFpGYbpHJo7oO6BOcQuUJcwS/7qzCsIT6y0Vv
T9jMJEZbw+pPp9bOnGvZvIffTQwF6OXpBdLsU3CMcZ14nHPi0PWtYMzzG3eoht1V
8HMMRipZQFMKrrz7y79JD8jkcEDGXZrER4+bF130N9NuaWk93PaBh262ODMF1tg5
pnyWmsFCSmy3IMP4KVlt35moIrObWOCo1YxVWx1AoQrb+tgfAnFl7tuwK7iGAcxi
2GmieiSTAbFrs6W+6+iZpFasglBBw2xdFXkgg71eG7CmSLyyltnRZGZD1BL670uW
dBHLp9kaas2hmhRZwD7StonMYCcD+BDKmu7Qjn+kgzDJFEXeNPcQB8ISdrHJ8y4y
Bam+0UsZCZnvOYpqKkoZOj+uuYpbdt6HmaGiAW4sLXcfTPfRX0o4kJUPIhETcYF2
+th/+YRTZD9O9JdGbt7ecg6seAEeQJN5Fd/5y/slkoDcfDrjcNJRXtWkj4A59FWY
2epBgoLg9xbD/6Hnsc+e3rOznLLaNxhbT7K5kZd9ohMsGorBFeX84VXuYxwANNl7
b8iWuhxXzVgSST6wEg8D74rtn8+z6zn3HP660Q3lBTAKckinLUV6xcHsKRPzcucv
581NvG45uo2VGiT6PrxpPmZiUueGuRwc/7wMfReWqynMyLLcmRMf0QajznxPNKlI
RbUPp3qY/+aJQ0Ko4aVXhklCMTDi4Dg5XY8+MBuNLdKRz9EZEW/U6i2wr8wnenQb
N7nvpDnY/6l5bezQzRJ0vIDqB5Ne3qQkQu0HeN2AE1mLJHrC8hYWGgx6Yde4oPhv
mWAiOhTg4GMyqEGa4LboOQi9/s/t+33/1cfXCTf0SmiFBQi5eSRuOeYVUG69LpF2
de10CdGtqdr9obHvVmRBk1f1WCpYidwDndVwTW12BU+2pcnoIlza8J50rvcC7ax1
BifxW3FVqyrAZAVeMEFeT9B7HZP00b79s7C9fwPIVIIghN1TWJmBQH/CRn/z8gur
BgjnDJzvDx8NgtTa7SKLXeAaDuptcOoR2PKL5hOS5jfpqMcEBjrqrD4p3v/Ig9+c
1AXT44r4AJ2yokI5r2RuhGXwIvohO+SY2aQTQAHEHed6zk9QC/gRTtLWXquaaYRE
T8pl35iuubUWUzeU6/BUSXYO4+YW5oyvkAIY2JUTpktsjEkv09k185LWXEpdXmcd
RR4Le9saKdxOprVl4HgPtLvEQs+Y573BKbfpRE5Q5hcqfK1VBgcJ+RQKABmdjcus
pLkamnYBQuvbzLnl0FjPsuyEY14k0cDNMx7xWbv3KU/RW+oaUHkLsdyHSwYMCjrc
fjWHISZNiouvbmYOGvw2jzbEdxZ1JjbFGfzTBHxh7zSKvT81mVOwK7NVusNydsPC
MvXNtD61Rs/zm+ooQPJ4/kGsaM29Dcm7lwm07E153iRH1mdf4AMtpt8mVdZCwZmj
Hsvg2Yd9eVcHNl1M47neQJOx8+jdtAtXItdG1M8wmexSmSDm2qVGaNBT1SZF66x7
NnXQogOjVf2ap6pB1H1mD3ACXLELBjmgHBmFJqgzkOB6qNneWiCKL6WxzUpMtfLw
FIidtB2p4sXRSm8bWDY1sthSGCtWBb1++xEntfNofGXJANP/XMcvSuIq3F8i6aAA
cD1C0QxrmnxqHGp2g9+Egpzol+xp22xC2tkKCtWJ+WsDEJgtn+9GSXXH/bKkBMeq
dzDZb/5DDHW0i7/p8nN7QWazvE5wfmWGZbrzpKG0Uz6S3syFMMApd+gcuF7N9Y7l
OKpdCSTSt9bh5Ow9HBiXDYPz7JuvFHNi5mGJs2ebJgLba/t+8WuMg2RLiIq121Gq
1MW80+RkgLLTtLGGcmznT28/qnp7SyoFmOHxx57tFwgXqjdet2G2Pw4MgggOrLeO
WN5Py+VCRwPL6JeFAzud8UbyQEW+ek38N62AUaGW7St9Ol7Qo6glq0gqBy1gmWm1
O0+Np4sjNzuwQ7ZGWs7rcTvOP4eFyP3qwwEscfCEqhf6nPhK7rwIBxF1PdbQEuNp
0kMxinPdDRuMCEkECDu0LGKjUTvRSYN1UwKlja3iF4pfiBaGEq5lTvK9nnzyJduJ
5MEfre+AYqy4e3z3q+MBs8lqEj55x0eu2QEUhBr+IEtI4jqh13j8DOZqGGwJLa23
qn51PBQ60DP+OghphH9HjDxMWDhHqqTz4SS6JQbbJkIpcVYzCWl3+odj2JeKnfip
HXbkh6AvbBcMRrKTLbWH/LdgOFRwQyYQQ+lU/a3PJf2/OGkyCHsGIohzZ22/fnWQ
LMiqwL96e1VmX+E9lHRxKEFyaVTERDVigmJnDszG2Or/Yc1liBLYWAkA0QyXRd+c
H7hQzYeT0o5uWPozE8nbpCsNpPFOg3cV57S0DC+cIoNCBiP5MgCz5sn4wtpOMyCu
S+4CbvLzqkmiC9zT0xO+6RrtE7sKwYcSk5hleKj6NYN6+0TdZqrDJ+OARBa+rZQ+
5ayyK1FFshnwc1p5xBz5NvzM8pluAaTK+SLXN4wEWhPAbRU5D4rUoqN45o2IuJen
7/vpFpMmI0eR0gt9pOYMpcRIyZfnZZnWFcmw0p7qlr6V1Pyq8S+XvAfPnNjpJrg8
csc/EAJnpgNGFv09oSuOjSPZ629NbgTNARA9C8m9zfnhqygvxhJh9BsfH6A7r0Tw
8iQcVzQGX3W2ym/vzew3E3Nz0u1ZsxJAhBWl68q9uwUoBaJqr6PN6q2mTIEiJR0N
hs7VWaji3v8gvj+qoJfwei4zJHjEhp/1yRi6F5UWAk5Bpm9yb9U2XjUmJeZWg3Fs
oWA32QrNpOwpAST0HUNNzwtMnZPxyU0b00JOZEZ0875ybb97qBYlTKbBlhmeMfPp
A9644HeCSk9yJpIzK32EH/0m99kWaXXwQdbdJZEwFYTNMT7Akrs+75Yu96OgTxnD
U90nVKdPA7JsuOxn9k0d7pvmqRC3pbcmAXGxD4R41BWomRDk7OeV3UExk2sPk9O7
Zv15EFxyc+KMNEyj0H1OlUyH7pKm3w413FxGbhGAW+7VWNExb+udp9ADW/5kaBVT
boK/MWsLYW9j2y5lhiW8o+ej0tvsOTo3BDGEPDGCCRzQxfwnBdwmVG0XINKErsPp
OAKrWWYUDuBGg5gEjlQpNHovxMUpub9JkVZa5BAvpBoeQL6YxuLln92cARRPOqmz
vvQ1e1M2GHPpyfBhDI22QOzzrwALcrMc71vmUUN77VsJoIBdr3gYiEg/p07eYBV2
SgtEUUPVNwYa4kGIwsyFrLLvSYpYeye/YfA0epIhHqvJtI30nkhb4HuL+N2ge/DU
xnO8KVdPL9eXzGU9M+D2B91u2dtinQbmgNNfZKNbgtJsQVry/SsxUrCPySkYSciF
a8ifAXC9WgyOJ0d8QYHresglLl8oR21i2xIkyLSb974Q4cVKGZd0ROK+Jb9RQI26
D7HVUvePVFjEi1SUykBLfrz4YzjPFGMg0ASHfKXfIW1Yb9eHvtmyykV/Og5OOPLg
zuoaAF+wjRzNNAhe6Yt1sDozXJT5Yhjs8M1zWgyqo5ucc7pfQMJOzuDGB0xkuqeH
XQJ4+UNdKoxAZ//4JZv+m2ANOKDkRyHOvZA4Hy4KoWsNY0LNodL9Kn9t0HTB/KBW
jSjG/PPIYImTQxRNi7ksZcBherUHqNEpfcGfd3nSWn2W9VGvGsrsRoHD8LBh1whi
G3pOuVKaSSw2k25vCfso+/GimlPKF42Yc/ocCnygUKBWgm3/8eNXT8ch4CQ51gzj
vRbSPohyyRFYOYaNentYVbJPu2fPzSfAW76rvNr3tMR15+O/W8G/BTCNjx7++Lt6
R6SGr+j/++uHIQqj+k4FlRvO7Dli8I5SSkc62a2VRcAx6QnvXMLBEPIfOnCSIWqJ
bjy4Phd445t3J4TElNONNgHl92q6xgyYNmvs2t+ajLQSZOhPBUCD5AGp0hxu9ftp
dSzC7jDujlZAdLdejAEPUNHVDcRKPTECM2UcSD82paZFbCLjKI5xXixx2NdbUCYp
iaBNrPpNgumHhsZCNvW4irGlpevV7A0kXMRJbfg5eZfHnLi4kuqdY7c85FpYoE/7
KBqgj8M+ReJEl6oiCkZ06guz6LOrJhqYrTOT804a7ZdBS54q/bTy2XPhUaVdhILQ
jijakTVkqYnmFDh03E7ipZCW+YHlI462MJc5OEkKNV6tsUsIk5SdvDqE8J8+VFn/
oWk1jxeNBzB2eUJfL1uMXgoFM5xJ8waGwtiaDT6PEBpkxMl/HAf+O99vtEA+qqDM
/U6T1ppqfRcP7gYAKBNUUkYMHFYP6/q4macLn0S8DKTAfkD5GeWHDS+szVd7sKQP
NkAQJjmYQ9QCiZPp9oXjW7B89VZKfrRS1rHac2i+l684k/qCaRuz4E56g30Ebybk
54+j8sWKyhBl+2u7gCO0kcVcK6GPn07qXpxrkE7u9DD0LEOPEgGcqxFKkEEjyUMX
ZGzXKl5ipt9kjDiIX9fc6Urv5YWKo5gTtSOt1QCrEH+7Tsn4q9np6/49PcB5HmDX
+iFnWx9CQx5MQXn/lZAOPc/3IMR0i+gw718e9pcMWEzpbbix9gESKEpreENqhurf
GD0abEH3cdQmhh5fZfvByTYyVb6g0Mu3qMLF6SQmxMEQPeDYdQvMZrePH2gYv8qW
qn4bFySgX+mh5b9WAsTpDfuSlTB1pDGGH9kZZuXs7czjAjTOWITT8+fTY8lmPsxN
jNIj/uUrH3r7rVizOVIEEQDmz9sr1oDzY4u3CJ4fC0+v9ac2KJdrueBcKH4nO1vM
o3wblf5RG+eNBVoDwig/7E1n/tpU2kjB8y0FPvpwTO0omVrwhcnOkCEwZwf7ebfr
uHBjTzDzChrJftA7MWW4IfBrP9dP+uKSzIc7Zb4XdllQOEKbBAQJ/QRHQU+BbM8y
fizAnukxkZ/ISCB/2u2AMHtiGHz8PXD6Jon4IPha2TPSwUBhiWLCaQFjW1wAEZfT
n9wntkkkojToauOShBP/rsO3Uvoj4MCogXyoRPtB/Xc6Hr/huiBAq98PkBXizGcE
eHTVh/nqmyZ+KaaEYFr/oIK7ID1vPAFOEQHCIChOMIvJkprAFxiEljpasr5Ph5KV
F6cDFgWIoIXWI1tV+Fu3yLrJRFCDHty2ersKkjKYp3DkFc2eQVCvdjgMPsbUIBde
uyrUIHhghUNdOJR8Rd8QGbGi9ZmCKXhUYZzBX28+vwAYWvKKgu9Bjk+zSyw00uFI
ID/WBHsVIhuEv8kJ7nH6YGGTvwFTPXWtqlCUte5sQ1xhR0F1X6+3VyZ8sv8r01ph
Jk1THjT6MDYxGsXv3kaeiFZuBa5bKq8HpTn5pgI6kHbIhPdF9X/0YZz+NEVRgF5n
11w5+wpsfXaP3uuTg4xJ/YPez7Sy8oamFoP3fWGpH9Opmtj/dAU52Zz1eO02iVzl
HtInt1K/+KyJOmg1r6uW8v/kqDvOL8NEuuUZ6poD+zAnsrg0BlyOFlXkcw8Y52Cr
4amfe65a0MQd0p7uHIuBlJ/++xeFSW6MJFb8o6cXYGabb7Xl7pTgMguMn5BnqUaO
gCF6wNprvyUmaCvJI9NjPfEAbXaxy734KXC758aJSQ+b40HbS0zNd3MMRB2U+ce0
WBKCaMboOUQy3FTuCrAcF3X3wS/oejcfenwcOyvWpBUPHINFa7XTXnlAwInTTtbu
mn8TNAoShjvrGlu0L5rjPf+m9DfWKDy4Rj7YssZvW//MsosfxumhHsOiTwYXyAz1
/vgS/IGtnEpOYLi63x6/pCbzNF7ELj0aqPzdtWWvhWTLZ67Qp0IRP97SJe2Gwsaw
XBrvJ6VGI4zc3qO1k+GP8FL+HUaX1VzSmtsMbI0M4mhJPuWZmsbeC2oI5eNn6Iwk
ezT1DXymLxuptltFNOJNNBW6LIRnSalh364s1PuYULunjM9vSEQ9UsgockVK7hlY
fGamZCA7im2xIwlXlIkvJuZu07T5rkaam/Fz3SIqaHnrMx5h0z11QIPEFDqm8knC
UvegMRDcqRSJl9IUflIGZNHJrMWjWZWYpaEGQUWOOO3xmsn2FS6KG4kotZYBDEvw
mE8vPaHpOIZ1lXjO4/tsVytjBFzvomIIyU5Bc2B4axx4br6POJIJnSoa+ARmEv7g
9uTLe1zE+ds2LpLTW/HSNL692xVsHGJLpHl592ZVWyj8NXTXvgW63tV6g0tALd6v
QeqfI3gNL2YkhBSgS9riSi0uunB02f5yMqy3xz//f5aMbqOJeY0uM5qoVPhEYqpl
olk51DPxED2PAu3gfJKehOmK+KoDmEdHuhUvYYQo1PfHUw/dhKB/LBpKEpzPGu+A
fOa12DpEjcwTqAVYvRrTUslMbME6GTYyGZEsMfCX1bGhC+dtlfEjo/u50nRjtf+v
Tbv6xhfpwjSzDpbQqoeWABfgmFeAEgyCuS3HEzINyVidrKGVp7JO4vfDrlGPUxZG
LJnYP/P8C9Z2DBHiy5JslJL52wxjV6sFN7OjU5vIqZcWxIaYqmdYMnBoyadMbkJd
Na+txc4RK9osc55LMoD5UsPIJdAlqASGXxKuzWba78tYGHj/3JLAPMxKc1rJOgQ/
h2cmgngkZzjB/GRl0Owwh3VJYq3akO2sT8ImTjZiZA3ezi4BArynGYdYQoBa8tdH
DBkcqVUcgz4UL8T6eVP98lEv0I1aaHTLR09vx4wIU+gouIi6cTn/72YSyRHmBMOf
0znKD3z2D2OiAY3/+DKYyjAk7p01yPA9HtPdpaq415fGfCHEThoXKwDqraBjX1f3
8T9JPf61TMlEEjltiPfPSJQcoKfOOY65VNq7asL+ob3hhfuh5HJOdHtIacWcUnIk
ZRWAyT8HlR6jyKpG960QxMXjwiPnfo/pL1NYPEWh/Umrot3uWFY+/3dyhKcO9Qs3
tYeZWM6fmv2fY1x92NAMgscVROqCbMfYPiq+fuyI6wO5O3AtYwGLidE1gWP7wbO7
dGEhY8PpOvJxl5vSkPa90iobFTZZibI2ZvRA+5Kima+fBtIew8w6pgjuB3LFFQ3l
OORCQRCDN3su5x7joeAUHnUm2m0FzIORqkoIB1bl26XI8ReplDeTmKlRt1zzkYjS
2Vi2SfnDO3lK1N9NHBsMXB0IJWh+ONTEq4MNjxfDwe7U/Jnw7cUiUtNXdktCcjRY
e6Z53V+tHevN0qBEHcuZqudpAsDtQfJ0CB+M1e0nvXkou8PMiIHObx/Kv/C4LW5a
WT4Q1iP6aeDB1JmKeBSNSN54i01B70/qYgnSAqf17Fh7tsyAg/7OlrsZfGn2z6QD
Zd7N+komTOpnEV6KYzyTOf+B1rgmBYrCI4/EgDtNoE36X5cHMQziPAq/FLlnpl/t
BszrKekyrVH891beV5lvWlXJuEXAjE0oJshlhT4Gwn8osUf5vG5ptLqI4Iembbf4
iCl/QITRbpcSjPXffj2S86zO/P/Epefno/QYtjX0NQ80LPfw49pbHvgARtsvliZp
xCoJ11RKlIpQMhrhqzB5jpCbmT2XNgmsPi7qWW/Gx52Zi46TM1U47yR6R6oxhtLR
hh5+vPs8tzCDrZwjRvOMmivmkAG/KWE7Jg5RADYPX5WuoLzkfV9yIhbebZP45icT
JsGlup0NOEmV/N8gJ4tW2cMbJ1SpUB2k8eN1bYmD+aF2ZeGmj37kNHA/b7WQpMwn
Q+lKGbEoZPK67xVtxX0SdkFs03+al76HfDEIwxMXeViVO0WsDYmjrgh2z3rgx/1h
OCila2q0w6qRjHXno/RgrADFzvqrDN81RB+uGS6ywMW5qBGllamdTPGviVDS9fEk
3r8o/HGTSCn7A12jihth+Fb6g71agqsRQJvk+UbMXesr+Iawv9rDJBLNN0hTTs8Q
HR2reBWphz5Guwg6/hKAn2buxL0k2lQorYrmMo+Lvvid+YREBphPalryvtK6xObg
zSKzmPYH3d8Dy/HxbjLULKYkkbqEY4NFzfKLFlXEvFmeKHhX00KIc1Ofa5t+3QoM
UEWYTqHKUIceSgyMKhW/4gpqmvxmG5cOvFABl3kP59++PmPcxWWW1RSYjEFEOEiv
Goybj5xVl40T0m/Zp6o1MpQX1B27evrjdcsb5oSrykFWzl1IAFZYCJfbcil27+2k
lC4L5TsQEYj42I1TKbwoKCE3LNEFjXVSX+eUOxRhAjo8jLGVHBVOwrpIj98vKXB6
23PXrxzZAV2TkY+GltVw1qoGU4NXmPKpIvNnhW9HPoqG3C4Ap6EODYfHhXS0zmX4
4n8AJz8mSPZfexSEw/HYvBkVYl4FaeKC8H1/hcLDe1cV+7hKEIoFqXyrTt+RiQ6r
Pv8NsAXPDA+fc+1jcSsazbPWUR1GwoSobeLqDGghq5rwbdJ2TDEoAvgMAtf2sjCI
gAXvpEEJpjGidTQi6wrbRbNJjR3HRI4VFbdFWrvBbua6K0PDs6hw6uAY45eHyBgl
9j6PBFR8qg/MVZkBQqBohDLvKenbd99lsBveFy4W8p8IHke3TSBOQoYxecfZbInR
6OG/X+cSJL19R9yU85ceapiI7ginrU7LJm6PoIZHXjdtZKvoa78lrxXRzaZx57JV
Prt96AEGBec5ERWbNpq68GMuue/xHEeGx0nZjPuWy9wlJ0zy0mE+C6HCpZmD5yVr
hJVfa1u2AYBCjjGX/4wtuLnBfMRT9xO32pZNU7JrY/KMXvb/ZF8phk5H8HLyR0GE
GrfjnPsngYiytw/KriU0h9VJZVFAXMrrpqwlcbjX7ZAPvVA2Z3sz1WPyyE0Lhp3X
L8u6ZNLrv4Q4BQT4AjKnEn3KSR+SsJm4yByhG+CBqKoYHyhbT3gOizsxk/Ey2SsQ
QJBNelNYL0CbGoxMUSVcZlAYjI4TDnchEvD0FcKsIV7qQOue5oZii+OiALnmWk1k
vXESVXX/fXs0br0K4AIGDUFactzlZK+E5ts/XD0VYcl3PobrqX55D3xQFMZcIS6V
o2CTwnNs725/eqGS+6njqYAQChpV9MzhiVQl+yYzDsAvzVrsQzNq7VEDd/rkM+2P
srMwPG/E1IuDc5h2v2VCNukhLZthZ0XAz6QnC+F7hF9LZqm5ctrI0JNCFMzmLRPr
fuwIMyjr6l5xh7hy+PldYbIyylzMUQ+/tZ8onns4oFd5ZuFj1DbGAMniQlNG+bBs
wqgLgtcvy/PYSNBnqZypQtzCt4us6hxwEDD8mLtNvhc85yfDHqaVjLalQ0InHJsg
I/9EN09ldI4ObPIhbIkp9QE5C0oOiRYX1I47j9JBzPgu8v9AEO0dMGe1cv2g2A2c
YjO06TgzHhNwL/celCqLvRbVGoGX82qgP6l7rjxgJCvKsyOPJR2yr5cwK8PEyGer
vZXmVU6m3gle6Wuoects9l6uYLUTrDyCi5ndkfVbyNJjuSsbwrXTIuPZZZ4HzB7C
oX1YlDYRt3q6TszWPT7QP/l0+WRKsbqIGOEq9gJ4ebtev2hzwe4F8h3ddVwbX6mP
7popKYI7HtkSTe80e5AtIL8zbjjmyRAdpN4glxmik4xwVqNBW6Fj+ehWCsjCwc30
s2SKcO3SyqF9rYZ3gkUeTQuUYCAoVKUKa8QvRIbTex8WNUHbG3mRXh2eY4xrO5t9
tGjCECJIh264LLk0eeC/D/uCk51WrUOYLxPRKFuFbba15HgzCARNhQZCMq2OXeZV
cK0L8oEAkFaega79M2ie/6y9TmSCyYo49rbWuxU+ORU1xmSA2IvDiyqWb+i0bUMK
3lwlfCjwEtnqfrDI2cctxBtDHFAK9sr8ys5dLyzxau2nKRXwPxURgqK4ilI4ySCc
iyuoUJDDMOeQz9hBlym0WphSbKOhnJu8gTt/28VANGp5rKn5klGNWT8Ey8csHvGW
UwvSqwUiBCYGVRGN++IAjKneqoZyWXjejovWbTcUILTwpPHLuhKotkyy8oynQMDO
WNXWgv5pkJvjJavXEBaEc19tfeJh+EiS9EFmfcVhq9SYjOrMJ4NAsE27I5H5hQG4
1X0E5yFoU2bzViJk8NdIAuQ8LjZ7SkGXh1fsLlTWTLZu7qbm8JSl0Bagpabl8Ijt
488fhiqjbUErSIkrXGGWHKeD2w77AVYR4V4n9lqLC228i5IkAp6FYzNTGhrn60sU
Zf+tAI0mfadupC9KLyG3DtzR/l36fwawJPO5VlWYVM6/t2bZZrtpG/p2cjN2MiGf
jmo+7PB/+X/qHAJKIPkCRayKVG2HdI4+aLgovXfHjpgqr6X9FBJRSfV2yuWXjNqk
v0XB0ZqKMjQeiHI2XtuFkhEH5JqWO6YWtEKAydBLqOJpcNBCQg2CqS3L5ufMgF2T
vRVWUPIIp3fHjOQbVgycl26BXCdMtL+dSCCXKiKaz4AwOyHZXS/M/m1aI7UO2O7y
ERAgIEPGOKV4xtuVLisCRL2CwenIaX8yRw43f17chW0yvxocGpW5b9Oh3g4JgRpP
fMuppw0rGjpb58spJ57l2+Dk5U8xGqHlwRtL5FaiwzrQQuvtnm/DR9FsxPxiVpMu
jzyMGvdlXRN/o+SlMJhfrvtx0JUUjW7Zvvy/130x3CUZ1Z+GnZCpETGUVymsDojz
pMuGE5adw8GdZC5FruGME7f3/AZT5oLjb0J2FwmPbYlJMsUqIfXI6kCFVVwVseA0
hmUK88hE6lp4v/FiMNJIKt8sPCBgPIWaeTfm3kiMwuWrWXx9HQ3pIOKByoruf0Sp
OShlmtmuAewcatKlC2+fj2zGRnyuWePKXsrzKLRb9fDsnt6AR12uWx3ynEoW+khU
2uSuP4opfpZlbIJ+b7QWVXKeUH9NYldwaWMz4iny0ISMRwztZo4LrNZiv9Mx4WXf
ULrtqAHZWtXu8RUa4xI30QS1a28U3sJN8MDALGk3e/4gFsDPxX6IkM9NGK/b1UG7
MXuA2MJ4YmF4RL4VBRFLNkA/yBLWSQGoZC/tltEZ7OD8qnfsljZTwrArMmdUb9xQ
GPU9Xk4iwhqbamTv+T/53RIdQXCL28YyHDmR00Fo/iWjsGbBNFBqa1Xp/O/35QzK
WQkbatOxfAnLLqsCt+2z+iNSeTy0qxWxvz/V+ECKD4PaZ92UCWQhFGQSvu8kqTVY
dK903Wznz8Fd+/863ASZsQ8fnA3Q4wfJB6A+dlGf40Xv9vcZhtLDEUEoO8wJK9gV
Qx313gmrAPmUMgG0kk1kDVOJ/+1ETJG/wks2xD7s41R/c8AV4niHR4GLemnDgpyf
ysmIBSq6de8CxFpFxykWsCbH+k4cqBodMZbVnq7gNyZ0KvEdHMdwIr+33eP3Eq9X
fSdVxh/KNM6AVI2mjqdFZ8F/K9f7tOS5lMM0SrxLW46lgAXXA4q/RtbX96O3BbPi
KekZnxFB8LcqO2Ze2OqxU94Ioa0ahQMLkoL6fmseZHqNYIdB9sXa6yuQVw+6l4jA
etmn29IKyk/LFZzqEQ7Oar0YJDIYX2wkIQpOKdZOIjP2Rq+Xbr+lJhaBRnLgy2u7
FKmKDw8mK6Xgk1uKiWp3PEjzWaG3nUpITSkwLZzTfeiNfyA7b+noAZ1iCOzwy6nd
sYyylYgGjWzCtqtxDUN+RbpZaI3LTKWmqowBsTTnEuA1o9mdhOhc69JQU2lD6fK2
4Z4NKacyT+0rO8ckh0Ytyo7zVzjgXLyRNc0VOOlL6+4eKUWMK7m8sHK8B4R2Ub3j
c46ZwqIF/rCGb98xk8Rz5uaGw3vzHBOHRGqmNQqJOZl9mRmt+ptVvzeb4VaIEU9K
dXxJSw2tsoFH2R/jdXgQ442uRVO6Wm7Dd3xJzx1Xe+BcI6/ScgStp+APbauf4Ne3
725Cul0fUVVZyxmtRqvtx+VJ/2MYMb0wXBl3/8rB8eG/jZwRLFO4rvHZG2itri7N
M106UrqChw5hV3zcMN7sBgajHSDwTUfBrOUDQ5tx79GiRFNJUAnNrXFv1/hKdA8V
a8+NRiQqT0/Al5ocF8uH3SIaVDs35nYBvXVuTQYGiKXmj44glcIcV/m5uOlfDknz
50WM2Zie1v7Gs0zZJnDV9xvhWhmdU9o7NVhrAby9YLsRXMgcng5zW3AspGFgMokW
EZfdB3F3UDq8abQjOBxd9pLPp583m2T51+CWfPMcWRxO7055cz5DWLy2ZPOxCmEb
2TNS90z1j3SH0etAiz528wKUX7PYw4Z7t9JDD3QQT4COI39VsWGYLw5aO1e3N0aL
3pp0I06VFCE96UL8etc/aGTge9hEpaGlVKSk9fsQnWc+yDsuP+qYl/1RGhI6XsIY
iBJxFoXK80D8LQRazZJAwzh/+0BKKLhAwjpzbhhd6vfP0/tyAUpNvBgK6J5gBLKv
WHBLlTofXGSpxsbDFH4vgRUJx59Ws53HhrXykKGFLcEjwRNZXbeFkXTjTB338zlX
VMrBEGcZscFiloIOJDo1P6FOpMeXjfapIn9uYAV7J7PP+5e332jiubEzkxx9lJGM
CMBan9vSViHQ4KCuAVX+RpiaynHEEK5dJD7d38EHThKF+ocN6woB+QCgtYPBs3Q1
cbJtCmpkwEOvpXnw2AwMf4g90pr4YSRSwae/u2JEi/NjKdQtYt4S3qq4Ve3MhG7u
R8GymF/g3gs5gERbI5HcdXciBk1+NdaCV2cfk12c7CuvseGMixIg2YJHfhoiy2T+
30vhbwr3EBEgSR44Hu79Gc4axtkuIK9qXalizmUvhOYd817qV+g3Q5ZqEu02D7ro
xGWNMxooar/9KeFANpfD1cFewPpRS2JlTDLb2rnvCqvvxB7go7pookDMbsIUQu6y
EywcwKCbJ6cmgttJWRFc+YLYtaEVWdt86hF0BPUxKo8NMru+AEbW3E8MAJMiRv2u
oqVH7J7nuIsCXOXiFd4QMFfzwFlD//3AicZvctcHOVPoa5K6HL2kQVemK94CfTJA
AxrX8VbVo7fPCphqbzuheNOYzsKN6l5NcYyLe1y4y/U9UkaP1hRA5zEh31hCIVWN
lwoHU8APe0xSA09jjzhWyGpImoevKQ8Fq46oBJ2IRvnG8sylyWbjZPjhY6NhsgkD
S31/xGwbpNayxG89juqFXC19+kXgzJBNyAhLx8KiCKQexmODmToFT6/V4IEKMmsl
Ic9wRScPxxYQ1PFNCYyXns7xniIHiklGFXU8YrW47e8W/FKb0tDtnC64ryt/pTu7
7f6Dd2TFi5hXrSJO+OiPHMRDFO+nYyU9IjGjqW3BR8akVKF9wEc0bjMYDr80E+DZ
sJSLaT8HeP5MoJSXHs0s9IwzMvN2QheeEnM3avYkbTu5g3c8b3H464k4E+kNKX8Y
GsZwKaf3k68FDgE+bZNleofW4Hd5eAyy5kN39e5YPlb7fmG7BM+FbOiCJTUg5kuX
EA6GvR+1XIBhXnpWxZjAlbYxbfnFteaA+Y9QBiHXV85YjRNDotL+kFxwvVPFiadD
xAvvN0uvLN3r5N5aZd+a/12T9/qWb4NMjYbhBJlw0U287BHwSxrJSfn/ov+H4qwq
161LQOT7UkQ6gjYJCPeuMbctgh7zHe7j3IY/rMa6ieOwD6BNC+kMxP2KLWhVcpJR
iMuaD6H18lSkSrnKXGtcvJcEtUzjIefkkwtUqZCn+G2FhOoPZZ2J5lpn99fmwzzo
s+Tazq1Dp3ohTcn1mBtW12/DWE4R25skO3Av6YuYVmFok9hBcJEKzO89VRdCNGsO
75TWiTQgSD3iaZvN9BKOt+8Nq9/ECW9vTud/j2hRv9TcK1bpNOMQD2Igu3jR8ryS
+YblSdrxwMTRVeGmMYeDGUThKGuufJK1v20tK7f12c2yYUPxI9v6jCD+WiJWo8Wx
yg8O7m/oPPCQSnh8m9fpZPLAUE/fdLHSE2PCGIzUSaNr1nLATkEXqs0TVIoDl4T0
7AHssUGcGBtGpub59C+ExxUJ1OPjMnl0x/bLcBZlsRtuRwk6pE/nrgX30KIQnf36
Y58HcDJS9EI4gpB35OqIPooyBAzxyw6Qn1sOCrxm5B3+oEWP/wVV5u+A7EKcv56c
dutCG4c1twpe8N6/cCluPZ9GLrq1pamLupuiFqDuCI/m9Op07nKzP7XZC4Tt5pcv
5TDhAAwNO6cFgqmOcTj2WwOpzbSXYXMr6mpYAtUoG23fGQWnBlv8+GiLpbxElBsw
C3h3EFaa6vQDnfcjPAAicn1Xt1ESrckv1jB7WxgS8H06acyD3aIrGbmtNs/cs358
nOMSxBeA2Z9H1VHolFN+kdYLzeKUe6usUmJu0QYbfop2cdGElcaMgD7tIrlftb1D
Ojy/RmWQMpmWSAoW83kIAYXyLHVjjN6Vsja5y6VyWkEXebb2YvWFv9AwsRy9uK2n
EZd1ByXdlWVmu3Ng+gcoRtmr/epu09sdrYp5nZkZZUyF0/8tnwExS4m1R9202lwh
uEjN6tHi4DFjAbdpl6L2YrOPtFnjxrpftaToyl9QndRiK7TPTVDB6/AFpAC5TI2V
ta1EzEBORduxTdvN1L9Ms/R7QtKKXenxp8SDJIXxgkgaciOgccR55hCkmEagUujs
5RhDwxxCrK4ccXwq+n75ZHHOLrzYjkytZIxW1kYZrnedKtxlJQtIxc707AfUBK9Z
bwaQGTBv1ZC49lefVYu5moxG+DGj6srxPocuTJtvAFWx/5WVTcjYC1gYaqRPuWWg
Js7hwQDtTiwTJM7W21EiagDqK5K7LdQdkDeqNm7WgtV8RN07hSbds40Z+hIED7sI
m35VAZf3xQPjGvNnYelXSrrx0hQzbLbe/VrykLQPKuI8cDNtbolWG0REAUfM/YLm
SnOpjTfXUB8vVsw+7R+HUOtPefxn706N1rLlDnGB3prcrNZosUL3sGhlHkIi2evr
4o8zPw5/Zq7oXeOgW2i/bXtB6W/bdALZgpvclZATLvOYK9Bdh3lPaWB9TifZ/27D
I62uukQTnkveW5i86BPZXe/Ct7hyx4sP0NmbrI8cyTQ5kZv1WvdjtDdJgMm20GZh
+1yQ7BD59gd/jOcH64aVeRye3OcG/TdeoTnbnDcA+ENREM+v5vCk70Yt318781kV
m1o/HxCV3Zuw4PryHLXbDii0j7W6vKk4ywgnNYUngjWwLfQXvDyWRWilzOcodqba
skrfjo7W2qdnk/xnRiv/g0tZ0FUuk3abQBGEnlxZQlX2Dg5Zl9bH0pauC6G8buHd
qq8rz4hAFc09gTBJmlAfJJVI03W5I4GcHAEoszr3m3B/TgJZ4J1Cl6Ui4deSi44F
bZo7OCr+uU8iqAYdbeRIBQFpkoG50iwgfcPQXHM8OtQL6aew9kVGWWBt8ARcZoMP
pHX+72ZrBuzr/2557xXMQlJsVFUn/QHlJ3+ik86X+8JoZvWq8ipXXO83r3Dx4fA8
Hu/7eKoAxBbBuAOlb3DbGkd83rcInhSlAMCl6cbXnPoHqyyS816KnhNzMv16rT8A
2IuS6jw8JXeyu/0Iou2SEu3dX/+Z/1Okkv9SSBi+hfyQgOCc4+UqrFoC81htLd0i
8tmKi+yn/O8Rh8b0NXDzoK1++3ArgXQ7uCBHhnVJCmyY8mW4TPPpiiP2i7CYRmZR
OpP32rWa+wyIU/AuLlVnWS+IDXnTnL63G3U4kig/IeEf3tXH8Tf11ZE162EHP2SL
vQXaeG+GVklllqM1w2Q3BgU3I+Blu+c6P3KA/b0nIV/TI1QRjk3+6lp7dAJAO4XR
RqZUatrvrIcWZJio42ewljrapUsiHtFY0XAM6rSBCKDGOg4SW5kWILHcWMoUuGD7
L8f+jHmnQ13S7c+7habJurnL4o9oTCAs9BqYE/aCSowItnG3X/7OYGY0OoYXU8w7
2g7707mhHgdBUKWreuYFUygiTyUMBwEnvpiT7YJCu8O9u1N9ZYT7ujkzP6YBAL7W
LmtEuV8iHPus11asVidNJU0Kotxqu8XQDepfCwTTOW8OpTC0C/P5ClKr2Teu8OEd
UPwvULgzgz23M0SpPBsBSp0hOBMplzUpNpw82qm0XH1fNF6yaWKJsFP70nR8OF+w
00zXAAfS/jn4b2OSYdZyEylLuIx7bP5QV1YAoBT31FPfexyATawxP3FOx4/H14qK
OE81kSD7vA5uk5sAtGCfIawyfE4ssPu3dCNiDwDu6KXuhdifgE6JQbXOxQwo+tff
LWZ+ruxvFPyssYGnW9hnOvVmWDa12/8bPs5EHRrJM4e2iwzNqpRewEJJoxpaB9Yl
9tnc1ebCXi/w+81+Ny8OHYd2GKLekXVXe7McxVCDreDAXbWHLZGssIB9UpiItd7M
RQOiQWBg8Rbt0xxaMZtxp4KqHPQIdvfafl+YP7Xe9d5Izq0E08V6KZw0vClDZjVQ
qS2U3cfDm1TJ7pkFRNNhHou8wClE3ElCYoBPq77w1tcpUuKUu/GJ77Y8VLkfQKdU
oTCDVlX1ntTRMwW3i5rDXyEuSOLHdlTSyhEweDjz/882MZ6GlkdCP07gd6b8RzMn
Pt7RaRzZdGlKENfGVxiiGqbOZMfGEwBHSEiJbkTdU3Oy1XEz459Gh4qZxAx1ElRo
Wblc8IwZrRtI7y23LbDttzRjJEMUGB2WGNyZQBXV80ipEdOLoOne4NNsEplIFbLm
WppOq7K5pu+crU0m0xfXcLivkqVVNHESQJfh/EKtZ7LJCuR4YsgjZS6COAUME1h6
9P9G+ZXhDrSjxKdJa30+zq/K0H7rep/iCdEjAbpy8t/IOn/nAjWdFk3StIRSuRKr
4/gPNQm4Al0hprB4Vlt6rcT26vY7Z9Ge6zvV3g4s0FULp7Reim07ONjUmAINTXoj
WLln1CipVdGGjvAZq04cpltIJkQCl5a8ZMXGrvVOVY7c9prMDmfVEFFBf+zocRAE
91U1YFJwOQmHhTlGjgSV3mGU3POQdnmk5psR8UbjLmdaTBd/Rkx3VGUje+NvOGn1
5tbHCZs/z2U10YhUzfTTAak3vphCP4KeQAdg72DUsKhMnwMgIo56qNQ2WxbBq0oz
H/lFfPnra9gHwrcPIQK0i+05BE8JI3Pg54HQCxb9CnGThnhEaSMN2VzjkiaaGUz5
HcIpwrcox/CEZ4DbjEBwNYn3qdUooJw+XAKl3cT5LMuUZlQJLK4Rj8+C8QiwS7Pn
lh0ud62lyRNkoxgt97Xbj7Q1MMPxHXeiZtLN/1HlFDXUhPvwR6sXrQHW0g6lDwdW
1fKxmwYInQXTq0dEuJpem1vEHp8NhwtSsV9L7k6wrXCtpnT3oxZ5ZzWvX28wrp5X
qES2b9G+p5XBy30lQ0ADDxuMtmiLcUYVdegdbhywikOHZkCR4fR4nVG976DjDA6y
Y4TPXcVwmtrK35U/JEbqnbDBuqwdXFybJHr2O4qSewpfsLSFld0niVMFrr2LEBLU
sEyO7ZXfejYsExrDJS1Qi+6p4vxIRipkgZnmeZCIG+Gd2q7saRlFhygZ6pU8HD35
yP4KL4653C7DnqTsnfT3R4ITke2dyckTu8ctzwdGIyHOPKbN+pfpgolPo9m3gShn
92F4AAelL/+GY+pG0jKMYaUXC6zTfKgBbE/M/KHxZpsLOF4Ac7w9VrHBJ87Nri8M
NeU9iiQOye9XTXlwAr/LwLOTHTZKgYypZfkRDRmru1tDpMqBEa+hdnjsVu0OqbVg
kM+UifePlJXnSaB5Qh1DjjFrXgdlJ6753SxRwYOlnJx31FU60nORppzvvBcNcPJj
SS4wUDUH3N89Q7ATHGEhpyMazmU798Z4wJc6ajWvSoDFjpl38e4iZFTVFj2J1l9q
gI/Gd+N+/mnmnPg2z4ei90+onkF4xMUqmXTkDBf1pvGiPFp0vNK/1ehFFvuX3iFm
5GPTsPZyHaWWccE+f45vKjERuZpzccBVqwadxu6TihjUaoU4ZwTjyulHdfbUoUOQ
ynywbiPhW/X7wjUOSVTxZHUYfuRa+6nUN8c4hBiIlx0ihBI4tz4rlkQ1rkL8rgY7
zgTpYgqLcxm5Q+ngrzZCmTLDzoGrvlHToxI31eUYjSlf7lGbGcAJ2JZnHElVGsqu
xq1/jw4ng8Cqui5mJBjvSAOYfuMyo9sccG6h/ye1HFwrMYuTES5vah3bfY3Qx3d1
UAnivkU3f9mCvavWRW62KJkRvjWi5oOSxbf8ONUlfrwl8Av68U1KU5mct/9TSg9k
7ec5WD4e6wGXMcUGRzhbFZCUhe668m4JFEuQYT3UZOwvkBFTl1G/dMQK5u4Onn/w
W7yfi4GiVAJku0uhrqoetcqzWg8WcH9SADTFSVCCDOfd19sRqaE6c7s6RpkIzkVs
FKAK6KQZEHSLrqWz5mtu+6+if92HiRTmPabDeQ46+VpJcEpqTNwq7j+Efc7980wv
5W4eis5nbXuEJU+2tgAgLCMgYXOKuX0yxFs09sJWJj2UvLJ7vxY2MOupSPHs9Eu/
Jrg9epeLX/BG8lYVLHYMELrQCs7G8Vb6/yFTtBaQRXC736Pi1AGLDIytEmk+oc0G
zYpKATixCA1AmWgveGOM2bjhP/ASAegAyMySnaVBthJm1cWTf14N7FkUecNVqbUP
SaFhU40GfT9zvmkBv72wFjsp3awXFe59Y9ESy83brMDcjGEzknHz+/elvy80Pg+J
cRhrrOghJPQYx7lTw3jpOxKr91ECnqrkIcBWoyLWnzxppcd8FbnAeGVHBHy+WjoO
llX5rpWwTGZM3hP9Spgy8Q3UUJmwdXWh2hiyBK8gZsg4dmDeHlezlnf9B+emaiut
zbvXeQl8wTFMM7w3sCWJDgfnP3rpTBaONIhQDMuNCPGjkzxquH+CAK5jlnXzb3y4
XXijArKeZPKxZ7qizHvMpz58lYAq1DwrdE+gEXuGC9k9Jc3hbLmnTC90kcoA8pD2
igrWmDTgSc31ayQBBb69jc5OA3Dnu2+ppaLzo7JpAmlp2vEu6A60jqqSSv5Xo3/3
jXTv0dCgWDv6N6JiY64pMrRL1wgBN5J1BxVTlfCqMlICMsagtjIxp8RHXyWk3oWk
UiGAEdVRV6VLXvuu+yt6j1uNS8jX8J368f+J3dScYyy1JyweIUGiJLkJM1diU2bJ
8g0VgeA/0mEPKLgdW3YFknApp1OuKRXPCMCBhSbA6YGn+stZIQNKJSKUOUlW7cqD
hoWi7vGz8efild8l0VcqskyoxePHf9MxZv1qX3CPNE8nYtjLf36Ct0YrVwKu9akE
+jlIHsl0+7NR9GYt0iKEYJM2i/WEYTlbcjIKMC7x8EzdbJ6R1l+JqmXnAqyZ2r8m
XouooUpH6uampvSShnOkoX5sk/LhYPKk5d2wiHwNogt0JfIpNZeKHtV52Desrrme
rvOO2E5oabFsKijzkNNq+YVPXSKPzOuOfFRTBsapetm8n9LCpjcPX8XBtvvV6Ce4
vrXig0BVloDBg68JGiJIH3teN3hFBqjxnQxAqR8MFiwEmVRB2CVw+1dQqZrJDxBP
qJBkDYo8H+aiHZj4GeglaA0U7EN6ARo2ry9vLOf8j9NXFTf1fTBZA1w0rt6uZoQq
XUiJjfr1ymc+kvo+YUx2rztii5Hz2gmcowO5JE68icysEjogbhEcqbqI8ACNrZmu
h6+ZuPp4CrTn0nXroShDmXLIetDHw/zvpMAA5eRysN0icYFyAhOQirlwbHUzxGvO
F/nceudH4+KFrs0TgTkr9Tc6HbJM9pDcPY268LU65/fd6KPKU/g9hHHQ11v1Pubt
kbQHNJuNj7tpvYMy7TZL/Jvl9M7iXxjBiqAXdCoia9gpQOvIhh9cgTs1KwqY8ToT
em/FWoS+b3RIT4Q4FPBN0Lq5641WAOhxeBldagqb1xuqNQ4lguAe947AYOw7nnyf
ee0hqAchgCItPq2Q0m420UFqucXOvSnY6QgvzI8hFfzH8UwjAGQI342BjDFVJ8DW
9S7hWdAuoS29QW7NxsZH2hLG0vjbRq1boCs3c6oRZ1PuPycU/ZkfwJiHBJW2zeBz
ckDVNSqDVcgLkvX4YwcfpCIgSz8PhJ5jOPwRFZGlO3LakcGzIAf4xwSPSicfrZlb
5X9o4bqyfOBNnMbA51vLTHIsHF8XV9fxl72uWLXtdDGNtgDHqO+uklqjZ8RXCrLu
vd/S+pTF//eFm60v6oQ4glm+XcOwko5f8ebiGrtNQbbttsRDiETEBDYX1eYHt22/
cxSLUXV5v6TSRMEbTCTImVOam6zU4ShW81Esz4JosMyLRB8DyP790uo8QUMutyU8
6KfT+vv9XPbfKutUmpztzEDIRAXvMlVJkrYXTGy7pz4A8djoMi5YNISn2GSFDEx6
TDbBl2To8yMlkCYFhinWt0/gzCrwUJbgEl9VZwaYkHl9O0DUIm7g2ksskXm0jOin
87zWcV/ebbOABeWenOvkgCB/9d7DfcGvKX4TPt+LT2sXFXSXfZrypl7vusMKCVPG
VWBvpuSdBEa1KWReM2XwYVie3wZY4YQx5JtIOKNnThw3dDrbVn+F/ght3FyqZHEp
MpDjfQPWrIl3btGEHqeNZAqag/pnFbJxT7hZt+z+sKQksdfJqlgAxjpZnnPOc0Cx
47HpejQrostwwcshbWnylPb5e+q6kplA6dWdk5pE9QmT48Q8AhOnuOxCCke8ThuT
3RCy7ChJNDRgYceEdTUt6YqhdFZGElWhAwGUzabZHFKPZaR3IFUc0HVGII5w1f15
Rpma6NqPPpRtvTKWd7cNbvUmpZ88U7H9XyfeITeq2yAXvFfVq0XDU5bjs52qSQ/U
ACGuJntMN+u2gSMAgA31rDW59c+8JU+hFrpXbK9iUGKekjwvNDRzo9ORnUkGgAz7
Ha6f7mHtF2Unt2GKWxV5QUsQo2EdQVfgZKIzlPJuFAfJdRv8m0TSfqvC/Y+8zJhO
U/MaExKfOOBkLvsjlVnhoS2sw83pyA+gGxjfbgtFuX6PnkhNkRvnyZ2k4GRlx6xr
s+SaS+Vu+sTEylrerOPvBLL5iaB8rdsKOxbSKQycjsWjcwUjZl7NzDF+q3dhz3Ve
TT3hqAcySWBl3RJ3Iwfk8fHrwZWdSIBZ1+/GFyZ5qgjiYVunmwWKd5qMGaTRLyTW
cqSx68B/abALXFuCSO/D+XHB2G+c7l2MrRlQ5Om0vzMfr4fXLNbDFHXXaLHaNztP
N6SxBtfN7wvydT5qh4w+ulabYSIjGQzLqJ014T5mrOQWHwK22+7oIxm+t1GV4wWF
ILJEzkvwMoDcQCXS0PeWGgxadMb3dXWMEN7osjhL1/h0TOIpKwYuWXKUPp2eFVMd
8X7FR8CgW15rITPkNwrfpk/1ni1HWgl8/dnyMKe+loXzASVvuRmFPjXs1T7LI1Ys
pdiEBm4UyQ8PZ+OGVUJrwZJSKsVNa6zBt9xv032m+tuGBFlUdry/GHWrHbqku+6S
42I8ctcL9zQO5HG0iIiNccsZNA/hYrT3Ib5yxa62C5ZVW6tMjOP+sH8oatzrPSmd
4Y6jTNpRcM9AqZaE85WvrbGLRhUABbgGs3uNNIXg5NH+IvdLeJMDRuc5JGs1DPFk
mdUUeP5MassoNigZMGvvCUVHZYrO1xUliY8c6Mm0FZH2Z+uAZntPOU9M6Uhg6/bK
1/pb2eUlvd7tngh2/4jqr9yvREkXnEsaOeeLCvKIvcfbwhsAuxOH+Wor1xgcblh/
dOFQNDV68tQVI1/9lJq5c0n8VFt5ZRNQ7W2HMoLOSOTzQYGMBIuDKQOf2r2FUoVS
ncw/CM6RlCyS8CtR1Kj3LvApVcoQ+pVqEAwzQ3cXldrCXad7SGGK+Dn16+n5Gi6z
uDip2weqOwSjWPVZZW7KhLEQH20hfdC3bIijYnL43RDb+J+uJcoL67lOl8qRljlJ
DhA2Ex5x3jEDY540egtlG6nit7N0WQ788fejXVrlk8SKgY1xpo+dSWqyGV81obNs
pW68PztsWtKnSk4L+IydJBZjOPKIFIrVjHAuEHzcwl00pP0e384xXleuPm+8g7j/
wV2oKD0BE1ejn9QWfFoaUvGBuoS2Ko2mDcDI2wA0WDvG3qAmO+fyadvB1nGc1mmo
cnm8yWgupveFV7WXwSY1thom2RpUQVhE3zDuMbneN+jQG/FgVQv6bcUhKJd3ucuC
4+5UIguwzvB1JpMicJWe0RAmyewNA1OhEt8PZJI3ECxqoQKetIhP2nyrujXP5BIK
dQhbFwo9bFiiko+mW65c3Nb0Y8E+F7U8U14JttPSmSDY3FeQZPwif7UT4u2lm4pF
6X55Yif3dySjvH/fUzA0NUrjD6sgoctQBP5YI4KW4fpak/6sopirLhOohmU3QgYt
gPsT6JKBo5JiiPSkkSK8uxjY4vGGAmgNrdA9VgYOl+lRq8eSPCudlOZtvrfnZ6bg
frBtfIxeB7oeJ6ul1YPhiD7xp24OKC8ks6G7uZ/WjZnVaQsChaab1awy1bZzCnYZ
seIdMM5qx5KNENOuWcSeY6MD7kkhTp2e+JVwP6RO6xdqPGg/8uWuGDcF3wvHhmkA
Kbr61jHgBsjuS7S07GRhuo4ae2oBP/4Mz/9GmcF5Bv465LClG8XLM/zQQhy+4QsW
F66jtecjyTMPtWoQIja1oiHmvbylbU0neWX34UJHOVg5bBbB7YfVVapsytdphhnN
GY/1bjFNhdzeTLsFbMMn6ojyJ8/WowdvuTDgy/rJYZsQnRiOXikzDNzbPqrSvxLV
v/FJgheLG0txoh/+mazITPyo+HK/Zj4K1f47YTlSHgGRMCYADEAnA7aqyMXX77PR
M+PFFM8WIDmTZTq1mGr/Ayo2EAEdSuuO3W0//EJ4O/A+EKmW/lVaMzorq6QKwzDe
mGD1SJQl8ZnMLPnln7Ghu7WLYE/wYQ6tSRyrNVmpPrGwcQGER0hTsuKaSXLykcdo
gHiPq13CQuFHG3jYx0Ibqm10YdSA7Lc53aB7YBhV4WCIVDfLesPnTONFxuT5EvF8
QLGqwBiHkf+NleUgy+x3nfTfGAH1p47EdDgdCWNA/mFtH2XuNQ88DRPvNKEDi0SN
nkiQeAQT7fQUb2WzL+nA6wl3TyiQPhfhY4OMs+EoG5TQSMdFPht797GPNUfHL6GG
xPJLf40s0kkXhiNZorKYV7IMDr0gVGDWdI4VPfj2OobUUVqJgivzKosqTKjGvvcT
0Q+HnLjhgfyu8UO1Fk/Ztx5kF7pRjLhH51vAbUr5ocLhChaj6nu3+a9aRzBvgOD6
UKvVtHdr3gOhB2SCcDSBOfyJMf5LF/SmAPNYsDHQ4w8UzkVsSyVhPCyzqFi0rgZS
9Um/CYOto8G7W3AWW9wJ4pPe8frpB+Fc3zycWNmSrY3yPoTxacjgKpxebKgm9T29
8VWeZCbtL5bcnNFmikIqWslnqWKlASaXff7Ky/tffzZrLhXPnlKTEUzTdQ1f+KZa
sELSxr9eH5cHqLyVQr83ftlT8A0OAkBvyr8YyYw1jyhhXpF5dK9Mw8TZBbcPII2Q
C03+UHzggRgm1pEpdZRf+n1Xi7wy+2WtxOG2au/B6equEFi6n830cVnOVMsTQkxt
cl79IsoiAt8HCcRqJtnA71bFq2jXSwUGje4df2GWKbn7BucShFkDidIRLZuENtfG
kPUfXUgG9nmcFafy6A01DdYBPAjKAsQF9TKsocbQ04t9WKePWDqhMb3+BXU4Vl0V
Hl//WLDLezf/tuL+ITvlChw0X0Dj16QWr3x6UMGbqH/39fbQCOfQpGfoioqJLDPb
AIm2OBawWAx2wwqC+DAjDbh8YRkTNwdMURjl2LmR1BTr9nvvi+4XdYpo4zJ5qftc
48djEfIRmEZyoa+mXy17gTh67G5X4jTjOa4wDNXr1I5VNp3myfLVoyJfHvQWA+Bb
CrwXHrYVPNw3BU99Aq8KnyD2w0IvgtVvGa0khDo2sGwpqPVIezdh38DfC7jr6NIm
eJ5aoGD1i+Kpjm8sgFFAe6hPyzPTotYf0nPGs9i6oszi57psjVvxtFJOj/QJM+SR
kRe8dahO+l+JbVZsSS856EhALEwHtisvQFKZmj/W0UEodP0hGzq7BLS1g+Q8wQRq
uoDApmSUT/WTSBq+U2oum1h8At4fgRmMz1yOzKiao1BCI1Qp+pwNp22QgtRGQlWF
ZwObK8eXHgmbQhndBD0tyono+EUA2OOWZie+/+qawfwU/qffFLyXojqsBXVrJoAu
9uGH8wv8qt9siZAvHQYF1pH9YKCUoiIVUFApcDnNqPs0bVYWjHc8I71zyXkasvWw
ippKEMf7y2FSDJ725+EdCsBEaHexvYNpSO62tcnedAV/NqFy7iUPJIDu0q7nQFzl
5j8yqH7xme0uVMtq/ALivdde6UuseVLeYe1ZtxJoeRuDfTu/3sQ0hn2h1oHzgp5P
/E8SQ/otzv9DmcYeYyBwaqF3jgltsX2pTlO5RBZU3anS7u2FufVyTrlnQ1syurWJ
r9E5IOPPQ4iwvsIdrfriav8v+F3JH35if423okhP2gheeor2NCbtDKDd90F0oxpA
aqiKeUrYSu8tsbAB4kyixJnA6om4ktskY0pilYpxqTsnSJmIXmE4Xc7V+XKrRUj6
8c5Nmt9kVWayIoa/9K2ItP8jYh+eCXqz9q/CvtD9XILTpMGzoXF+fFG3R0XGcBFl
j+2DwFz0w45aUM5eqG152jjX4zqqKwhuQiEyFI4Zw9Fzz2ZmEJq4c8pUiI+9aIm7
73DXASrIAJtqzFa2UF4i4YBsjOfaXbemx+2oASb66f8jQIQl3fboaWQUnC2SW7PF
zAGOR4jFKkTICou3mJG4aF0V+VenUc8a3vwtpTX5S0SbepnfVFnX3IerDLlhino8
kGBkUIWh2liKHQJbXGKYyNG97OUZoeiceeZJYf6HT9lGgs+QKoOOounctqzNoYbj
t10A7SOszb7T87tGUIsgZL6uX520+po0bgx2rNqDQKrFyaGbwQxUTCB3QBK695zE
mCbEUsSVBVFGEClElXPjwBrgQxrtdZflH4pCa+jm+xGRIsu4t9elfMxf6eOdaXuX
I8VAkopIXzmXYSauFW64i7hdUSssTblLBX0kOKbzI2DFaJab51DArW3TvEKdpTdz
Vl80pzzBxr6IBsnAq6vz2kPA2DC1ceJVxpfppIuLl/8h/Oiv0+XrkMhtsTVrx/Kd
CFHKuLGHEUQUPlOpJtYt4BVlkEknHJvHimHGNkWVia/hrvxTaIinxlSvpxJEWbU8
pZCFaPGrJfjMdRLBkQKCZK5p5mdSYoHg/KGJQF0iQvxgybSIQm9h3QxY/S5vhPWc
Hm5tYnbbDLZTr6J/D9imCo72brnxjePfdIZMFHoqSzpWipR6I+155FjatcsXiPFK
G4c2HLqzWsqvQH/GawbhGe5mIlFjWML3Hv0zyrQFYFjKFteMVP/GJZugJwh23NyL
NaczBYRAmEaWUpxn0+bpL6RfidwsDzViDJ43X/MvdUgVTKJcaUxQvWEyHiFN7U+G
vIkauXRxQTqefr1cwQZtGaddUSz8oC86UjvrzrEPZE77emPrnssYvUd4AMqpbq0t
o+wwnJ27TBY6r9HhkfC4Gza2aCLJbpadnEKPmD+VLhjrK6nzQN61MFaU+Bs7cIDi
e2vXXTPaJMOV/GHFsK5w9fowzGMP2O5R0fGfLxytrCcy6V51EtxmSTM+kAAkZWhT
aoz7M+jzuIEJBbp3R/g+kTQYP/y+ZjRE5Og1o/F3aLE/F8b+4RY4MyFJxgJmuiEw
Lkjzc4qYgYWK/XAFqm6XEAlY1+CWemtLGa8+HkfakyPWxqMTSt5eFavVoI8N9rfv
WXZPJlxMLPNbEMO8s0u6iX/IW3M+cpSDkXSmUllW4VsKZMKErOUfm9pvvmn0vFiy
fBLvVPGdmCJx6pORtFwCk0XDuUfllsXvGTBgRFBKz3YYxo9yfge0RTb0ZKUwNeI5
Zz5FfTSAi/TAK9sHBA5KEwXOC/JWz/CNjTL/tn0p7ACNjTxVMmwtmVZO7e9UNdaN
Jr9O0OxoKyiqHqL42Gns6y0gHsGAsP0+lwuVTq5uhU0nFRo3L/QXoHgAxpnpCGFj
8ARQhv/zv1JDWcyIQ8cXG6ihjtwmkLjtNu7wAlITNkhdsPSnNkzcQa2Nb357Axxt
d3eAj3k5ZpSICxnRgl2OqWsPTd9sGaDXMormsXoJe5/5VegICD1q3RVpIXSmSixM
vzmu+USt+z6AhKhdJrmOTjBYX81FgNvxDlhzBHcDs03Txz9Dua7WvK9zI8+9AKVY
m5KA4KiBRGVCCGQku7icFpu8DmaKwI50LHziYXiJGHyulnvD8KgyftRVHNTX/S40
A8UqD8xyzfwugCcpPt6n0YYUfLmmmz0zBhlzQc0nQCFOv5UxtncLvpbr4nI0X6YZ
w/QwK5lNLcRlQxMfNkOEQaRxyoLfO14cKAkK+0jEydBQQFCJoHaFnkm2TYaRShx6
Cp21q/D6dwgMpZUY4TSGIQmCItA2DXtcH1fT8swv5/obRVYJWCqy2MkPqOWZnlQ6
Qfyzb0kvT9Ru+RRyBJN3MwKRxpkJvOol9luj0KrGzTKui2rrTSLQiQbZETyAVdZC
eoYqxqMHQStXaZ1O3y5yum10LgRf5J2Ao1re9n7K3XlmFpD8S2263TovwjPkAUDb
gQbWG4gasEcU+tGu5J5SdfM9zoVbAeVShMq7VVl6E45Wud1tQZmMcrdfJnIuKC0E
XdTPuIyqhcjiuex04mMre0XmGw2Patlnri3oOlgjS3OnGkOD5esalJ1Ta9yewYK0
VsehwLBuXM1OxG1ozNbPPyQo4oCHKBz98Y0kXCNvUsFsC/8n7zc+eId4SivXZ8jq
j4kjaG6bsoC90QF5jUWTff5/uQSfDCK4O/m9uWD+u/Bwva6bUaLF9SiNv+lxaqWa
8zfsbPimJtl+39vMWp22v+Gwc8gd1jVBo71zKggdj1tNCMUwzs87PodLQaPZAKw/
la0Il/aTz0uRjULLoiiTDC241+gVqKvfFUwyL8Hn9bkzPOQEsoTZmjsd2722kHnR
Fn4Bobz8QXPGp+j9j92L5E2IeblfIH1tHZS32aEbcfNAbklKZyCuzNfdRH2zinqP
sudJ3WGG9WVtbiF9vCc6TCxFdOZ0X8anCyebcLbiszA5k1K6UjDckQvVK0zdYTXY
Ini0Du2QlVIiDdRW1ASeka1C3YdgCd4jp09Z8tgh0IHBqCXr8G7ZmOw4AGdkn9yI
pMBRKDWTelQbc1PNhQO+04foAsLBMJ1gvoz8urpfNocXnfw9qCa8QlIQYuZeyXtU
lyA5i9DKVd5qecrMFmdmztVNuZWX72WzJ4ydRUQVP62rUh0oZ7F86Rc3V2zgIyka
Fn5MnOm/pQlBPjLCqHLNO+j0xxI4x1w90oYwXmEYI2wV5NOXzPC8eL76t+GRuBil
78w6apFGqtpI2oX5rfZFu6IzYRWnJa6HLSgxxplny2bYCfoXZ8bgTdwkxUjVrbV6
DdwFMEnY1rNFHyg4xohihro32aN+gr49axBzkFIQYBnsmZFzO9vJIy0lkQcHjwh/
11M79Gaz5uN5Y6Tyih+PB2Bug7NwsajtVwebHhscSq9cDDIzn18V5hrhmAxKzYrP
JoUq8F+yo4KTGMm1n9oDsWFm5vfgTc0yh38b3XZlTXUbJraKmKESiZSTdzr18bGs
IglTCyUKffky2sZoCU5B7ng6khNJwRi1umv0H9nqM1+kc8/7+CgmvMLz7g8YBmOe
GS8BHVS2bt8x+djlmrAjzl2Ex0nQeIDIIKk6J4FxnYDycOvCXyZ9lQHCOMaj3QNy
UCLDeTY1KKCFFjLdtt/HMB8RgSF3wmR68XPoF5upkDMcld0OBOGry+fcPjced0QL
z8TKi1rKIEydIl6xR6s2HoKHy1KLnfrElw1L6jBYt/W9Luc1Eue4cbnEt59KsIK0
XMRIJEqy/z2qFCuDXs06/lbMz6tsvAbflBvtK6xmCM+LW7/X64xPlAm7GSUGQMqq
OCMXaM4MZhqQ/WdtJgNonivhMX3Nf9FGc7T/F5QmCttxT8/8YRdy6JJaKtFTHN/4
2T6uvokq1KAKwot5LPBb/46sRvR2qboJ50TGewVTPu2KdU+rT2SyCpYbWDyIs32u
sMr8KYIhuYaq4bl0t9XIXuRtJzteSum0QNkkI3yv+rQDbp75y3VVl6oa0afwkVWL
vS7CyBYJYQKBnqMiXHm5MDW8whcjNUPA9hqJ2LlWe60yqQrYKAWHjDaWscAm76JP
KXG7pNs1QCMfhcig96xS7hlt+wmrQQrgqT9b1+q9vpkM2Eeblx/ozxtsBeGuuUqV
KogXdkhqOklHijTXcQLDZZ/YksvW4uWPuVqV6Q7K2OSUMC/hsxFUr/VC5VSSJVEr
NcZ50Ni5BaTpiTLZSsC8CnILnh683H54kmzVhMLC5ilTYK/pL1d9fQGLJc2KuNkZ
IvrF+p/t3FG/3/QM6bvpPMzk6zxcvIQR+CS8NpXYjTnmYiSVOVE+2ZTrfl34rGIv
qmGGKuCtYDq4fg51gNlsFDB4gHWEnDuV8hLqSyx9m6PHrd5vhHLiO0P8VEdK6dKV
D/r/jmWt7hCi1BJiCakmLhqhjw11GVLn8Yy53tMbaBbXZx07Jyu+KUW/QGMNdv9a
fIy8GiZwYE3T9LHfXkZAQXC5/5AN4FoAa1ioqIrwKcBQhQTh6CYD62XFyPryR3eS
j0T4nWVUuSSsAqHtVVrvsJGnzoXZHOxwhXAk5gKORK8rSqA+Xpc7b6fvRMBnODTc
49PXjfvVR03X6gtlbIzHOb/pb9UqjgbtaFKO1499xzyZ0Wg4SG6mL70z4NHQye1g
1i7SQYQ87GCaBjlLuX6DZstmwzMrIE7fdbCySzeBrjXbJUw58Ql8OnxbelM508Ts
4s9j07DBYQghEys3qUaiV6kL0Mip8m5VdTawcIM4QV5O9hzrk2tcYANp8YAUV2cS
Ibd/vYEZzyOlbBeIQWwRS7WvenLFVuEeUO7x+9tDfyKYgmSEHxanUfDdQ4CDxeFU
0OczkGvC34VGH45SXGu1wkLN/hoOqM+NceHawlk8ryCTbtG85Bx6hbLOcafhNnM6
C34kHI9KbI8ajzfP8oOxHBkqNyDfjwlF3huNi4jxQo9I6dPvqCSt02HFd3/cYUfD
3IvXmaCUQpkbSmQ3RXs/ZzFf75YMYRFM6rk/xEbmQC5qIMO+iFNn8CDh4tkyiehc
jaN859NG32VO4Lx8PrqdzIj4sLldPaVqPilmSZ23kg+srUA7eBtbA3ZPqLmA7Mv6
KtbVvoj1qTICB/Y8hVRlEfWPX879sDyao5bjOoA/Q9+acdRkMnCI57degDMPFc2o
a8ZjaVIJkbqJq1hJCiAQqtNjowYWMhHha7GHVFUgJByXcuWwJTZP9chX+7Y1OQvq
2Ra3ucLRW4+IoM2oxyZUkfwgv8EFRbbSKLtPzm03EhLrcQO01s79suSMyp6WMeJq
GwB+Qcmx7nWClo5bezZQepJQi4k1b2QqR7Md8OK9Kd+nyHdvK1bMF8fsRnsZ3dHj
5My1FHtrZRvkPedbO/veVPJR8W8GUqluJAOeZqLp4jAx0CxrEwHMrIDY4we0GKQ+
1w3U1xYZ7nT+s3VN1wpxAfaOPQWNa6Vo8XXvGMJnrAin0G6eWWe3LZ2KHAKE/gNP
klHXiSrOHUAWf2LcSZ2RFUc+C2tpXkurYxyzTD9zBNV9PbtX2Hw59wNokzfIsKWi
lAVFc/NjlNQAcGXh9/puAdvR5qcZu/f+UWTdV+lsb5Xd5Ezf2e/y9Q1OLZeRPDiU
L06b6WuND2Bqsga+YFDihQ4HD6AemKAkMHNJoDqZM9TRlZQvFrD7EhihgrQk1CcQ
jJNDRA9DjmkCCufZkF7T1ExyXTaI9uDhiGMXHxeUehH7kGlX7m9Y+T3Xt7Q00k5W
d7d9P70GnFkCFRL3Zbe32F4C/pmfDyCjok7coO834QyTM49t6EcQigPI8GZn6EHZ
pSw7M7aqNQgIxrkpl1lPY5InWnlnZ9rdo6u5HcVmP59KnFCmkcvfkn7g4xJ5KASR
sFJcet9/orH4trAUlnYCsymsLvk78UaJDFiaGlSEAYsFhAd2kngkCJdmxX/a7SJe
F+SBv1/gvW4nTG5ErK8EMrsOJPhdpvaAZBN/oALXyGgU6O7Jnxf2yknlMx/xS95U
lmaMjgJuN0uZ0vYmSHzGYrxFxXzzUparD/cStmAQfjuJ7hiB8iNJWC7fORnXGFqV
m9hZpX8GeuflyeG+SmNbxqYgxqdWXGUogZ4kGGJ3tPSKvth8UlQKui1Zt3Q2T1dd
ctsgXmUNXgfPHGS46HyZM+rNLA0pmyBs98gek7kQwRjR92v0j4lQFDgrg8om9xJF
c3QQmB2J6Oy4V0oJtmbMCPsTN+9n9tqVCtUqavFi88KLU5ob6BVNa+lRvgFqeCGJ
udtOTaiUy0rV+qX/dWq/kcck+7xaHOEAVxu3VK9OcT2feDqg9s0t5qrXJV8kJnkp
tVfpVDF4cwUfdPjSBgAJ2LfAKCDk3bX/C4T1ON8gETJgJHoloeBsiP0alWB1vbOw
ErPer71WuaKFG5fsaz3lMjNpAJg+098iCiulyIogm4x55tA9k99NXecx4jHJJUFT
277v00JXvGdvL33BEzDKVqNe0Z9e0l2V89q9aWFZaUSI85wWeecRP1cNSFYuHItH
etjmd3MZFgwH2bH2La7XFuPWwx59ZuUsogYbLlNEdVNjZPAktOcG8BDeBn8KyaSB
ytYmehK+GcdhqCl5I+wW8pSwgyFpg4DyUDoV5y43growX3ON7wOUMOujIQ1KykkE
7oe6jrUaE17+APWkcKzzpQH9rhGOHtCrazDFUOFgUlUu5gY1n2Cds7ucBC6EZAPi
B5AzC8HKCjw9AkqUErRnDSxAZF/CvrJTCRFRsMDIhJUzkQNo9PVubo9NvEyaTq5I
CrPVCaL155Mvd/3JSCh0V4arFibXxWOGMsxahqDfibKvCD84UZmy00mcpC3au/MN
e/JXnSbWQcBvIbJSF3Eeiio27bs9IWO99fJorgLYr0kwubon/XssTt8DfirQGyXY
qnHmhLxxGekp8OyXBBK9Qxz6ePkUEUynkHge4YeZQFYZMi1FgJCHyVfyme1riksv
zNxFLOumd3wG8w6rl315NmytxITostDhDyVwGaN2Etkfow5bbsq8x2lzFURgWzLN
vxTfT4GaF/tg5MyswQr3FIdR27vG6pjN78YQzwiIgwyAracMrPw8lw97SzITRI/q
+ZLe/F5U/qlbvj5niwDRv3rZkippecP5QQknLIB1uAzcgEAh8jglkpZM6m1VIIMD
Fp6CrN7rBZV6IygPlf744fMnIQtJoXsQCPA78aQ3M9pPWRJ87leEUpjTHxoxAkc3
DWpVgW8/aaM9YOo8wQohlqot3hiw1gCfh8HeZPLLzsUmONG9jG8jEOnRHLosBOyV
eA7VKaeIv0g5iiCdBg7VPcitt2IjTHjidXsucz+fuWwHvtnqHCZnlr059/0lxSzp
iu5wfRPfhweWanES+K3tqZ3y93bxq+Tyy62O1WgHeenfb+CudTfvarkNBHZfX3wX
R6ERDuZax5qT/8Hf4afObB4c0gJPm/qH4c0GkiObxnzbsMdYFZUCp/yfp37y71Kd
7IE6+0gGAacX3jwtY6RBsXsHj8joLz6AGQW1rUHwet31ysR54U6KSWdDXqvpkuP8
gNPMD6z145jAOyyXjTKbukkE3wvClUy5gos14RK9Qwl60pyaxjEKC4al8CTotQPZ
v62i5ViH+ZjWejoh0fVqaD0pguegCp4Vl2jaVmJwk1gdfYalwzgHMPcj+VnEemqZ
I6o0P5L6Hfpyf084mKvCn7v4JP2KhhEniEt4zIuvtCPD/a0ukb1RCtU4aozhj54R
CngTdJi3EBCAH0nO8Z9BXhIXRiL17L6wwhEZS5DMSfUroZdMY/fC2CqmHg0ZJuYY
7yrOtQICibm9LDgjbp/QTKrzxO3KSZ6gwBjSVRbLbj1juH9BPbU3rtkOqK7dze0K
tkKsmO55zqi6I0HBOZ1oCqXWjDKNX5QkCf2cOGwakAA3oi3+5HjOwBmCxUNWwH9N
c6GJQWPkb+TVIGlExOJ2CV0C9UaBiYGbFyJSOANa2uGv9C5g0VoSk8FAuaZDJ59r
rDQRsoaiKCEq08UhZFPQJwJaYC+p7xAWUFdwImIlkJFlHiMiFP+KrRlt7z6VG+qZ
267Gl/9TzEWPCKdgdci9WGrzB2uCkRy5UmpBAJVxjiFAVCuNMFsq5+X0vPbpIp4t
eeN0fLCETspXW3LqynVyjtwgSuoplZ1IJLqG3P0bXC9ll6syNBYLChDhpZWZeCev
iEOObqfkUFCCpmaryeLTwiTbR6d1nMR9n2tbDZnotVWoWeJSasEkTz8dvQml019F
ySUvtYcpaen4pbrfPEsgNlQF7HmhW1W33EhfvIkcQa+4/rJpYRhfUis6D3sYkz9d
TcpS5O/yKPkBZCoH9TV0ZgBlTGm5PLu5fkClFUdBcd6U98hjnbiXKJTO+Ud2ifXY
VqV3UmnHOFjJ//kaXi6niyM8QE62cAssSG+P9wQVKsHPphwKkSsVga15pBxdf8CO
p3JF9P6roMyP60+fXWm2icN4nxMH11g/LqzFi03T3NSGGq06tLBByGOmBQhNGF3Z
RBUw9zhJOkUGWt3aX0WhM6f/Jxi8E7h0UQ3n6b7p1M6r47gUJ3f2JxsjSXyxV/Ap
GHK4fZvkdsP3Q398zqItFeZ7zTYZRNIiux7mktZHcFM9KxMKrMCIJv5BoK+XIpF9
fq29QPSMuP/XOqqY3ac5qvQ6tmBjyenKq3LFn8dUlC4ShDBhHIosWmECMtsCs3GT
DdAr3Maj5qiK2k7icrJ7NFDu8cRtKC7Em1HXcbvr2iiMnCblzdRBwgFK5Fu1gmHp
VJIAGeg95TcJGlxlGx5o+EM/LwykTIadMTzysIvcsSZkLWtoLWl9qkSBlnIAmnu5
sRPxgB9+KvYZfQPKjxL63ejjaiis3zteSluw+AYS6nr3pKmcak8nwCh+SsbtozDG
UC9EGDMU874e4D6uSifhxuWt0pkv3ZNbG7vA8WIcjIFNlrQr/hE+/AavkmYY/pbB
dzrtgYqIwku2lZo22Go7TId1I7f/XM03lbNbLUbxV5uCbJTzSUsf9V1mnDfn6bk9
3Bm1iVpGYyRx8yLBg/2yhuNR7WzecqNJkd9f7Skx/TuEtbWdCtTSX+yn+DSpfUUG
3PiMPYZbWJawRNlLgIzj0+1Annqy2s9OUhlDe1bnGh4wHRli46VYq+YyHyfVjCff
p+DJgJeIQunTxDjsEiNTp+6cBzC3EXwBSUiiFYtGpzqmzbGsZTV6hHG3JSbR5Fqw
yUeSXufejQ32ADx/VJGQUxsVA035pavq6KejqoZyq3sFEt8l38NjIGGIEMUAbQWY
icyjTXJ5p1hOOd83HB6uUNOmm7dcHquYRVa/xfX8P7OMDlhNTAzTpVWuWasj1AoV
/C5YqeO03RCXwRp/tFkj8g7w3JM4RtHhBse4tla2FQU2jhZlBhywks/pSBEbBgzz
ddF+BKT1QHQcMXeC2axLqhEPWePCVamWFE7d1srRcsPZGc5tZIUMmUyiNTR9qoaY
x+I+GOgSscdsC09e2SaXBgZqIpQcYZJj++okdiAcgeEV3HeCECEe3HcJjRZ3oP3i
wty2eDg0dnWz0N2tQfUI7FsOEO8VJm3VacyZFNkX4ftaGNGt2joN/fx9tiop1i/J
URLi+XoUhyGis2oPDDDiaQA9f4Imwy0UtxfxDt+x1DBRwMDoTfOyU6w87O+QsmwQ
hldV+c9SlEc6wsuguHo5Io4b0DLE2vAaC76RqJ5hwRZLr4MX2xc7H2+ZmLhB/bUC
TSsJPPHYMr0PaQeet5HL4TaElLDxlgAof6hHLCbIP8cHrgOky8EiMG2/F4x8ZQmJ
t0WFTFHTGRUsNmCAEZ60/yHB7AT8W2NlGiVa9tp+FOoXSmC+xS4AWk7bpAYEqkvj
S4/sXCIh+ZdEwn3NcEuzhzRiEh+9Dk7gOZ9Nxy4l7BxlZM3VjkdmgOl6DVXsPWnv
rsVtxYGFWO0mq500byYSwwAgZ/iAm1lTYNAW9V1kRJ+snER+rTVU0oRtuC3YHly7
dIjsK8r7DX0rvC5VJA3h35UlE8ItTkUZj4lS/LigaqKd6KNahIxsklyIMacQcCQI
QDSygAny1OXsGK3xWdxud7SbelWVbE2plndfTUj8WN9EYNJVj3j6/lklWaDS77oO
CO3hscFH598u5pIhcUKYXsEFj+dPI1zoq2KTNVfiTGE8+qcWmhXCKlSJAOOLecbL
qXVLJTG/NUJ7i35inIMa5G4zXXQrSOlQbePv5pQFKkAUTYy/uRdRFqPCsNQP7bOu
J9AeaEo3vHjZeD1rc6/H2QzbsObsOXQbjGmsVbhOGQvn9sai07gkqdIkoT+fpfZb
RJCr/r6mRJb5pknh0H37HMo5iSa+a8qfWIRmCEk19tpmnlSTXjli4+7fSMiz1334
dO8emCIGgzgHtQdpmxFVNZmdqIyLXSDWF47Y161bdTFB0DzVpE4JDZyBUKpk6Qff
1pw1gjd0cNmIdHGCsc/IldOxKchW5HQGE6rCP682+4vBpBUCuhzQNoC8YkQrmrS2
G4uuLZjiSVNoBLU31fybkTQLiPWBR/iSk1Bp9E8wa6tcnM/FCYSGcTCpM0AKXq8O
BOh9NIbEg+aG7YhQhHat/P+J19O7GNu6HRLbsZ4SH90/R4SjIRE5OOSCHWNDvqJJ
PesZ6MskNSOn7wFHIKphsWSRUl5Te+5kQ580NfzFw5bgImCqt8f1Inl7POGfWeMH
wq+fPYQVm2q5w98mvYkX7b8gdAYYslETpYhcw349pRtCUcLHvRvXQZ5cSRqrwCwd
q/59bdiuMdCaZCq/YX/hxZb2T1Cj8DsO+ef/EevoN5baA9vBG0WW71GcJ2KGSmBv
z8N6FzL5faUBGuCdyNyc3eqYJF5biyrf25+4V4j+vwfqz4N6FKSlua4SmK8FiNmF
Yn3m41HSBT+K8Upr8IPNimDw/sFhSlUOH6IMqsrbo1mjnCivYJOWKCreV/U7v80d
BfJpweL8m18tGqycVPp+94n/T86E8lmJVX1784ULs1klmk2ff5SZn4v4PreDBRet
Bghco5nMhvGUs82Zvl5qf/+VsKayVkKJhciJkCrx8/rz1ldJSSi7MfQOt4HsdHBC
+ABS7nlZbJGQIRI0P5puNr73KHYVkFWF2dbw5tUiSHpnwkURiIu+9hqWWYataBM6
BZh87p9ePtjumXT7GAwfrmly0hT2AiOZQql6cd0WtLC5awjaGRoBnfyGCLN1Im5g
m+9+bcpLcy0TtF3QGR50AsHowF7sL2rLPFZ/wYEcgLWnLAUCLluXWm1+hy5AVCgs
+nQ5JqGL/ogpss5oGz3cqBA4g7xNDX9qhuchWhpw8rCQzUN6S+CBYePeEy5nqB54
OlPjp49Bj8PXLcfPzMirGJtriOYSJ8Jq8ZcJ4czxH4IGiMnh3Ov+BawaYlfRpxFy
5J6Y4imgO56r0qKfCa2xlQ0MTmzCvnpKXypYmg4goaUDuZTGPBRy0hR8ADda8e5E
irbVxC+ZiR9EQvy9w6iCFfTZVlsJw3OmXW5kJzaUdWz8KOdVzTTgOMp2nziWTWeX
Gv1rKXIeizNfJNj8nm7BnYub5fCua7w3QqpdViiGG8nsAectf+mRegnsoajSgvBj
SDkib7GGHHfcTQgqXRi/8PZZcnJfKEK1ZZv+9Q526mYJNzodvcJhY5Cpc2ue0qAW
htwYBQ40OUdhOIpdunNCC1MhJ1/qFI33mlTVr8no6Nagg22pOUhQR08vEeq9Zh4o
SHqlJmlYLsIzazB3r3O4RIGJxcH3pXKVQ997i8FMfmY2OB6LfIg++4hDD8fbAwHv
BznjTdtIK8NUI9qHUcfhSIkOMbg6NMdp98Kas9n1DSFSsIllbW42nDUR5AZ5vCZo
0VtOva96rYFVHgmVJZznWlWxsoKns/Q/Hzis5hSs8ghPhw8T11vZlBUzcfSRgfmg
6b7E5HC9P3CZ+MAyuqsMgjzAboXTMCaKysiVpENkecKeOF8Nile6hFGM4iknwh0m
5azKO4UMcPLG8GgU8B7y9XhkXg6bpBnqsYadYux+ZkM95BD+Y7gZEpTFWi24qPYS
lwo+IfxGBWZpJycVC5PCcl4O9mttAcdKmnm9g/ALmLdr/DNzWa9y1UKTVoafjce4
S/J4AxA+FeCVGgLE4sxkY5NFC5dsuqqi+Z0p867I6BHtRX/sfKsTR42JxZqiS/wY
U12MEbLVD0kvMGWypesiOnw7jR5fu9IaBS/YVV0JrmIEH8iMLFyLnhEROGq0OJSd
WCX1aRhWgMenFUNeMz96u3nauBDv/ba1RHI+Hn3jJumZW7pBW/71cHZVN2l0IU88
8rARyEzxvyREEVLQoCe6ke1Z81yxV2yz13FLFdAG/O/kKW63Hzcvm4RUNigvPjvH
LrwM0lUC+cFK4ASlbtEcg3me6+lB+IFRrBVvDCpTiyfwX6anvQ7c3F69qXbUQxmX
rjra6JK5EGqBfTz6CjJWzo1YSSzjKgX/pXcqx0qlLGLF91xz4fKTJn//EntLliez
cDtgORolWn6OjwE2liQ/HGZZEjpyRr9UAwmi8/uWNPa7dvJ6Kl2fPkUttfRbDFzW
RiDhm4fp+F4eXrjuqZ/n9gy+P3651QOHNq5lWRhXWltUVI8DPLHjp/7VP2TYw/1l
pbK8iM5GHNvxelT9R/Lkp3AFzDnY+eU4VPDNoogOIb1ZGaEEl3aERHVz25A/UWZ+
ggiQBRviINOwkY+OB05VFcVJ6MUOOQQv2g68ZID6jLDL1eO9H43NiVl64jdk27n3
6zeWX3pbyts/z2/UFr0qRnK4MXuKeUsl+s7lKUOVXh13gSJxRx+bV2W/3lQlp8Jt
UPWVuVxYuc0qG1EByXDs78P2NhCRvKlkF3VW49kfS+tbl8q7ZTWwMHjJ5dtEA6Np
tWZ1w9TqcY3Cx4vAErm66oc8aqhTIBXqpw9klQh6rADgyuM3qnBhoj9VkRkUDl99
tbCrUY3sBeLV4rhvLD5oAOBuZVOia/6WOhvRwbO1nyLXunBQsqXTcywGVUqRrzNI
7R7k5mPPVPR0XOplciB4Pf5C4OEMS7SDMhq9eeJQG2sdMvwsZq1uQKIxLaL8DmJZ
TfOqrlRHafvNtxHjhhgyuateFwz8Wv4jrJdOBBHIXWCHgmHThRWfnvHr35loUty/
lFmvkxjGEKbkUKrJOheDQBiJ6H+6H4JU/dunOcVhnzA87ckXM9qf0b5Y+B9gEuzo
C80h9EIfS/1Ul9yfP3TE5Kz5yrwbtp+RDV46o+ParvC3d5yvSZzBZ1vN2ASYPEYb
VL2kM4B0DDR8xPyzWRqRAdF1EXeHkv1H7UKfhke1jtsPca8tweAWrsH+6Up1v7m1
4Y8gPKzWpQhwRcXqpNtWQbDdrn2gNsdmcxrt4CnrLJ9hWELlU/kbJW6EAYgCjkZO
/Bby6GfrHarj6VLH81KTIq1R+Ml0JfXRwgWZ2VH9mQjZK5L07AXU+ffGLSYdNZ07
+aZSPig8m35x1mI5/4PbmarlA48+eGnLUc6YULXPmCLQSJekAos+7QCBHzRwbUsb
sCxwZdq7gcgzt3iM8FJfYW7Vf4dZi9Oe5CNJkeJ9GazFAZWMxhnU89R6j2+DIDmp
F678nvLt7RJ6HKC1TIPK8r8Wkr9WGnWEi8iPCzCbHXoVJkpbQXU8BKDOTbvMKOTk
D7c2XwKMnfWiAFVHRs7FWe1oJb/l3a+7PQYTXPDJ2uElDFs2y9hUoJcBuQpeteL4
/t8bYzF+0I4kJ5Z/Ft7xk+5CoCcE7mRHbL9ONKUdXhS4qSyY7dBdhLNgUbwCJIX+
1hO3d0zbIDYqNHCcT8yQvRruYbNl0Sfwxpo50HxPA+p+yqQ308lmnsKO7xLThQrG
ywUyBVvjHWY7fZQjxHXk0PYJkvlBdBtixZOjhtb1rZS9k8IbNhbudQrP+lDEQUC6
LcIGqD8uowimlnyKJzplZs2pqzsty6g81wWeAeEgjootMkeUvJL638moUR7sVUSk
M9VS/0D50sLGqot5ESNddApmBTKTyiMvGI/bdnxY4JM627gRziSIvGjRMiee+/ov
JjxzqKMgwHSAJEw5Hi03XnIqmcxK4jCaAM6wOTLmAuLQ4qeE9jkLHNDpf2kbXPFV
8U41KXTLyw4ffZyw+CqKZa/1wzC3KkLnVH53ZxGgsiMHs8mfuB/7k39dPDzqMaYH
oz4tK2WVsEoaRXpQZKDWSvEooXVZCXMUwmdRHgl7Qddhic06hbK3+LXaGN6b3UXg
fd63QEVz/4B0DOaPCyEIs2mieZro/9pjdtX6Q/ccs+tpEFVirIl6v1uixl3jt9ok
JW1BLgH0lrGCKgpYOP0EeCycPDWMNBp0U43QfwIqJxx4HLbN7pXlGyhxPsDnTyGA
4W9rhng0GUzBTE/CY2LY7rL/tXh0r48g5XSGyMp8DPNIdgnq2zb02RHFQjij/Gkx
sAjLoI9iVGlxTwM4LO26CA8Nc+krxd+V5IoUJv73AeE355EODGs81QD0k+cjXPhb
rOAooxtlLR/uJijlG8cOH3heZihxPKe7TwsO+lRVCVEdRYsJnx0JWBcgdv/M/ojE
2KneLbPXOOSmiikoq/oaaoPn35wzUxYazTDc3In9L89IVBZxnfCsZ++B7b7nZg+r
v2+f0qRN4P9QyOdU6gVbLcXyNs58PgJGx7QZGoUZP6RtQR3sIdbfBFVUt92/TK0J
FhFfUxhVIbmpZXrJE7dYyfLjnLF+1eDDdGDYQdsIvksZ0LFpp2/g6mVxl6UGk+EU
COfUKtWy7KNTfkO+HbLNbz03zSLDgzfvtyvBjLaOTYylhj4JhRX/6fQrW/7W6ihs
cAZH8mNzoX7AGXeUvEAEekWHReQQLRmNNLHFkBRUJhDCc8TqscH4pWa/ex1H5xjW
EHQB6Dm9ro2FTmii4LTn0qoxiysW+xt3zCESW6hAFTZeyHUyN7aVYyOnfxpc1sLV
mYQLSijGl79uzBo9KXu92/7SNcyXoNy1Bh+oNCSmfx1trWBv5/kwTyT+cMn++V3B
IhZC7kqry7LdHd2Fs6fyeKBIaAOWGfmYS3fTGJLYHXZoVTDQ/MwVSdtUTWmx78kq
2NH7xuifVZ1RHGauQZBS4o5RP+/0btxgcQsgZe070tGDj5ZmFsDOIXBBdQI9N5w4
F1osmmuApus0U+49kchOyqBmeP9nncluyf7v4zKGAep7RmjKJjB7KAa4H7XWHE9E
6+mERA2e4XV71yyrTKG0L7IleCAPPjmOlp7v+NtF3hRpnxxOAXxjCkQqG4uEcu87
ELNczbbtHW1eWmsNd8aLkcul4Ct7o72sNpZzwweCzFt7ZPvAkYGuYO11DqIblHTe
mjC2cJlS7ZhluBnMB2ItKBdDQiwsYOMXBItrzrW7LJgrb42pf2BQI20ZXzh98Fn5
gntYPoZcgcEfzhcNQduRX4trI7VckPWSiSk5I8czCtHhJ8Zzyfs5jnGhM5t2yHDV
ERiXrrvlRBaQT8//oLURK9vSw5ed0Rt7CxYhv7+pZlpDtfYace9D6AY0DrEWVDb9
vTkJFlsi1ukmYEmv1upX7UpNwz9/CZawpM1JSRFTZsGO2dnXnN88+MzwihQmtmN9
HNIqgFJsR4pYi2MfAdtojVHG4n23Yy/UCje3oZVAGEMJyaUDR+XD6lS3PiPuld//
FqyCUa+qlR9n7ELynfsjHhg6SfReU/Uy3HFSWnHyLwxKSKwA0n9INWjf8Uog2VTg
jPdWAV1dL2+SRi+mDkxSi61f5JHbVUyhtuxMcVleQwybB5Yl6blxmDYxl4Ur9sMe
5XuQFMOVytbxHiGfcjJUfb3bcnvHFh4ItAFx7TViwY3nfH2Ud1gPdBRBhHAdiU4I
kK94dOS/rFswV2g4mEyx0CJ/bst9TX7eJJhcBsS7u/M3Qq9bw8aPGew24bj/Vs3/
rrEDRMVANqdebkJugojAwlab1fYpjQe/BedyW0w9as8qM1i+Bm9BnJtsYKrkaAzX
vzMFvZP6tqS0fsjq+AEuDZGu1h5gz+0Czh1Na2zj7QjFHpmCgQPVt79dP6oDoer2
83/+DRtorP9A4xX/NBQgrFSfq4ajQ5iTpgDHHXINwc1X77D318vJr8b3jX8V21ow
YfvHqCwP9Ax1/tz7xWamS3clR2/wnUvDxS31nmrIst03H86P5LIwocBisytQmgrb
UCBNyOcp7qT/M8oLvDXrBJWvJdcUowhhwciuhAbbWCZ6c2EcSxUBjudd5Vqh+BbV
C7D9dEEWLhTUe3pAV7bJY4J1jntY/7p8TVUdCUhGS9DSFCz3JfYczYdQ7yQePYD6
f0N9Be/qQFBJwEP4MmzaaYVc5T2VIjCBye9cHrBjm+zR4WpMqa5IQYjodO1YQOgT
K29pU4m0blqGPopHUcjunI4DX3cajtSRLdATicjECac7YBpo9AI+k6OHS7pUj6Km
1ClPqB/nxgpmwmRLL3JK50HXa9UuQqBwjUgBt8DZzd1XspQhkcNX0RmQ4i2Q7Mo5
J78c+f4zM9V324Xmpmfq3gwW7v3arBK3OjNyDP+DKgN/xgOvx+8v2iLR+jIkFs0o
xB5Hr6Hex7HrHClzUO5801NJ8jtAwWOyr9OFfRuKj/D8hed02hxQEQHay955B1mj
c1ykvkEKT2XJRTTcAHCSChQalBKVPoa1sZWH+Ae23QNhaGLKCOcuQPkhGE+VBeN9
ZM/llc88wYmK5Vt8iGjBXhK5kqVZluOgXFD+MFeSS5MiAkNPjDfqYs+cBI9aaTLM
yWhAUGBtJAcmVVb9Q2nD9VwXHIoyCrvFABIIVskElWxCHhVqXgib+PVH3+V9ZFub
bmN+FFIMVaGWaryIdyB9CCLfnX9Zg2urcjg8kCWov+wbvOV4M9gCPZAGXmwuCghg
8rxQ5xYXa+B9IjPjzjVdBSkZ97p/C/e7vMgkzEToQDVHhgflV20PBV2K2sjeQuBM
r24w5L/sN+E43g3S1XOPLnHw5Lh56Ty1aMjMvA8qkjx1ya80AXPCCjioZBe1AdB0
Q5gIY+ssySI3Xtt1YjqXMNSTWYSvdqnOGnCsV13nUQZ+W+upGiEFHs8NlgRiQBbp
vToFwh9gA5rPGSWU8yHVL2BGyRpIULI5f8J52RB2mJrKTwreHLvmGI+Iq/mw1ilw
K7pAK0PBowlbKhSxDYjm9cnHR9JIls9KxJzolJRQ7ckC5fIs4RREbp/eJZ799g4X
rzodKmKsLtDDs90JqFNVtUj+5Eo2Fj08a4QlTaLaSx6PWWDubgW6LrJBbYvZt+B9
LOx7mgY2gZJhuva3TPQK94+ZtKRyvF1qmMQAyZQ64m/CHJgK131IpicAF5Bw+Un6
+L3J6keKfMQ6Q6vhUTAzDuwcKVH0zOwJ/vTvFu8YyB5ZXmAyzMy3IvXS2HlkLoKy
L+Ir/vuB7WRb06/QYU/JFdAa3inhJBQtxMj0CNK8yHsxYmC5wm/1JFPifxAFDJf5
t3oud2Cgf/Km0wua1sRYrnVdcMQEQSihBlUPtcyKZouX4VyjBKrtUd8xUj7mb0Nr
LhLlu22s7oWMwyAv+YE6Aub2fWRIxvfCLL52lRdwKHRhB+oFw3cLqISnwqhcE44+
rxSpJlxvj0Nt62LlW+CLOfTvoJs8pFgKfBL7JHcLZK6+pbovpTKqg1uGQXX8cvVr
0bwXF3krZtqqP0Pqft5m49rqmtLkH9S+0ngHaCR6KSrUuFH+E3Dsg1J+gF9m5RVO
oYuk1CY0XyvSFSF8O/f2+eNSwh8bhYKoGNInNGnuPH2h0ZkBSPSJj9mztQkqumyN
QjyYqwjvW9ch4v8YPKwo4knzcxSM87WN3FvkGlcwyTGYMrGTcr0uVmvm05NqkEJ7
OQEIB+hz5PozWqJAGpLilsAUnI0X7CvUmbfdQvTITjeEuaxdYnyNfJ5OrshVdedj
ZGSgZMu1KYKqefAjDMYtS5xpiugJBQeq4KIGpgefvZyRs2xbz+bvn4NIcPswvDqd
6hbrhCD/IzvT0s9eSv7EzDolhyqrMbnHgjOmwN98u8Y5mvHveEBaW8RNsFoflK0D
lR8Zy10kyduN00Qfoi67z3Dnt0R2xuDjnk9nzfQuFMugIkS6FM60jNBN+5sNx02/
dew+jLpZm4vUhBcMLHSM9oePP89nmJC7od7zxHLYjXwVWN6wL9SOpAAdrwxzQDYF
ZpxbwR4lKiowH0FjOV3Oi/GyZfydSw7pB30On9rJocZ3SlpDKubuOCvvu1GsdKcy
Od+XKReVvFDGaQMkGGb33KrUbJ12aDIuUfQM06f9sd+5JzjaJuAq5ujYIDsinBqL
K14GQF61rtzTNSwA4RYktVR5iltc2Uf0kftGY5rpO7dNfual65fysmhOq1L3o9Mq
HM+5qWeBmtdrINnw653Qz4lwI8p+4knfJUMM/Ow2BPhatW1byln7zJ84R2o2BthR
rUJKRlmlmqnukr3dCLF7o/XND9ZwqmJiuprqOvNrl0QETjjnBtFvQqQCAgo8EEAU
WzSr9XSAYKDn4vsbE/UaGJVl62hLBn4UcosGROu4rN+IulqxtOiGPS2rvjm2x6x2
NpWdFRLj+U8swmBVikcOjF9LVoISifj0NY50tkv6zdxhsBNclPmkBufegnR+dVSa
lHECOawu4M1CAIPGhwlfveZKzBYuPw1SgRX7N+xhy6zwlaG9UX1mw01lmJVFzBoo
dSxZiXz+tGd0MZG1LlWJzQr3La+lOLdbEHvmUuNaGXzKh0qlr/xrox5lkvzmOU+j
9EcDPFDfas5ee6PG0M7148Updpe26PxjFpkqDZET8dVJgORLnhClEqFdaggMVAFA
+zrb3dx9CxdWQAUNBOM4NZfTL3QAg1aE2QSIzml6yQSj6k6arPfQF6sYE9r3/3UZ
vQezmQtq2HuY4wdF7uRjLO6OdkJdBJgLwb3JQSOfXSIBF3vRJxeiYlaaNCsWLWeR
qcuXnpMSwVYBV8zFD8W1iGV9tg0LACeek6ucS4/4NS1oNYebQOgLZqSQWgHdImEz
6YFZqEmBqQYKiDsU4+PjVupqpQcwdPkVZh8gFxe7fjqt0UXl6W8pdKRkRID4CyK7
k0rZSHpZTOmk2r8ru1wYmIIL7RrGb4JnlH80flnl4XVH27zjs5WLNl1mLwjzFpIo
e1KJp2mwlfgjwgIqjlu66YrNFFDdheDAxpk0vuFMCIdOc16eejgSsENX/kZ2Rapz
rMLOUv+cBO/fwb3SQ1KNweCQTSh5tUg8TUwDUSQihd7z1LyfgtkICh+yF5rLUDPs
uVI19Il6ErOs+U+2xu/wmY8Gg+7uEZ8SseM1r98FCMCn/8d3qhnHfz9sRUP0btPl
5Qb4JczhV69DYfiKpRYwl+6Azq+15T88U/48BcJb8ZdV9ulR+7Q2QLmlEN0Dej5p
WCU8D5A5t+jlaBvkJkfwZFKiWTJHQ6Q3Dl0O3wrGOfNkRsEB5ra8kYJMeuBNJMYj
u5jbXNCr5xwaxAyPC6DwgZQxSEhUsYKWJDtW9U0sklurOQWvnj5bxKY2U/o0x+iA
GiBGUAq7b50G+YvX5t/hTkgVJFyOxv2ArbxQ0tMwn/MZ78zLXdDCkTgFMAaTTI5o
2DSsSN6l3Ybpaajb/fcxTlXRCBqehObknfwRk8YkJnhbCFaGAYANaUR/rct0sJPt
UpRL2CvllD9dx5DtViYrt3uradTJi6d+0r8OXt3vA9STLWBPYJKXudtP/4wTWNNx
YGltSvWvvgYuw4luM6+eTEXKa24XruO63fYsWLHweurIvfXqcNGNaLQ2uF+hJ3Xl
QrBuM2AfZvh9K7SLvpzNgp0CnryRjxA50GqmnkRBKyTMtI8Nfg2Q4ETUK29mkjx7
U/sxfDoRbqchbsNrRIs/DEdNrRhhK4cUmHPiUiXKk9kD1gIjFcXNnuCHMYkzrYsi
6dzurzT2xOB8rxuZ2GuQ3kh9zf8db0e6b6Tl2dN7sIM1qS6XWZEdmD5FHDTzFoOR
/QxNEgO/icIx0HiEsi2S1qJYww9wA2i5EY9sK2go0G8RexXXu8KwO9GCo1535LVk
21RhUyQLkx8RUdKT4EHkEszI5SP9X6/fs18xPIucdBXjwhEHeRjB5TNTG7q9y43/
WFlbnSj2ecrls+9/CYoOh9/O+LXfv0p4uEHdLiszJZShKU8zT5Gre0iq1fRmsxGb
mDpil2LUZhLMcHxGz8U7MAq6yJb9XBxvojFXyolZL0wf70LvR93cX4XtsrmcuTeL
7oZKBd5DvOD11cgKjXBHLEnMgSOUhKIAtWOpEjF4QLInaM0e338+WZ5iN8QWfiNS
V3f/bzJH2Nhz28X+HNtqmrFr60sd7a6AzQa39oMMATjGUOugQpyOnSIi1URtWI6V
xttvrwNBFvGGd4GPblgkMP/npwl+dfhq7SpO+NNplTIUD3FxT/YNHQDlRn8A2RtQ
1MjTKRhqNOiDuGb4iDZQA3kffTAfO2vik0jSPgxC6JrGgoHKUqDy2ztZAuLcwu0z
Z5FgTBJFQNHqYDaQ7lmGq9TN6/ZRevWjhKdgtJwze0jEd7bZd/fFm8vegXr46n0R
UpjdeMvNGLfgbAjJPfme71VnKw/6erxeS5T8SN+Ux8xk0V2Z6KslYC4Bn1GuDH7j
r0ZEP1cemWC+284z3PxeUvHEZ+zxWOuO7meD4C+7pLk95Y+UsDtxuhPOvHxwa89G
9EzXCA5GqnlZJItYeajLVF0yJEedNZcPAu4rRpJVANEV18aiUDgAIkG63u9VE1NX
uX7Mdsp96jBxadRRhUNw4K7TEic+OfzU+6CR1CXV52GogRHQ3ztn3ULmphft71j/
kRZvsriZtdF58cq3KegFD6NVHSiYEYRK65AoZOpZ3SvClMbh58WQUD1KptNOO+nj
wFndm3c7P5NybcWEHdSzpqGJfHQjC0h/2wm1YWFof+OTg40/9TgVlhRprt50Qibu
0BdpkdWVYKB39pNBIYl18YIhMfGrLyyemvN4zMSLFqvpWUiTwYgRMfJmWI+9jB3l
KpetLMAbYwPDjurEWOp3xyYgTuSllNHk/Cznm9d2mB9c9hIBWYutsoOdHoynFJg8
Y848m0S78owrIeepPJayuoAV4eoJ9pg+GRx/BAfqC03YIt/w+VpXvYNJGDrgo9FW
k0Ym+NwXPLo834S6RH56II4UGJsiNuT9kXetqtda88fAZuv3myqeLpYC6GZxllbR
5kMVq8SwS2aqmFInEtYsoEVbJFdjq1tnxZ1BAUziciETTBUjMVDVSOc0Z91+AwjN
uvkJQB348qpOhobAIjxE9ok/NR5DDN+mHUVY401kAAz7aN9BNq8h0XLJT0lXVkEX
RPo0Ruq66dcBMjcMM9b4T35cv4yfZLRo8nAu4WGEv6Ll5ULznJX+Sk+sdQ0MMIy2
iNaA7o3Q7ECEy1KqTPXpV1MDADuLw40/6GcOjKQh3XUkGd+UN16GWUcIBzlk2GR5
r17C+MTvDJtTnBmSaOwTsJ6P6JBFkRRIlnRIytpfmaRuN9WilkO/dMdy5kAsrjdu
oQ8h3s0S43eu5tFAo3naLQkwd2wyv0k+Ll3SrYolHMMGjRT+xanlRx5tkCwtrScM
1INKI1f4xQ/4wnSNS/gmCj+wcVQygsDqPp+gogS6Lgg/6i2+218cYr3xt0yTpawr
mmO8Ad0ZiDqQPKAv0asiJE/Iw9mNjiD6DDBZbH9t4v8Q1ozEEPPJhpGd1inBlVQs
UWHEnksIiZaOKYdilebcOr5maSLpiC2Tq+8YRQsd1SIgmlsxwiZXguJaQM0TIcgn
Fr3o9ftpTgHrcyXyk1w3HeH8Wl5TlCpJLdSK/AF0u4/Wvt1ePkRQxb9WtwRZaeTl
+A7Vs7qjtgsgqdyKAuUC4SEOThI8X7b0P3myIcd5sv2Y39IydVAOuNFB5tahjIu7
o5bJl+GzKnNi5l1ytLCGr60HFPhlxbDv9Pg6X0VmrEs//vFr9ouVPqisweFYAODB
kpYOlzI8zAgrppdkzXJ+Ws6TG6qU47EWrlNcPPK3vb+9l2V5CUSRRGgFWh3gEHvu
WbuSNqoEK1FwKfvd+aTptmUjhQweIfHTDZbUxj3cafQ7v7+yunvOgjN22memUU1D
gCW50EDidhgs5KPeozxy41HVAykylWHkNC8hei4q7e2F+WEL6PaUCNbM0mVAaruO
dGC5upUbrylJVwFTwcoNYDr8lwMnkyLgMwmmYkpUxFJIwDmp9Flp5Tiv4+fL1qLP
P3xve0EzstSjVaEa3v6KITNjfr4tz9Y2v0KfHXLyoPLs/oG+yac2yz2BJjTW0ShN
bCMbWqLCVBuRXf190XlHJmJ3SzN3O2+xV37jXaeLkeJRttKGshWE6UrlajxJ5wHv
V5OwCXR237A+grMiL5oYifHOny2+pdkTwPNNnqWo/hu08t1Lngqcn9/zt8lcWMor
mtosaY5YaYiun+wnFns3KPHk8+36wy5oT+SAG8kbG/VIvN2UY5zw3f5JHZEnVzgR
K7xJGpaoAYyArHjLxw63+VFJJopX7NsYYx1kB2FIut1OnZ0xiHakZxXaUzvl9yeH
iYhKpmcqCq+M8sFZwEqGa5S2/OMZ119ITVSTdi+X9IBTcdyqz2kN+7ThDDujzfAn
xbboMfWNCcWI+rIiu5Hqc1LSioRDoirRWlO9OtQVKDnLF+4lY/waVVReNkq3IHZO
FXZNtFnIdeeu90EJatbGaYzKiFVtvCcU+RTueptZF9cDu9wQExIwIwrgreKwlcwo
MokxH9EqUwJZpEWl/kUhjkJdEPVvFeO9eTlW+T2nMbYbU3JeFz2+T2ORlyNiGM2N
p5mU0iezAs/vwWlHHnDbvGGSALsqATmvUsKmzp2jUvxx/5rp2d+7ZMs+aSjjeQH/
NjXSmzgfdD/GHYm9/8mdvpLswnBS8dEAjy2oBl6Yx9/jIa0yoIVTNieswITWof2E
SSVXdKMPiIuslyyq75I6gEBpLx9XWGthpy5fHUzXtCijn5m6EWJXMfZ3iALQq0RS
HVwM1eMxqIhvWwrz4b+19+IUbioj+J60Z6wxoiZJSSaT9bo/pUQVbaipV+fRCYQ8
hf4NRUs6TTo14TSpszTRg3SxVFhUERJA93tnUt3cm/xwaocQxxvZchgLwuiocQQj
cJoOOPlfODifJ1ulbleax58Vmn6FhSpbmasFnZYozpCqiKa7MphMGWsZ7DIF4Jeo
YH+MzoyINeGoD38PvKqHCAwPesIEiHyNpTX5jrygUV0dgABFvOFxEtLogElEt268
ZdPcNvnlN3RNDJ3XWdNPNd16VsC6J/56V63LALuksmT2S3cPMrqKwem4lmoo1s5g
ilkx1cEVbp0GdiR8cmwWnOiD1H5Dz8fSHJE9pAFi84GzSJjCMl16BSGWkHcBfEgC
Ds2K/e94lbPmY2ajpaVY1BW7BqdrpV2uNrsLZTBLaOPd5kAlXXDqWP38++vmdAxF
jqolNJZkjV3yMwUbdVOU0TplBPz5uhO/BlM0Orvj16+Kv67uah2fl5GQNoGtHcjy
2ryl4xBTAhJlmCjQvz2SvuG5VDchnDlFjEUohG9UQUPNRJlb4FFROW96bhjQVsTa
CkOSTpSnotpax6w7m7ktdPEoTp4M+gWpcLMOelZ7Jghn+prQaRkgbvlCKKL7NjKy
uXBs0F4/YugiYgwGqb1gETGJm1wbt5Iqg/Co9Rrzn7voNotkvj/7IgpagGtKzIjm
farHslTTyMhl7A7+IG9G139UX4s3h1LFyJsBUKDax+l74pCKwuGVNkX+HMJoNxqi
mg7ssoJN2arRUvxixcEwXDCJx/4Lz5AtrctV+nnHtm/zkt+JOtOztzmSCH+9Nu+g
RvkDa9IQmex3Vu544jc8s4R7/MHGIrjF7cuna5aro8+QHYuM/T5ctRM4p6vJj5VL
aG9R7LP0bF59Jtj1CwffD9ZxmPbp/0iO8osM40DH3weyoRPKZalTV8AYxvJCDTuT
fIQIHsRVETRKGGGULe2OnES3GSSFcZCVeVDWlrAyPgp/xz4pKeQzHDKYj+MeLXci
CzmITe9j9lE/9sspsZFsSsWb04XZpGrR0JCjY8IiIfMHqDtBMdih2m5yBEuVcy+j
NBrMXcBu1eaD5jF/FjzAPSJukQ/iFwxhpRl6dN3IwY9Tkb/qYkgYCr77nhUBaTyN
2njhlHnpjTQV6Ov4/DVJXAqsKhwgTPvSgCfqJ9yB37oXUdjzEM3AJKG4siai0+Ft
oRo3aOtzAX0mqOJse3eoAv93cxFF4EAiQ6lw56Ra/Jx7AKf+j0JbolfgCHb26vUh
iCJaF9NlGuIdxCzqv/Hy77ic7Tvx5B7s9aI+prByNivMtmTBEt3ZHkE1dnd9gaoH
dsxvF60lfWLzmcU2d+M/MdyZbPUMoBrjSXBx3m2yl4xodCKuzw6x2jR3T0UbG1+h
N+rYDRqQU9T0zYHjMuly9UnisrVnNcoMeRWZzJoqYbwl5Gk2p74CGv232bwp5rRM
6u6EqNrx64swR5Ti7unY9x9IvmMmWT6NVxQ/t17DZ9sqG+zxMrqTRT4HzDJkMz6x
EpEeF4/WwyZnB6+Yy+x5dF1FkwLQ1k2/w0lmPbT10z6suzKBNIj7fCe7QIN9YfY4
5d8A+qhXytePDTViJlFng5Bzw4y7FMZVhS5iz+lhcH1q2j3GQNNxXOL8xoTn/gAS
mZkgAWEfYmzqnIpa5pgf8TZriJQZNjbAt9Z/N1clGWMDzEbgVgzUDghQSsMl7uUs
IHlKV3HkV+YSEjQi/bdEXGk0xQinmUDi/QCdFcudLeqmFKhfZg3Jngj2Fc/E1Rc3
XqooKftr4ooP/OKzUpON2Cq7V6J05CP1liCGtsRjYsvEdiHrt0IONlmJULBe3R3m
sIFnkM9BRsxINoCi5tQUyK9NRbviYiCa6e4T2reUo5bJf//0GzH9RCf0gD5Bqvpf
h/Q+g2RfP96BWYIxgAOtKOy8x4Uj3ajY+/h3bB75MdEzFwxwvlS7snm7/Wd4nOHg
88mlas51AB1rT1CEkrMLaHgf9d/o7OihfsMtVySG5mAulKkJltyVSoTiFd5fcrAi
oHI3RXGNLsBUiFO3K8kzPUCGFWOImwBclPKam5VoapYCqRHveRJ4NC/rybfNk4Pb
NJs7RKBwwOVGz9caLRbChlNuAii04c7nwhe8bjIW9GDEDCTQPocypvMNRjB27jug
VEQbaw0YHodd3rOrxFwnDNBz53H/HcAJyXTgveSbojxa3H2AwckNwd1gkXYiC8sb
W71I52P8ZjgcmYvfpcsnui7FclYUHfW1hmavck8wfxIx03w8RjwQNg0YkDKRc7vn
G/TtzxInBA3/JCW7Pz25RB/vhgJQ5xueuJmebNkdrIf0qMWWqJszv1smyyfF5xeo
hLnocd8qlKkyFrQUTLj+VP/ubxQ+y/Y8RoubrvZwSdRhs3SbWdHw2VgL4+S7bjLj
hEM5CHOZZFSWl/VcVc7UkOzQVswySeRUEbH/xK/9/xrDyGntOt8HhHDwLph0qpWI
NtzVoadKI1nTP52sq6cBh+dKidL7VGSzg3xPNmwow0ymqxvOBq22z0D2XxwoLT3/
QL90TepPz2ISPQtLOnKgaoC0dwjrX/LZUgRWGCjna8+tokjkYOhuxy4KHVOTxbDw
YFQqXTUpY4ByuaT+MrUAm/B/ooy4Owtv/9ETcmfJKrohR1K43abvh9Mvjw2bQMxA
PR+RiX7iJTLmqaKhtlAn/OUins9z1ScxWHvm/6IHUFq1UF7CZyGLMr+w8urwu07T
sVe8HviFicR/sm6WZ0TbZ2aEKAhbT230uSNNnzaw3bWhDGnRF7RFqD9zmSShtDs2
kMh1+JM8VxBJ0T6cke2nfDR/6Z627298IPPH3TrQmN6w7dhYzlUfrOwaMQiNM1Tm
Hnz75/1nBbnXYLkxt6nqbkl4HbjfM+jJZiwQ/53tmotFfIF6Py9uYknziVLZl4u9
gEYv9Ov51Velx7WSM/eC2kJ936ZJi+BGYJ78WRV1gWNxaRrKMniAfQvjp+P7tYWb
ZoDEXJ/RxYbeLhlTSu7uhTdPBdumJuOMfRcljeoetC8md9b0KfU8tb3kb9AUsVzN
Jm1/RPv6V7LX8S3lFSuFNL4RBDblzaXBrtzQ/IizTRjDgn8oF5Nft1+yFRuVd7tO
Bafj3sgBXDEmIEWrmlCFJ575MT5ba2edOsYk2bu6SxZQl2mdP6PKZcv8cLy+U9wh
nb1VNF0EA7yDYBQmyYNHLDgOpwoRvtTwYCCwDtlsV7mN8gOGAvzwTeScFy52sl+a
JrOES2UCQA1wjZdX+grN8g1BYsS2OBs3rMXei3jgBgjYZ759IwDjo0gXTDtCWUJC
+hblgNvwqHvVbJQCRWlVH3dY6RGlx5zSvg6mXr9h0pudYswYm188Ema4sU8e4FGd
6TyQVVqpXi5QD/LoGwCITqSgYApZoNc9TDdRYw+wU0cpEURoP0V6IZOT99s8DF1U
gS+r+S7/Fc6v9OpB0HKOVYrC+O/DHnVDc9PBIe6fhlXdDLS7UyGS1KCverDypuRX
qlncgu8hI39zn/GwT7C/X29LcA+SWIizEwW9YnZqL5+vGxqljNPhnNU4aolUDaq6
rLzD3GQPg1WwD0C1X9ONMnK0zIsJk8Ocl012viFNtrXNaxAQYnP+gLpA3M8PAo3G
rzMmbLmOXJSqsX3t8scDXJLgBjG6i38VNCgB2XaGgER0lbPhiew5oaq5S1r0y8bD
AQrkCnBkaCmfcLJ+d1nz5Dz+z0lHHi0cmNq+8r0g8Rtj3KL8IQH53XlD+C1nJw33
EycupFA+LJY2KesCLW+ZOV3DsOseUrO7069yrxgeDCK6mdRJtLkL4Vk5n39jfXNv
1P/jJ7e4LKi7FLzu906BPVLZDWun2Ey1OyEW0cxBC56ODo4/KQXMjoC9SE5VwEj/
waBz74hYopToneugUgsDTfmfpRC6UgpHePus0Srs5Sd3bvlQYshHV6vcu2j7UvkG
GYsG+zFgzv061HVe0rE5/hXj4IXDlQUynRxjGKBOJeI7lT2zf8QSajXK9J5lRLtv
qGmYd9MSoerxgysQU8tpHS8XJnodjhRavGbKXB9ab5Pg+pA8dy8gcUORJ7WNZUWW
mc2GZuW+5WLaaYJqbuMZ66MBvl+OlNiauMJIhJXKdw2UWqi2IajIrkriZdUgdP5E
Uh6KEbmHyaLqf4s9HCeA2MPmL7zlkJU2oteCtgoEgqZ4iYJsPN3W9onjJ/1U025L
W7NbYF3xBkWYk5T9yN6q/EeN9oTLk0V2tBlAXq7rVguVQpZrmV9qLzPCwgvsoa1z
P/J1zvnQHw/4nk3/0xG8HQ3s6rKPwrcUkX5MkYPSsOGDwHPBh8A9G+ju0P6phNUs
dNXWikeNrxk7hcqOeStQ8qpLrZSiY82lbsZY/XgC3vcNgFLEXI/fQe8OF6ZfiacM
PKi74zTq79kVHwsqnJI9fh4TKls9rBdr7e2i4oZR8RmJ7+HSrYcVmRrE9D/hxN45
o/QJlje7kL3EtC7vzSRgeqbtggoMN5iokoFQoHlDqWzEO2e5R06gnnxKncJrxkoZ
WYPxkUOaTiMAduAQJFmNq1i7m0V5v5DZOGn8iNZqyd/0Ivv7OAgXcvcPef6DRLvn
pevbNvnNj/c6Z4EDi+rBCDTJ80EQNB2TzTgrFcUADHgjoCkNDKNwKdMUQe5OKnPP
ys33AKxD4MIsvZShlvwLbuXAzMfsOZDnYIzILLKlf1pHODi8Y/SFAlMZlTxW6uRN
mNGKpZYXS6kwji334IQSlDRK1MTMHUXLoO1A0+EmOE6ZtrV1oxQQ1Zjwv/RAqs4l
QxDzvjfgmHM/fMr0NleUk8HPR0EEjqyXkExoiSwFcMvpgXHQJy2rrUqXkJMNnQkv
5Cxognc6OWWeL720HW5YrgvagXUOGEXSaaIShJ+vuGBLFUudznp6HJJBxvMN0LRy
qmpmjeQW4Rt19sgXiaQRV2PoSQOuTKFL9cgtJZgaQB7+XicahxsKnUirTOZs0bf/
dCzt7Av5+oXtQhymUw5qs4mgQFRJttYgUpC1hNZozXPw0I1rO9qPHdZO/5SVleF0
UrxyQzgVlbvh1Mp/KRnnbGMiUiUIEyaq1O+9GB1EOAOD/zNn/lHyS5rltnp88Knx
aCHkdEeWMmq4jVgQCwWK65k4heUH5oDwDuHXp0wh/eiU0gYxSi+kRJDxW3QNHJXb
5bFDqOzYs2ANznMkWpfXvMVVkuHgKUneAjM5C7zBai6ElEQ5ABuz1V661tfvmPaT
OwzDTtGU3hrH2ldvXmhF+8FeZx2B8w5osTxnp5L+jVSq4nU1KfXMDOk9ykv9Ddpc
/e1Xb6MXaQBXW06g2XVLEo4o5Tmk2Do1WXvoZGL6kkslmhH72BQ1YAiTCjGaljJz
Ab9Y80lzSA/pFnfm/FbX5jpZIkwREAGc7VYglclDi8aePjutzKRfPZhWeV+jLt/P
usteOVoUbAYb8/jOZXr9wvYkUoAkwz0X9vHg4M68ZlH0JqIoI/u1TCsGwXbp8krG
/2C05TkGqxv2Dbso/mlcMkYTZoFYg7vA9t09fQvlmodw0EhoyCHSzoPCtlLSwTt0
T/p3cwkbM9wY6w1VnC5Tvi+Q9X5KphS6LOLpEC6A1Bnn4CI6pl3XXrzctqV8fQ9u
+qV7dG48hq+UEDaWHE68HHC3vC2h/L7wVOntjUyQA4bYfRV7uImvB7FmhuvGc9Rc
C5O0Q2X+arGn3tTJs00ZZ9nKbuqcum85vLrjWjsrvBgTfRSFiYEN1h5thmkmUQIa
FyM9xlEKEXaYOktsLN/9aidF4dz/hilCnw9e0upC1og5Z4RK93ZixJEs/8mRd7Mk
hE7saAPri/Eukq6pIZgour3J3u2HCSQBHuRrgKHXxfLIzMZs6Qc7rFbQzxcNn4vO
mX7sYBtzrserhvXk+1Xj9jPsJmhfAzOnMxK3uULtDKswH8UQFzN8LS260womyoZC
ZiJAG/nEKojV3ASz/KjTQgjjHwexONowIWqRhDdnpBAVrD3TylxZ3cLVSk+GHJ91
1x+1bvd77uty1IW4eus/AEjgKy018+Pd4SYMsOlnXpqs4yKn7Tj/9uEFW7NXQk97
ELl6DFeF9uQXoMYR9pAS+80GiWMRnJN618E0HHalkqgbjMZ4I+EZghZbGpRZLDOc
l8d3V+6arnoo830RqlFMs+ATjD7BE2yqtFz45pCtwZkLVz4xXAd1Xv2TVaHxrC6W
xp2G6d9AP7PoW6kjLqa8j5nrs7xdwOr5cHMv98sBPIDo33LFivX8rhpwobHv7Ndo
tmtW59BvhOgQpia1EhY5XS+V4arr0GL7mLP6u/0hPzjq/Oty/HbxL/dmJB4E34qE
fYtYHvQyt+1oLAaVmmqxKR3bcMccGU+qt6JijkscWK7WI7Wbfu3KmLA88irDC4kM
8LXngIn95iJjpEeoUjcsgxznJr77QOHOUZaBCDoEYujHf2ag1lE+ABcqCfe4ZPk+
e1tF7tBsmSxJ/3E+/Cfn4iGFUEs9FaXrGPAF+LctoZJUzqoNV62qwbtOcb0wxHOP
cJNlq0NazGwh4WMAjgn+8YyaTZzLF7XNBvwxBK9HgTqHPpxes7nTzVvQpkEcBGZS
H88ARxEsGJdjAbluZb6G9azgpEQBI7b7xArMHVd5Ep7CamCqK8baXiw33EvHweCc
GK1bhUr/XTWTyCnEEG/4AWx98DWF/q/2Ev59YOArECReh+lDenMaWWdKEKnQw/ff
qkDeLLzl7lODSu1NF52ou3sujtU1pLSRqn7E+SL4AmGI10f3zd0rwNJKLBKyDkgI
HulCX2z5LEi5we0QjiXGdZyhM3qA4kLR2i2wTM3h5XPVnujlb7Q9IF2oAPVg7Sc0
F6+f4dTctEbW+EWk8mwZPsNUhEBpPqmB2N6lEQhV/lhWzG3hi7t68//q8PZAJ7YD
s5fG78gUXyYBD+Sl+Cc2mlu5a/xkMwLTTUHKdsxoWoqc+calQ8EQ96iQruHAR/Lf
1wgkYApm98nyIAyy4BZFFDc/yf3aL2UaOG7OwNTZi/P1TkJ8jpEPMICEkSbsfWHL
m5Ogo2UJY9WZfcNEWQJT33b7Bey65L+mw2A5IS3tz0uNzOJhdsfz/LPQqgIgdIJA
KTrW5VF1l4cKHmYgJfbcK5ivrzXqMTOnK6CoOUKdY9B0zgb4UY4PuurGJVKa+Pjr
oJ0Sg+xhzlsgHn0XhMpa29z60IrWSnGpjJWuMJBH6Fu5QZ/26gJKwWXBI19NU4jv
cyL1u5VmneBvMfetLMc5QTt0FnEU3qJtRur60bc5qYddB1uCMu2cFNwlksKUxDJX
4DeZLM7KT1R7hrnoV1w3iqjcf/+q204gHrvUVyDIiJpvlmMlsuLUnDrCEsMKrF52
ICAKZBFVSZF3nDZHDkKO65R2Kq4RQSY36Oiy3OvIWKbyEtYTuz8BjIh7Q1M7gXnK
ywxuos/VKsgcAZzD49RE1woQmHPZtKPV/CgXQcbqs0Ogxbg4OKz02GLD0AmctB09
bJ8+9zQVvROPVnEx0kxMFJZlspIMZqNYvJN/PrFeDM71p7HlrdVSeYl5zEkx2WVX
fmbyRP+5nW6gIDaSNOIlLDqPKPfr12HvRUHi7jdLEN+/80H3W1yce4B+7jZHeFcL
RH3bIu7J/Bjgk8Ie0J+QUJNw45jk7WflJPq7osC/RHBKwPIF3dwwdFQHLwLCuH4C
9zPnkdRVCUCRJo1kP2ZURnNtCBJSZu+c5dioOdQhWaDZeCfnimP8nlg8jWoewVf8
6YIhQM65qsFhViJqLBf3CiqpqRNwmihXyA0pwMqBVZivouX8hWJ1WL4lMRsfQwmP
mOESPGw6OITFt5Trwesg6QxI3pM2sflGtvSwEs8ymodAOD3MORRo8SqhWEBSsX9l
J2618gF3kGBeNlD6arEFoyn1++xcboBz+iBwRomEzG3Ssjv/pWNywn731NJrJkIO
RqOsqh+jJ/9cXiex14DaIR9vFG79DLmUENby0gD4/dec2mPa9QpkZMecWAD2/NYt
GS1Tp5McwbU31Z2WNXIn+zXn+MuK0YtWjs+BQwOCDePsP3QaVPvzcePhdBNJdVs7
dwbcZoT/Q62OntAPWpqxp/lUy+sWKlZmNoHGXS7I5UuTFNlgll31XFf1Qc00K6re
ZDGNWXOCrov74qsmG+60y63MgTLs1kTbOKW2WwJ3NLGqSw75kTis59bXKFtubMXD
RdzHIVRaxwF9Gz0OypDmqLmjgISiVSMqJRbbp0VYI8PoNCuQDQGthQG/hrQ2KEKm
35t+Rkpg1cboW1uwVWuz06NCMu4Wg2uKd+CSDoM/Dz2qJ1eSuK1kqKeTsm6hRyI+
/HdiJuRPSz0IvgYfRCA/OqfpjI7BtCmOFYYTprdXghkjZwvrvC1OiISjIxKGIxZo
aT2DJgUiZwevSdEGXF6Q5cW3WNjYb8cmTP6m5D4itGIbjfKW6UoJaCvtjW3THMYa
OX0VU9La302lrULpdzAdybuN3WJ+ur/wN9msXli316yjsqauyavNJV33ZsTy5RNp
AdlOf6z7OGb0OMeLcOjDo5382cQACDFxVC6y2TVFfw+NKUuIC4YTfP13z1/sodUj
A8lH8s1SHbYI330UwIn/AH2+OBp/nS3ZtEzy1jNtBcf/3PdTrwm/p7RqePjLix+P
yqbshYUfvXLTmJTMyV/PcfYiFGbfh6Z4bzyNxeQHktcpS70jvnBMvznIJuFvrOGP
G7TI1BtkWDoDKuUq6MeIy2EZQ4jU7TovsnFRwC3NMFpArl+Z4Ye36VhNVh+bWrbz
/n5DvC4nNATm+3VY4/TW/20GSq1t3vnzuO7L+I2NLf3Js1n81FOXpcj4LlAq0J0h
JVpDyrvEcgs+j0spjfsv5tSFK8H7PGfJwwt7+BrhsBWrVu6xPdRsxsEVWRUCGF8B
5tgHze0VbaqG6jS2vnQDP9oDpUMAEIt8Z/1jF6ytGdEtuGHqo2UuqoNCDVor335L
TtgFLjSbCSgniwl8hEQ/p3venECP96RXoGLN1OWppviS5EyYRwLonv3A+uYFIJRD
nv2JM11Kk06t1kGQIRK5t3tvXzWWN8JeHbFgOlVgbaEw2XRtWlqNNKMTise7b/zn
/tNevJ0KwzBOYX/9uHT5g4rHvr9cRyDIqaI95HHCz1YbqyuQGGVnsYNlp8kko3GC
msKEqoTRDNr7npqK07Bk+Otpx7Vs4Y8Xl3viRN12tmhrBjB5lFn3D4gsTQKTq3W0
PkMx3bGMTy7aph5eX9X/7Yf27Sy1mUg4j+7ey5STR0usfjsNKZfd64gMHwpdg02H
tJFuZBXp8ntpmPnnu0zYaXwr9SvueZdHtGGTNqRJQbeb3V+he5IFAiaGptX9t1Vr
C9f6rh4RtD1Npej7XXzyP91myKTx69bcRiPDqkjpveiZnwQj/LqUBAaC3/LSJ5ka
sJg8eEJHkgnMFad6rU5PJc2AqtpZmtC+D9F8YIrL7o6UKGU2o01b8W+4WrUpmrF2
phbrRQ4IBh3YLJexm8vRENb+dD9H0d8YKP+dq5BeIvFAx8H5sgjiaLjuSYlNprBe
GmH7SKeK/38x0/03ZJJtrdEQ7eabGyqQ17VV8ijB8r6jIIlH0errhPTWGdgRlckS
u8Xg49sLg4kQevM+avH0jH4/HRQtgZ1P8KMm64z5dqtLUMxnzHtn/SZhxHREurFP
8qutwRRJny8Y1BkCJNG7aYNygehQjTVg7ZcQUSwSabFf5Kf0PiY74+xOCNDeWBrs
vxFJLTFQQz6oTZMdPzk85FVpL135aCkBX6+ebYrnNSb/6THPE3cCsvMPd+vgAmCk
0cRYx6c6IXdJ6vYL0dYyRxKZ52q9opQenfvz6pXDuEq9bTGHwFcDvxQ4rSRrOlcu
+/FXbRqmaAIHR9SbJahWw+M3bx6kchvsZkpUpOMOczVOJnmmWpP3ARzNMTcLA4H4
aVUqHEp0EJzUFlnSgq8z4QpAfUJ/slc1cQNWLKIPg3EGPnEWjHql7V6nN89+L/pG
F4jUnTX7kDbnj5C44CyV0tGwrlIWQIzK2S7P/g5ZeWyJu+Z17C9W82hNI1TjSU7j
PR5CDI6gcmoVAX6n5UP57jRnNABcOWBBbuun5KePWk69vUrX4oL98B6RuThO5SLh
cB50tG2SKfnq6GmjidsM08jbvjcV3Uw98RfuXQgPVzAEdcxPWuctTQqVLV9Ob7iy
QbeQYSiUNTc+iz+5OFS3FfxvpNI19pfzEkE/AAC9vyHPgMUqOILNqKrsLTv1ID51
bXFiZplvMeKXkpj80IUGVEHQlgBy1vOHxK/rlPfNK2r+fsdzk6I/boNU60AknyBw
7GHrJhIfOlcZdcWNDW2LxokvR3Dx9fLo4HYH3zEBKi27QYZ7CaNRas7zNPtVwtSY
NXmN1QphcxOSJgUuiXwSnRYPnOWs37UPXJg88ROzrmlbaJVEk6erDVEPgB5Why8f
GJuZakH9Wol6dK90/pBMAKA75IjD8KwcmlBVf//bEqybw9gJiXeyntEc/C1tU2cS
h6/2UivVxlEsAGHuatmdUhgTbz6n+P+b/o9XVTOTvrehB5CmmUGW64OHPbUcpoDd
QBpge5iPyC85BFG1sB0q6rnZpsD5wevKMGWr+O+g+ZGnnzEH8koJd0heICuhaPph
sSROZwlupURL7o6g6ThRWmR7DzH6M5PpC0BoL0irzSynfxgFrFS4WIYEUrfh3fx9
vVf3I+rFzyIhJxvaH9nrHBGa2PmQZEb0Ku+oeJHrZsJ/NMlG7N1uanu1zvYh/9bS
zA60+lgcEauASaXNEje/5SZzy1kbWzDvtU3+Ah+IkxhTz7JewmFa8+Bkmo4nXPCk
zL/B/GSB+aZZoWv9kxkwXdLMo/YG0w2DCdehTqDsRdMi+Xg1nL0IF8E95FGvlkmO
2ZUeQJLnbobDTNTvxXHCwJYqMcKpgFZ26ArKBPhLQ4vwUC/h+sIJinkrdTZ2Z+7N
E9PP7CnJpoqPs0er5ynqb+O5ekc8EG1176ZBmoSMzQVtwYKzj5mPhYUdqOHHprvV
QIu07tIinus9ysQarjfcrYD5xH+XTVqkJNtNPpmQc03VMK0xwFOpwwd6PLCydFiH
lugaf7x1iq7c+W/HSh1EknUMbnGQjBx09z0LbBSL6+a2R072NGekd20TojASMfLe
GgJfL7cUTvrxwjtqzAfQdujhIXW/BeMEmkqP3OjMEyk1J8vd4q1ddskYXJsrXRfQ
EdUvmHrCQY12fu32f8UhN+gOoU5HIAMGmeOG2V9Ou7D28F1cM6H1P8+NOlm2Nfni
Sc4z3rWgx1I8ku1/IdNR9vTdER48v0tJrbSAefwEk40KF2m8lNygRfcpd+Zw5CXf
oeR+z3OCC9fID5KEcObGlp3sO/tAiI3qpkCbPv+TwWcctdatmwyA6z+lqmDCUMg3
s4sQKWyCH1E1h7/lDF39ERAbXrpPYgEtNP/MLOoxw+a7lPYITqT2EXT/x/GlwiFw
OR8w90B4ehHP78ZxBDtfKjmT61SKS/UfL+SlzTSG7n4fUwoqhrpRqphBq4ZQZ7KP
kxvm+jOOb6SQtuSmDmX/sH3+LdiJ0PxS2I17JzfEUscKEHviaUAE7cdiyJ215m73
62Zop+E+bcRDPJJfvT5jP/JbFjkAlaREMe19ISM/oYUM9yy8RLD0ajmzrZOE7gsx
7+fUB1+wJUB21TA75Z9/flESDec02xfrf/PDZi1j5dZ9oz+HmyrmxmOTK8AM0Usn
v2uvW7XroznMKIZZ1Zx+GmlJWr11oP/ZXE3HWoZI65hsHz12Iz2rqm4HcLfIEWGC
nYp0bOuMc2s+wKfKVnwSnW3ztaFMFafsvxb8E1plBkCT11EgLtn2tTZXOst5O7YN
Sc4MEkkcK+qdh+LG7P09zuEB2re0or03hcPvwy734cxrHP2BGrSQVw3FuD8D4UtQ
8nCmQUSNycw3JAoRPT+1SCoxSRh7XtxvMhMth7YOlr8ZjZfZUJz0PUeVy8Is4QfS
+ECooDiKoDVCXRrJk3q2jSYua8Hz0GYOM/FEFF3dZTqpVWSDGSWGEe+7psuLOix8
QGrXwobxHtoAAgBpKnhlxqRM9RkKCGQMW+gJjQr4/XRQgevCqXJXLICHgPXleRv0
yEfW573bjNZEtnX/yyTWxnkRWHgr7a9DvFdzz+g0G/JigXpdTakVpwq4JL2jwH+V
UnKL8eMcSpDusYQXUOKtO2tGWp7xiiuhH53GruS5o/1lsjmvvjudCUcJcXYUcUod
GdajO2cuCucjQQHfpCpu8vLZU20SUNLgE2dhVtU+347S/Vv19KbbYMZNnTGJ6ris
xscSsDzTOHESSa+1GvHRs7u2+iQb0/s1QR6+Sku3PFxYq7e/QrQnitWUs84UCI5V
qaoz50lUHqD2qkP1eNJTj7qDax6hb0RCKoSPybcCEUNRUtTZUWqdYhwBdk7+hU1j
NccfwYVgsb7M+h1sfZyAGxvfQDCre8jJscDIhGfHqfyyaZl78QDPljVdmWvsEp4C
Sk1jD7jnIwb97+r+G35rYhH6XGaNrbBpWk4IgUmXDjCtYAK8tpJgtkT8At3m/szs
2u7t8Q+ElI6Ya4dNQ7NdWb9Fuo2+yjoWwjDOTFr+s9auO7v1Mtd9bg4jAxwlPhk8
SasRwJvOKprPK/zgkTh8O88/zw/4t/7mWg+SmdvkgEYhuzBzDOpklfCvofmfPgH7
b6yaumeAqOb4w7EAnzdRgQ==
`pragma protect end_protected
