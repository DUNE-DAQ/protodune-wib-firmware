// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Tpat+VZXNI79b/f+ML8Ug2ZeTZViZS6xs/z0I3LN+FWDdZzoWvxPk7a0uwSS/AXW
MyevrF0St7ypou37UZofK18QO6n2x88+yNGEFX9seD50SXfuk1BXbrcdX1hi2LZN
r4QwJXgyoLSiy3TdD2Buqj4Db9ouanw+KlleWt+hd1E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13104)
w8CRbpNQjnsKttdBaC92DBtLsmB7LvYcON2UWkUfLv5hIZ9HEwMn+t8wdMXsrZGy
eIDAemHMv7emjcCcnUtKyAdz9v6WmOsxztcGSQSoK9UsreatL4ymNqNAW0M5cek/
+7moZLWz89oQ0SDso6+sPFM7LFOAtpVYW6I4fjIbcY22FpUi7NrWAm4i+fM79TN6
gMTQ5IcZ/jwjkhSbbR/0/IGu8rm4qhLBTWHEkZwZhy6/7in7tg9qLMtCMg2uLYjo
v9Pf/ZbdTArPEmjGB0837bjBe8X5O+8KPMuIWG/Hss3BnuhdHpmxXlTwR6Bawbwb
Aaq6AnMDCdDwtlKvFHCZMrFftxOP0DTD+802DMDZ/WDCPFNcRkEkgIteKwKeXVWx
NAGylivXx7dEjjsRXy8/e83PM2+w5KRYzey5UNRCja3W2c/ZKtG3oW0soc1VZePk
wX4LJJGjKSh09XXbkiCCsCxgmGOswr+x0lmctB4kshUJOpS9KXMybLjQXd4d7caK
XAwszPDn4OVsg73elM7J643Phi8YpsoIV++pGNjNi8w/eHofrURCHVZHr6pDrY9p
8AfWiudGebJx6L2oZ/d5v+IZJJnq0ZCdANbxuhPrMWgXG31nGkp5YmRo6DrumSQ5
g5J/OssvitK/Dpq3CXR6cbbniFrDJ2NLq39rr/5kzc9vbFzoMbiwMtp2GTkFL0pB
RUTUzUoOVAUPjqDQVWujdQcKJOj0NYlqctjsMW3+GLxkJJAj78ftqQQXkHwNlUdd
cVvCz3MO5IJXldG1MjNc87LZ33FipWVCyXLl1TXNPYRKwpWH94WCvTyLtEqT+P0S
01cqU9s0Cq9FvV4EdhNXiaJZYs0ClINmsYWUGbRadgFAv4cTAYdW4VjpF2HEe8Uu
vY3oGs44kImUnqFm3+qI9bOyuSD8XX5d996ZEAXQ6vo3FhGARgqKMFiPyj+cOHO4
ZPuY7ZlL5DdWKSLx8ps5FORC/Tkm4TcSAeNo7ylVK+InP/UWww0UtatpNRrs96jz
rcmUIpAf8UtV9VFw5d275GnSGmCTDwqBTjJr8gRHKYWG7Z3t8QOZ3aYGAjV+PgwA
jr0FlVZ5EN2IWagMHvABg3V/il4ODlY0ghwBt4jYl4vNmMtqpaUshggn5mecenCV
4HYxngyXzozGBDDcTHOxxE4rQki9X8+bsPjBE8KOBP/AcMqwlzJKJs4j6d8PYqWK
o3PAdG7c7lRNTuQC9UgP6kv3UIb3z35F/SXGQJA2jdJD2EQ03MJaEAFXK+s+MyDy
fZcx9CvF6d1lQ8fOJeRG6vYYb0InoIX1buCuqfC49FuxdWukLaLb4ABgeF3ITbrG
0CSbY98ppDah6lwoNN8zQUKpXNoyaByoemFxfM0SCUBelEXYKDaD6VWbRV51wkSK
mfPODckVZ1D9tv0t5VsybEEdeCUGipBW+rzMOufVPb3F7zmwLicOWVB+q7tPYzvn
UCbVMOJZgBBZ6DlGKbPf9AxHMlH9ymp4w1PBSm+ZENld/ZoUYhVFyogy38xAvdXM
xM9GjUnQfjkSG6XfqjT/8HiwJI0YtPHRQwT/cpv3Pkb5EOajaUUEKgVBFjYbJi6I
M7RcgDEqnlFLPHgrkbU2yXpAMxMWNse1UJpYuMwnPTZX2w/icQJM2in9dNJVCEej
kI6BPWdillxrCQG48wjFDdsucmx+pO3awjFGQoVZJbSHsm0uaCIg6xMikzve814z
mDOTcXnclhXLyCwupblfHZlJ4W2aJSjgBhl9bAPCqk9+aFn9ECJnQMkUy+QJJFLZ
bEtZQ2kiANnv5E6IaQfH4vnq/k0nBry2IE/r3rmSqAanXT55fHAl62reA4J8MbFb
Pd77m8lCdfh+8zD4w46ee7R8+33CA+ja/z/795AP6PObOASteLS979rhpnQJe0Of
R55+u+o6wlBs2iiFNRlNftst/m6SHz7ay5sxX2myjmXEwBpnem6UiQDmVFWut2Ec
lcC94pDOfP6X/pTaJpxFxJQk3vvaT6ISrFusIs9GWzw6Mx7is6RJiCietzOif3vl
Vx8swltRvLjl8r7enHa4QSDk4/NVuNTRVG0QuSBiaa7Ejmw8ztCKJe5x53C80qDh
PphFBjLVOEp6mp9YCm2MFsX3/yY6OZsq+yukP0vyi99OqBcoFyDU7UuQ34Nvw3p7
pdWatus2ru5ao3XP8X6KnMJCtFwmnfmI52wVw+paMwmfDg7w0hZ+zmWnUrjbltky
s7CQCcbBScUx3+l2dAwO1UeWPNX9GqD8oR2T9jlT6bEAknVGuY1DrHAoPujCkSAh
7/0tzsshKCgZH6BgnbroyULofSQvAgAC8/wXxxnYCRxXkwUzaYnkxk5AXN87c7f/
E6MrelhZ5Qyvb/nYT5LRZYrm/IaC5N3Sr8auj35MJl+4yTaYYU7bx3V1SN1F46nC
g2yDMyyntZMLqvXGAV1qh83FGp5BMZwZDH3kZLrYdbTVXwQ0UYsQ0rx7sJenjqFj
5CdHk3MARVdRXAIPcxWY33uf9/RD4QPA3To8dS1JZ629SbCqC8W2JVWx5pkJHsQA
7s9dyftUrVKBLsC4IYAA1vUIqMGwf4HQky9A5dVL7np2fvmjApuZp5Iv6Nxa47aZ
OVS3SSiRUxgg1WoGo/kJowg0OSBSpI7YDEXoWs2bJMUEuAZ7Vrba32V8kgoa/wxW
Wa0PhEdxyQAdBBB4QgCT+tTkhejMIPVs6Rp6iIG7F8JbC1Ebqy0eHX7roW8eN3JT
ME1Hp/vqDrNzFlJzzpz9PwfLpR4FazuIQ9Sqrzg93Y4DmRAX2lS6kArEKCBveUOo
KADcn/q7MBsKGdOMVpXI7CrRqL+1aGMBGRh+V0RCOMmervnT6h7Jcns0tQWzOtjP
209kmxpREv8Rp9ulr+yb0cLua1OWf7HSmCJy/ZpFp8B+d9DNAVL33zmS2XciHpkS
o0iu/u9ec52SRvJNeXPqiVPu/eMh/n4UaOuV5ra+Qp8lcNga5DR7C+I42+s0qvNZ
1vkKTmH7Tl8Z7fwvuJoqJ4U95oUak0lHlnlxY0nx1xWZGY/osNvSjtZsr0oEgXK9
Yrf+0DUEIniiwNM+uZbbo5izqHwVueZtus9A3RA3imYPUgSs/VBoL218vg0IRtII
mI4ocazJo+wQI2AUG5IUFJVUbG45ihIUcvljPwZIYob6JH1yWN9bA5UZXhaA+qF0
VDJQ/NA2gHTlKrldCKhNRwIMyGgkYwNITo9WDcxwZjhRGns3jLdHw0Na9R9x5OYE
z+xvH1cybccZEN0p9uo6F43Agw36jfDsirWBwhoiZF716HZTh0b8eMN3+my9Py4Y
FfHBYfNNyduj446S7CY1C6Vf8+bAx9IReRQeATbwmlTmcTVLzU2Y/7/Hi2TKpHv3
3s8QnxIrEdH1/Sj5M8vPugGwILAmo4HB4REW6sWUpiIWOzSx6k2wVybLNgwrfCk/
zWVrJbY01znUJhbHgUQWwKrPI0micOfv5CD3GUumxmLrpBBX51ZqoodhXdXh8IXh
UtmM/+HheXHR7k7EqFiIWCGHiXIyQWyjpOIh02hIj87aA4st6ppMx9NyFNlut25b
WhfULlXmWs7wkm7OyaM0pCf95/pWHiRVK0ZGF0hD1HyC4QFuoGNtR1cxWwn/z2A3
88A4adtsDEmsxV4u0WTcULpmOV/cnZaoc+vErK5vWEEXwtKfi8mZ7xMgpGqo6oJJ
cujqa+/PP3flPTZx+ONvD94PB+UT1gjMu9uyvKuISoAr7bFq7e2YnTqlyfgoskLA
uRl8Wkv6gzgiZuoaVuw23DeWbHBdpcL45fXPpicAHiG7xe32JMVZ+bfvJ2Ys1R8m
kVG7MIkTC5b083z5Vwq1AWT1PfByp7aabCHWKEHNcWhtsCeOTbh+k1VkX+cwD6pG
TiZXfCXuZ1fexPV5BfSNclqjEcxKZWVGXexpfiZnGSrtdQghHb5ngKb+7Kkh/sXQ
137UFmonbIxG+0acbXM/WjRAMCodnBcmGW5qIK3RTsElTlrnXuEukzGuRR+eRSoi
FogGaBd1N40NalETaE+wjfr2p5xJ0AhSPiAvFfG75LV6umi9pzXjOjXQ42/PJS0y
Vfk3lpUV7kkmvaX7UjuTL60KQCRZNCe0JpTK4m1ZweVqf7MDAhXtFcIrOLFabl9E
4BshRIyM7zQXfqE64cuPgK9lQfLbvf56du9BkcOscwBuRtSYU8nqwY/UscWL7NF+
6O4wFut3/mp3Q0+5tb436oN9rhn3rk+W/PV3MbQ5R9l5Adtk5LTtCR0KIxwcQnn9
flm0QhB5T0m2jvYuUxfnxUBhglA8wHyUepUa7SSC+k4pM9DcJBDVD1WkcFXsHbRu
Rw816qBHdxFRO61W2/EfMNjdQgNs9SlWAH761ztBXN4uTapHwtYVZuhMIJba42nJ
h/DCiIbyoMxA6mulMELkmEx74pKy0YJKw84ll+Qc1PCtsP95eOrZz+B0qWL+Chib
ivXeH1ywGmLVAE15rIdt7+RQ5jlAmY6Xi6cRY0y9ypP/kFFBrxcvrKDNSbyb9RlR
NMFS97DzwkVnc+LeZy7b0VXzBlaIK2MUwi8+UZJItmQZdBaewAr3Kmh0iCLetkgd
rm38cZGeSXYzo2xX8VryA8sM3Xl4+06cK0KZU0+slEwa3pkQ96kmnF11Xtj5iA+/
/1JlSszR5tIUY9j3EpDa5fVK70mhqLdUpSpCkLoDhB4p/e+s+xhEFhusswsydbbD
dZmx1Yo6QRzx7GVmk42HyvhUSOHtWMJnEajD32AbRe0i79ai9thWlKzx0jXeUR+q
7DlCqezDetJJd9xlls3CT33+cTwuNIT0CYkxpVYNRvE3r6+kR8Zt0LrjacDtReUi
kV0aQWHa0ZwkdaMzkWlcv77rnH+sZUa1OBW/hhEf1ci6KB7qhS1qZWV3A0VCz2cG
zNRI0Y0kIr25cP4d2VUVfa0f4n6EJwoXrspv5MW38AD+S2sfkg67EtHHjngNia1N
tNR6/tWMJP8dnZq1K0r33UMlE0+GGfFn7eEVjLbXp7cSn/T6IVhrYq53zCxNyqDZ
TSkIKZIdluuK3rCQiHmWQJDeg+hbM7Gk7OriyOn+Cy7jIUzy5TidLAhMlBA22Ob3
ZO/3fm56ZbVvnHJg0NONWISHWtNukBxsBpN+VkmckCJYeWNla2I43rc9mUu63HQr
L14vXZmSZ7k+d4YHENHYtbGkZ6JlgAKz4C6QYxxqapXFSxkK3AL8Rz5sFtwpxina
PcDZ3ViyzC3ziXglJDlC0OBi7mEAdKNxXC9MjGKYPzYDROkeyhz5TAFPfonu01QB
xy+jNaKMGFKCZZMnP/dn1r/dCbGVk+BbX1R7zcDwNhvd3840BpfHqakZM/T5/BD5
q3VEophmXXufrYGqtY+CMrmNeARyqvD3Ai0VcEprwakb+nTkzi978u7YJwq1H82V
Ckv8Enfi51282H51AMUuzSDYTeVuqBvpmx573ZLrv0E2E+tGgFurOYWof6Zbw8AB
NJIyZL4UXqrwhODOTQb6gpfxPAAGJUeem+YLJPk5WVU6MKaaBHn9sAHxVIMY5BcZ
H/W5OofmHV0U0mQjF4OAlhM3mMHMdU5U8jzdkI6XAKZ+GfyI1KTZCB/HVuY1UEBy
SkiE4cXZDS2wMt5WaxGptx1/nj8IZAN3kakLh8P2VtIm5ZmXRrSJVMnQgqZ6ue4G
UsKolQxj/Y/0pAm936ZOksFPB5dycvd8IIuG5sqjiClv2ZoaUWVaZ84TOLXb/Ojm
AonkZUeBLOC7vAqWhasUShKSrPYtKOAlQjabqJXhel/C/zPuGWBcgJSuaZ7zztoP
wv18TpPlCRvotAiout2RueelDEEHgzX/RAE7nGOXzuDgacbw3gj8M/TjU3tknCAG
jc4hTUCLRIehQEKcwGZQzBmryrZKYH0FteC9jh/F7aX+HtqIp9q9VHMGrZt0fa4+
omxKc/qZvjfmhbwQswZkZPMnO5SIk1/qIEflUGt2Ke9Z7Rv7Lfc0oxjz3oVvcidi
XAxuL/TZoGY0KyVfQKNdcVXqaCoImmRlBeZ5T6gCw+6ydyBu7w0/6bhnTijmZhXR
As6CkVmOzJT8XFZFaZHb+/NffC2pHR3GkjnySLOZN9APpwXLI+aQdgiKGn7xmRa4
QTRiNLuQOnUMj7bFijqmCVeFk0v87tLtBaPS8X5GTadwZDnPTDgWV29K91BNEW0Z
2Cd6kDHp2hcdvwZw0+N5mbVnHeIc9TXx9DyMzASNx0PWu6lZ7y60FtMyskVSdJB5
6ZXSIiybH4W6i85171n+5BgOiOa1AVnaEg4g0DYc63mi4spAH8hJuHEi7qwHzsLe
Q/hTBk37P98qsmoadQ6oh+1/sZBAf34yq4HtXhm52GiJYFQiokYjm8hvvWWdSngS
KFonhyt0hDhPLomm9njYgKh/glksTH5tk9Jq3HYo/uH/OLkv3z2tbgBfqgsQUiX0
K/EwARAl5wQQCIalpwy2TBM82DvYjIfuS2X5KscJTTmdYMI4gg8ZGLtdNU3wPvCX
sqnQLpI6IjjuUAHPb0B/ii/9CWcXdOOC16oupN5ngcYtxuadvxVNXTQZl6az3NcO
pjENdPBAi3USNLmkcBcoUK6ogskx5ldnDyQ+eDoLu+Pz1Gmc+58lW17dWq9n2vfw
y9L/QN/WHMEeSYdrah0L3g6YAgNKx7IHSpseUjNL30uwSbn7dUxp6iqnaeTh8mYu
7jBG0luA3eKS1hgBjWVUm/we7ZZMC/oMTJdDJ7V4q/G9MlxNh+B1ff7pXLeKk7bx
s3VdPGqQYyveJmPlSlAm++rbjFKWeoiDND1rlGfGCt1h7NrAeAr/gPECvMDfhdHJ
o9dRvTI65vVUGAm4yQyLS1so4MIFUIGxzGzdgWuI3+Sb0qV12sbwUoK0CrhINrm6
7xybDO8fffB8CbneaqAQRLI1MebCzzQcW6NUmfi89hsKLP0lLQEKwK6Saj/4gQWj
BsZDj0f3Bgz5eJMKJhl6+kSABKpGASdv+eEWCrQJiwlP9BBqqWDI5/sJu0SWhotD
TSRy086TL4D2Y+tG/OGVGll1Erk8sSUP+w5hRaAGscfo+C3z4xvS/boUl6oCJQPg
aBIhyvViZ6B/Bn2R8xJl6TUk+IP73vigGQCVtWwVlP8essyUgY4TQcyllISf7Nfc
w80TWsjmRHIDxEC9y3JxPiVdyqIPFK61qlez+H9JYNyCOwJUJlOAkHTWv3qGPg31
7mZKkMWHzDfJnX3YL0I0NQF/zBI5ofeEdyFnWJaHz2P6HZ4uknw0lEmI3FPmzPrR
HdZ3eyuIIWeE3uKB2sYCnKVo5jaE9tnm9zaJ4fCmTC/xHlZPix3Sofca1ATwdO5t
KDjadbK+IC9QP6Jq9s8mhzWpRETSt8Yb54QcUqSm9EGOTYncS2guABprzaReltfE
umP7dkHB2nn25Z1wz5gkyWP4673FMo/Hz353uvUc9fVaF4PeMCM6SARDUz09wfr7
hQAEMKCUU6eqxIfw87nXcU/6/d7CTEcvqv98S1qaGf1EnbB8JmIiydZUPtsnPLZG
Uuc0M2leEGcvsJQnwtOz9fCwLst5AFWUd3GeXY+0tBO1CkRZOudueEZgmIuDqNGB
EdWu50PdJHA06tZGOXx1Z22tIEMPKGMxFdyqS3P3FeP3Pj1FDBKDW9wfd2/2M/bZ
cKX9jnumQVW/SOX+96vfNAxA/flCYrmru4Zm5+FC0Bk79tmspYS0yNTHtCgIk074
cfjhgfbg7tbPsN58RG3gHMT1/k3XMWCyUX1r1KuEhE4aIXQOsU1/rZ1pm6El9H13
vtrPW/aoqHkvDq36Ey1W68/A6g/nkdq7xGLDlLGe1scgNvpjmpbtdKblsbX+ICsd
iUap4/eTgnQTndM3DV2enomyofBM4RdC7/AQWuBcJhGlGoN/n3dhiyEOQ2TbmKDP
4wgvT3E/eBAStMuxWTlTtQ4pRlNjsN4f5gPBXColw4088pz6woUT/fWfkizDmhCq
Xp76hef9/1+JfD6Vs3LD4sloI/Eaejsj8L30UA6prlxxONXEfAC2ASaap7X/llE2
AM/O+8CrRy+an3lJavhhY1x67Ktfc1icIyoY9z+V2x3j2GZEQdUER14V/hziHxfJ
GO5iRz0BcgwHrn92dB6QohmYD9PjlL5VyL+aGynnsGSJh/vxPcns4Zctf7EMLBGW
ywC/J+2FEae0IueWWP9Lek4qCPy+9c/E4kbdEPBViQUmku0V/fAl4A/HZfau4xYg
BBmqFClBumzA+q3/2x8pId2d7LuTf4ZVeAyzlOJjUlXRH6sSggCXzxjBKbcHZibH
TAoODRyUhoaYJN32MwBEGXjl5HFxEH+UbJ/AGrw2mupeZNfwfceDz7U2cVRae1nC
jlbWK/yXAkrC3XBcPvAWzkdu9zBw1kS6KnREL9DPJq8mHtbMR0+Z+gB6a9Uhu3Jy
9GZN80seuNRdW2LxZ3i6fRTCBtbBQ+dh46mxI45HWmFUXW9nR74OAEuUNTvpx49l
LfDBpeAyTw7OUBKfL71ESeQfnr3Vsn2pAPpbIq4CxisMtPJk4lRYNaEI+bWoR2Ip
ulAYkvUlorleWXHuwL2ydslsu7DSAAcw7SGveQ/ysM2YUQBgCi5lhbHdLHlG0pqV
19vHSo0ErvDw76i4e6/LPJMm8ttUdeqXb46v/a7YHnOs3lIeizgJSm5zJBbFNeu5
eLln/h/o/T3ZtWInb8KS5X3RmBRP8J6+obSGi7nuaiWyDdqpjRwIw6BHSOOkYS0D
7YJAXzqMCOzdVC1AXr53nCe5qdLWMm4f1FfZSDkrsFXbb5TWMs+tnMJ9gXr9Vh8H
l60R3RweoCUN39zZQcAb/Qm58mHY3yQXYtu2eHL6oJJ45VF/eofqclgxhct24bLl
DRHO5GqjaxT1Z/D6zRPUMnU+Fb+yzhclPFS17r+wl5Ak8IkQFpxb/Atp5oscLd1h
k1n4Ale3QgzGqBrzFdFGkZXRDuwPi/Nn0Th7FPSkPUXxmahz8i2h6iE5OrMNEtRR
FM32baITdfwCfo33LlYKJeU+aqkqsmr6pUvKZ6kQclfeSWjm/50oukoqfJ19krVe
tI+B7U53euNM7psF7PJSg5LzHd3WVyVeAMRjw91rqCnsoeCGB30ItQTB6XerBtbB
3e+tLO48j3H2cjWn+jtt7BbIxa0XF7KjkJQwUnSW79j4WnEhhRSgcHWDZYcby3Ad
HLoSe/mUbcFky1BHlgNEV2QPJjTxuvSQC8F81h9GQCg7jeqN2I66PGMaQ2lW0iF6
rxmhv7rX63y4OGLs+TJ0UBvbDG8kxdjIvv7ufGvZd8wKiYJnja7fiOqm9r1ZZk3L
9B3qwLIAIFB777hIOUqyu0CefqAePSFTgzatlGWK/6HxSjaDhSWcw6ypIrl/WzMm
yam9HGQiugsJWGr48EVIT5SWs2e4Rql394zLUjWbtO0gkPmNYwqMqRtS4U8QBvfm
K8iNkQqHsEfKZNG6hU5f1QLvldUNbjad3eApRnlXCZ2IasktHSr6XsU7ipWrAtVD
1sHEaWxOqEJ4nph0wyPV2+uPNGjIal0UYh4mKC2gCIwsP4naliNFFe7v5yROv6Dg
tcdfKRJ48+YlObwVgLOzLO9tCKqcM/z3Hx7xZcWuMS2HZPg1uVp0eDwkt8zY3J2U
3zEkch/LCtVzfZmh4GruLk2maGpYm3DCRAsg2KqitkMCzetOctgKl5pQ6DBq6BGb
R8Suohv5Q6WLm9kahlWdNcGDBh1/gjwRgsNM3mHZeK4tlsqTx9sZKMOyySRaMQSr
us5Ioks3dIcmTNyGKAEPmnnvWr01KbDOUXKywzydvy5RdZmBJ7d1WCaUJ7AJjtsn
kpbfTlSNYmYjXixSdTrM9PXxC9CJYD+T5Gef6l/1dlEAS3MJRxOYvOWvJnEtlote
dpJcHwbaYurPBCUmhfE7ae9btbz0gnSYD8tjJgh0epUPdSwOWu9It1G2O6+HVKX8
GP6a0nMu/fle4X1InfnPckRytv/u5dpKpUTwmPi+rLEc2d5V9xipHzaKLsr+EXgt
o9xYzzIAvkT5y+G2V5YEe5Y0+qTbEP1VG66/G7ilooqehij4e6oW2Hbs1YVWTRkO
BDgn8JgN8N7wytdXxWxGGup8jFkwY0qJqoE+rBrOOvh99QONcZVZFPREM5KtWoYY
eBbY8Hz1Q9PqY9Gx5Y0SmmLbkeIPLbMvWnnEBwssP285tYuscQtsy5ighRKwiZBT
fmcy5c+aqJ/ZpDbzJ83NnlbX2kKx3S1cFZ9U0r1m2hkYlKoLPs+6YFE7xfB9wxlr
Xb7wBngHiUiW0gcIinkZtoipc5f9lOkHahN6I+aLbsK0EK0yK3saZOVRvXlR+2dH
F+MIqul0EVze9IUTSe9qWd4tGmbJNFhSC+zm5RBz2vjMkgbvyErzbeJQ21XNSn2N
3MuUBKfAWfEMMDNG79F6k/tlRgiq8H0rZ+359MJixoX4C/mE3mE7AB5n0lVjobQ1
6v+IATmGcbih6O+aOU5lhQjVP1bEllW9RAPYftlxPcqGdpnzSTC41h9uYB1N+stT
VqSx5J6gOfZX8F2orGFGobQ1LrMT74m5XWSiSaFZzJ4VESnmHX6op19eBge2KeD2
g1EPnLRIEG71S4orJeQ0ECOlA71SiBUmfXkRU0WKdCbcsbhBuhf9sGuzkzBkVnX/
270klmwW7jrPIbfYJ6ABSYK94P0UopzVpCskMsbzLzBI9+dt59dKGyngPAfqq7WY
7tSR5KTZsZqu3amkMEjJ5Y2ML+fV+Mn+QOKmZoMeh5mNqyOT0cawkVfEe0mlgbFw
98o/rVZm3dLI/5EaN4Pk2V+dUYFwKKr3FpoV6DLjxqrfFTBG3eFa/IuymJh3CqiY
V8V0rA4k5ezwcGOlLdfF6RWRQQd7Is7048jMp6Kn0jx1+6DQRcJvObq0DzTgKepO
AB+W1a1srTnTfCg6HnnO1QZJ9qePoD18L9d5GENJ8yuOXF1ASOjP+/fPBzxv9txd
edhedfW0vzmrVvvtaB8qQ1PMKHHQpKGRcsPj4/h1nThdoWf6kGSRQ0ORPB8FiKkr
giGqT8qp3hQRJpNIMVfUTzxTPZu5bLy+Xx8trXkObMMRPwsEYfIhw7Rf39PPpxH4
+ACsjtgagI7/lhUWb3dbt75fkhnVbajdrfr7LFvkjYRxFtNe7ybPz14ZqAi/i07V
SybtFvUYHElug39cTxGZU1UocKpVn6dHrAt/34NF/xhJpVtyII8G1yr1JEtnKDOB
g2mfE1csHNdWogx3csqGV/c/FVZkzt5x/q26ef/AfLnfMcC+XOSf+WQSNDRcGXFT
BSpAhnz1k0Yg6rpfqog4Hi4hhUsa8LE1f8XD5bENcpM1IJhA0bu9QsNb5oziTRSz
yXs8X5VHUeC+vNUfzgyutY3EsFrQoTVw8byLRUFIEd4baNnJWWc2/m1FcxCFtVPo
kmWg1U+f0P2urXPuOfTedstuU2epMZdtWSrtqnfmsiaUbgrP44qkLCW1Og7IXAwc
YFLWgAcURbsM4wuF0r8cP8G/RGxJNz/Q4g7KMsSE9JgXp39/eyOVcplZvuQoJ/wS
CLzPw129OawSSzQhGCUkz5p5k8X4EY3l9zy7/SnolSIYp5UescGZnxSRkCwI1K0u
BC+igjzGZl2nzKZ5VeMUEWp6+kbQUZdfepm8hOzEPQ7ijxCu/fv2QuKVCBUi2+Qb
ntlTeueg4NksJE1uDMmIG9LLk3/ixATql3kpM1seCEidNi1l0chz4OfXy0GoEr+t
m+ok2d5oRFb488FitmNJRylZIZK6HqhGzgvmFrmiZ1N1TACJWLwqcP6reYs0RD1M
fFZOjsg8B975E5cDw1iNDY4wTfhxcCDuy8pcKAxNp7qjkzznwIh24tgTK+HHoCj7
kL7JIgFAhBllFLNleOceVOLhbzckUrqQieFhLUJKL8UslDIrwIfSVsq9FjFDE2Jl
WHPYq30oSD+oG3EOUfgpufFRjKWQC8YPP8PECz2pkLJFG4ga/hqZ/i3wO+Ewwqo2
h2MsJA0zz/kaUUYORJt9GsuWf72Y7F3PPPtAMXUr/Isv3mkJJ6lnXFpraFZ4kWjP
mN811rOHmGdgewarZUiJ5yOxo9vTUSL4WQhXl0JI5amXM1KrI8tM9oM408J45tza
tW18qDOfGJTWz6k38EyBn97xS7aptPGSXAAxpmEQ0RAcLJplPSGAYFeRvFF6khky
wDHwj2Yo0r4MqbGBOsA3YnDLZxIOSsZqDIVVXzJT1vdbXbwlGxlPVkFzY2kbtJBj
5C9/bEhvoz2BzCZsxZ8wCYntVFFk8rBncUFPhuyCv4iYAmlB4I/5HsHv8/sXTKb3
8WGJZVGeTNrqXQF82RpscoPS4RcYK0qHKTdbpSW8syB/BKixTIXSyOHogEqFv3BI
pJoOzUJAaIHHdxPcpKOZIzUQG0zmQVdJfGqHR116QlXzwJ5jZR1DNVzldin+edYA
3rdjLvJEp23bO8ptAWxqNTMO+Ank78oEA/s9RFcKsA7CymyeLD8hYYE29M0FBgTw
pZvWQLs1WjdGclTLDby7QhLoiMQBUD/1GyY0/TE2fuoUsaWJB0te8BwOieNAa4pQ
RfIbQSO8JYXdo6L5PjsnbdmSH+bpM/GugRnViy4r5dv3p4czyC7ddOYiaa7EIixi
VLQzAzpR8sIEMXPR6/GpNeJub/idJ81phnlDhKroD3cx/YUH+LXAtCZI6X42o7AM
f5QFwCzmRO8voTioHEaZWwxk7yPpHBJ3SMlmyxxJmrXf0Is1Vx2cIblMfXu6FlzK
NfcO5kmmSyxlQVsJDqonWo2KH2IpDGpuWrGlLMLRjbwYOIofUvKBDvCol66jKrCh
xNjcp8XKnhlkr+/fhkir6yKFCb174CyYkOBtA7B0kwMQcv48vOfanRkOTaUbQWFl
wliGTeC0jTV+yxGJT6VXbN9NOMv6mgZx491v0qlZF+acOHojvMwFy2phfEwbx8Em
Hs4X0FyufGeTnt8VmBA7Ts4omsW+yYnCoLI7wWjy9AmRcKSriH0Y2O8gDS5aSNqK
dl/XiLpvCPEn/EVEr3ZiXW2eN4fYUo9FlA+jiiBpODiblOYcXrzWCj/Brc/hd8SN
7BjmVy9IYQFBt+PCqeepMavplWWId2ibSZUdmfip+oH03HITF3vAG0SjvqCQU9E9
jmPpvmelzrk0dytbnJWm9A1J59/HM3LDRFjKPq2zQhOCI1RZ4aJEtUlRf/szh/UY
FC4kVPissdsap8/KrJtumdidrX0p/N26nLgnTRwkeEZRfgAwPYGVzoAPpphevtA9
FA5iSJmqT0nLhN+qaL9K6rFrv7fPdPvihjrsL9jbULL3wi7EXraXBkAcmlJgsRfN
6AnZrF6oEpmj/0hIZ4G7AgIBMPW83GFjnhJWJjFiFp4GGufY1hNPViSsC9K+ksud
GIK2okJvEySLFB95RLQ4Q3XslfUEDjrh9CDZjmoH3i7LXNxvqGqnsWpFV/BoR2Y6
V4v57TTWZERWInzWdMAZVAVhxNM06HoZ4v1RzAGXkl/cQ2k/V7czTv3Krhq70THa
ndU9niiRDUr4w2PYoJX7l7QgCQ1YCk7enKOX0nZkDiLqTdOvsc1yC9LS0ybzq+Xz
DXVBUQUXwdeEe3+lTvdEU4aDh59ylpnXd2mTNi0BIxbrn4NSt2tMuEbgn2MmPlLr
CagcMjpgqmVwF53zyPv1pgErQMbLbErwVJosyD32MIJUTlgxqPZUVlIpKbvR14JQ
Ifb9St4Yj5veoRIcM8MCOxJ6G4dhy6/DDvUTtv7KHG/t/S2RZjgk585JsrpCapYO
TT8HJpuc9YbOqgtUGmJJMSGa3cT8y7ec00qKR5Nd1FH0XyiWjZepZu39fsZExGS2
CatDY2jYouL9sLeE3dQKlb+1junD+DF8Ao9nYyrpGmeTP/VrNQ6yCzkyfsopCKOm
BwP4T4xbRBID84wQGGkktSpCQwZgANvDxxuitPyk7a7/CfCrv2rMprP3Mn2c3pYa
RhE5bMqOM/5Zhw/B2oz17KgBq2C9lFv6n1a4ZTOu9TBrXSJ/RwSZ3MC1wRCRg75z
FfauNZTUjZkcUGC/ixga12L5CQoB6Dkqw1AMlCI8kX6vNYNW73rzV1I9ispZtYgT
C6ec5MOq2XmQosxljQbpimvV2YRp7Y4Z4BjOZPS+KvHjF+v1xl7KY40i8WLAU8lI
CVIhmTljbG+sDq2nH8nCgM3gwvglRTCMNgNvw7zW/+BcaVn6E+rigezaWWv9yv/S
N+RfP+LOy12drRS6iBaOWG4G6AZ6EfGc9m5dCPUcB97RuXepMKAh6UghEYMFMcWk
MN3mOvjtSethFVZD5YYTMh2CFrp92ywQPEn9W28XjYF3bQ2Ep2A9MQTjfFki6nBK
uaTnzC2H1EjpuD0sKWbIkOa3L0BtvpKCrJRyCH6BvWcXLlf8BJmIbRPKUAvrHmkD
HPPzb9jLUrjjFRK8QoYZ3jRTBqTQqw5xsO7XMzjohvBw06gyFsq2zEpQa67nh2Cs
E/ROYiclMqufKH1VPcVW0hRXE4ClPr4ezyY0A00QG7uf22Pb8kqdxkGvClMRzvZF
Gk9RdEEBUecAAbH8/r3164EvCXl3g6KlQCozuXEX+l2wdB4LINpthUziPPDb4a8y
/zcA4Q+X0xKbw8CiJsvntzQyW5g9c0oterTycxp5rjZUXLSRXo7uZXuxVf5fZBxz
0JzlagYkHVQJ8OssfPreeGiU5NVC960CCoj64Bd2y2FrdDyKwxQPuzs36BuqZUDo
FyOflB0Bwi24kw+KSE5YxvBbg9tLpLBRczk8oT7Lx0heA12N93sQXHTWatULt38X
Aq2i+zXgivUI/PBFEmbIcz0iauevmgvJq7Ifd10FIpPDMAkt0a4LW71Kr/mnT5Ve
X6MYzaSv331zkhYW/5dxRYYQqxt2swtE7kGiVn0N0lHZlo7H35POxPyszAJxjmId
k+//AwVNU8Qb2Ql8txj4EAoae6T1M6wxLRlWazDVkPsESxlXdhYrSyEVcAIUF3R6
OSpafJXxMEc2XqYve2xjnbK9+KrI96/oGyG7dKXssNP71TlUwisI6NF9MAfzxb7q
VYV73A2TiqKI4Cs0FnO2YZBxO1IdJ56GtTcVhgj0AVz7XjxKAH2SoGNhnfM3TMDG
2FSOOB9lPDhnxd0K5YI5ntvdr93NvkkqyUXjlCSY7fixqzxoTyAbb7zpf1Hl5BB6
Yx61Q+gLfuUbFLJCCjg+XSjl3gRq509YbjoP3qYItGqSkd4x5Ys4jN1HAjMai39R
W+a0+5NwNvlJcEU6ibv28WuJxiPzulUZQn/46dxdK5wE+xWucr1i4a5QVUX3Z9GP
FA09flsp/f9Y82f7vA0hUPgwX1RQMb5FW6HJlsevHtb8FHmSUs3K4wTx1ZTOV9vQ
rZqUxzzUlnbGz9JXxqWgd6EmK1O16/KQGR6H5F5jjsjmpgqjfx64MSdKl9Fy4hdH
QDb5Oyo+d1TOxmLKq99wPnCqbjqAso64M4Cv8KalafxXjs0aajCjEXflSnkkCjUi
libWbZBk8I03cz8lUxoDtPg/2PyfdO4l+zCmy4j8fRarCCbMKhKLOW7RaXyRhQzp
82+h7p7qtqwyI2KBIdzp97785qGNjfzZLBLZi64vmtM9TKe3gzbnsxzPB/A51sFU
nkgjGR87C/1QnwNOND5uSpo7kgHgAGLxmcLfIWIsYHnShjep9nevuhylCZfy9UYk
YP2K7SdJ5m2/ITq/8uY/Fp8fejIcH9zcTUyrbsWRTLmIb7yM2kJbL1uUGtR41Uct
ad3DRPBKgRgCm19ob1tdHaS52+1PJ9IXVI8SH8Sd6aimpaHwux53gQE7LykozDQ4
28351l2DZIqRa6/BUu1Z7FzcjMCYkqutsIwXomlYflo+MIgNAqhu6ZD95Rrz3rf/
qaa+5dVJSOVfolEyCOgo1qkXRPrVwnkC+GmEB7o4l357EeIfwHXH8YlnO/KgE1qW
2fGR8HZCkFofxxjJS/O8ph0vfb9HPG56OZOjPoR5obBPDC8blcn/tVuFzUgYrWYo
qhxOd5p66j4TTnGk0ZAH8HnnQPgA5WGHe4npWGk91t2OdclhAMvphByBQFVaRASv
m/eODmv9fRzF+jp6Lu1locYR6LlZw47mqq3W5HpH332qgdEiVn38+kcNza0qPKYg
1UgCGASmB/sQFVrtFGiFeSo50/pthBppkbEcq1g35ZP64gB8cNOCqQFndAGlbiQJ
2boG2jX56sa3mK62LgUOXrDNVUxbIUxOnBlZBTb0+QCsSo1NVDP+4BhG0A+/+Nlp
7Edx3GdCpQKrzs5l7s+greQ2/gt6+qxtX9V9jyQzACJli0Hg4q23VBZ+dPcJZRqy
KjxarjJ3/rXKaFK4F1svxhZNiHGGqJCCwoMzY2iyqn5Navt07MKh9rKR4biDZaMc
v4hDDJdLv1m8xqp7O19WlOdIH3qVLAR6pMIFGp6V6QusCyxvp6My1vvaKB5EudT9
Vemx1x2U19KbbQwfmH0n1l6ZjPzBhldRDjyeTzTGolSn/fpYXHZWKH6kuKQcbdjU
icuZAImfwXGxjsWU0puJKGKiQ8+yjwTg7yykiVABI3gm/djTb28EcGUpY1wK9MdJ
y527sNXOVqr5PldBrkLo4sC992KY94KG+BgIeRWmrZXPfMD8UqtGP+sHjoLRyORI
OlxvWJByt0nLq35hKcz36/lo4Xt1l/DUTLJc7/4XA73FQjUHd5M5IL75gnbelrwF
SpJr1JIWztAQ2TC2qDvnsCfyPVeOvsf/iNUadEyFP3IhelKe1ebmCsvJ70AEjCw4
qP7jvT49C03jaZdQHulN2aZT3c+KCJ+sZA53pscUyzyhE8WEBW0As2Y9ZW8CN2hQ
6OXH5lDAL06g+yGV5F54AwOsG/7W9p1jgN2l2s6cCJwQjLVO3OV3jhrnQFK78XF1
BdsnZvFVLJQXbE0w9hkzNiQwRDKHs2vBRYZJD0KP8pml6PYnCDzuYjZZaaq5LEo2
zWrdszKqICuFXKWPIHLOFPodWwAxrUlEZSO8g1Ic6PA9PaaHEurFiQ8YD+fpNgZ0
hbOEo3ax8bpJupav0wC/t6CF5q1NDPUrlUVrwoCgkiHkp6fFw0L4Qx7eg7S3KqWt
dtIfQadQd+KQX/Ur57HBkMaftX4UDfOwBHYvO/h5gDwxNLhSzo0V1QDx16rLi2XF
v1XwBdt6kpO2UexSj+Zm4aEPZEmhpn/b/Go9N3nva8My/QYNIao048e27siheXdK
ISypBB3iu3WcaI8mHQRZEZeNHwv6mrIbzaipTCnLy+4mt6RfGuX+Ws3GRjxjM42A
lsWq4ypfm27TCmwOzfAtT9VYy0AYP6lIFb5nmJsDz/pjJ8HS0s5jfczsAY3UQnJ9
iWtQVWf+eAPeQMKS/SjojOf7VDiJegTuYNcuRN8mKF1+sjotuAvy8A8Obqs0CVqO
`pragma protect end_protected
