// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:43 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N4p83RJkjJvAq6u2jyBv5EELsFIkNvoyDh4jpItrXqB7chjuw5YTbPqsZHKAfWDO
EFjNKj8o6krTtStytRnceApUGONdz/hGuJQcNWC7AxHWQ1ssOJE4P74eqRxQSq2l
02ytuTxoitLBNhgS5xgPh9YaUYjx2yITCebQDUhOHjA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15600)
rxX2TPJT6JYNWv1f2/jfYoncWndXUxI7a8X8JaDpQRa+7lTwLu8bj54GqugIgX7v
u+49SIj/qBLdsPCnq4rzK/tXIlOsDbZ+J43tmNV3Db9fSdVLEomJZwg1MzACaL9a
r4R/GraJz3tpAkYDD3weBe3GsumcvKET6oG5dTFxn4Vd60VDsHgz99OUWyUGWr0E
dawy/31PsWU1+rkRo4pM33f1DzSrWQreo655djuDZSvA4K6LOwNG1fM89Dsq8/PE
cq3zxIoQGUVk3bmYFXAKgxJjrjft1Es4VmwvexHtvVPDbise83KmqbgJbi6kArXA
mY4rk5iEXHtwz6CqA39CGz1NSV8TiV/khmS02gyuIO1vkPEgpu9OHK00RUoQvEXy
5vECdY2LQ8cNJvzrnCQyEcXNgc95z64ODR1kG2UczM9Ep87ZUZ8TbKsjOmILSiPf
XAO7pXkQo51sCkgs/Tsuc+107ndaKMULn3oqZIHmIn7odg9Vfa6lRPr16kY72TCn
aFoCpunKh/YW5iNK1ap5fPTpd76YKvwaAD61PbmimMtfcZgyJ8Gx2O7fuTuCKVVO
xJTs0d4w0GUhNwhIsnE4iEM7Kj/Nm6I+DgcXJb924tPrP0EzIPKvEzEaDWOv71KR
h+gga0W/SVBA0EBw6QxEKLKTtAjkVG/CN2ii6PlwDx8a7myKIJoLbHD94wV3yGWa
ppHhxNRYu3ukdi3bY0VyY7sjIUErKJVpZKJvBxaIElydeU4vKHCaA2jvyLhS1vsm
e3ZZ1CQDs295BQSCHr2nCbvCWf/zD2dqF6amWUpufULOQ/Bjtq374hUvOGtlTtJB
CeqCkrv7Y7CGh6V1QbWrVt3VAtCTruagD4kJBPvGCQgTKV5D7OgZAF50UoZmsxIh
b4y8W18hgKeXFHXE+xvByICLDs+YY0L5TfahB8gWKKzjKKAB7e15Ujzt6fKB4yoN
5Z6M/PMrXBSMx6STMVc+sDx1E3YIdg9HLDwvtXGVchwzEym9QrR5NiZTrgfMEc0o
jOiA6CE3GQLgdmV3NmTn2rpXI5iiEgC2SCJg+f+wkV0ZJgdr/qhLrEOm0HBKyhGJ
ybQsPLD4VqUuibh5n+NYbq8rovuZeZKaCRuqRbwqpCGbwNFLD186Hcxi9mabBfqw
uW4BUB+RxhWI6h06pzJjgtRNqlTWtpoapiF73lzAHvUld2+rdmmbXVFlcYnZyGzz
5NW0DsKv04L/HBi542lP6OP2HhLoNjovLPAJWXqtF0yS6/OKanjO8FEsOSAu7Wa3
QyeeI0/DkcdyNVu96akSmvaKMHDIPoCQNEgznuKp3fOggNePcyy9BbQWhQeXJAta
6rI4M7KpFJ/nw+yB8uuno076tF9gEwZXeqVRq+BWnItLizTZy7OXdkhWznUk8sqN
WtakdDGXgION/CfsqU/r5SGPNUw+o8TBN5UBxfaJsBqlCggIxlbl2BkqfjuFzLeK
/0CEuj/mC6lOLg0omJBMScmhPytOjopTc/KMPsS4VN/Uz6F+cmY28g1ZGxHc/XCx
O1lK6byRxPJ/mTQwl4tyNh4rDsa88RlU9qKydPzMiSHYRa89bt6dGtr6ECQmTCSp
UkIAU3Cif8kLuIIp9j/LuPyjK6JHkFGXaLdtiixX5shgL6ETg1LhcOKeefZjlT5A
2JPDY/Iy3KHzWcXp3UlxjhO8W+COWW240Rbjl3QLFnXLkqRENM6PtjucIPVq53vp
XOkMUF/buIYLMeFmMWI2IDIlHVhjrC1uEE+k4OPz2uJv5n3/MOcTI7Q2JdO40B/3
Ddcp55BAGsuGHYRxIKeTf72tsO9h+BbG2y40+ohozOMv72zAtngZ+yoHkQMOo+5Y
R85KyHOjHfE2o+NdYQD12VwK6M03pa57okDt3oB2R/Qr0sjDaxt7YQUEBe6W+U2j
EyaQ4Hin3ZDfqAg/9Iom5VDnz4Q+ec4UlQyDWXeiAIPy83tGMMCqSNycqZysrGAQ
MpQsK5xIk6fbRkH8/KDRs8fT4X6HVcLUJtCI0YTj0Nu4M34KtKBvPlN/WMw9oRiz
BBUTh3vL/nX84PJcIuaJZAEp1wEcIC5HOrnuvGsURBG+s0fRD+FOeUwNDc8pagAE
m8E11l9RL5DEhrfNCJLI4WstKeZ2JRt+y9+5Ro7VT0ypzTefvY4K0+ES27mN0mha
7tCQ+GHC/p6YKIE+SB/j1hQuzHEtngcV5HwDR+CqGMQqg5ni3F2suDIxLXEfvQrB
2Q5y4tUjBMg2spPQWrJvrn6cuceE91Y6SB8BdvZSh4zjIzRZxwwjGLJKRDZpVxVR
bnfA3+KgzU7Cgc8pdXATek7g1YijeVIbYpNFNY83t+ywCztcLvgO1cHZqWgKUSsZ
9RiyJwGwKOT76wrVEGdLEno8Ns8Mw5ZuAt6+DviUYq9xcMdBGzgPdJURQNFxu+Dd
ACjYW2L+PXjt7t67MN2b5dX9bP4+c1eGhUi8nR9+v1c/aHZ7v4CsvMSExNCjWqsl
wxshYzpJs1PwQtl0ndCTrqLzY1Rc1Wmm3Db1/zSe27ijIX39sUhwiAEbbdLXlmNe
99k2Irctn8LYHb3uaAmQWAkeGnYzp+YlWoStpHOrK39G1Kk18cAc2gM4GbsFtDxs
JQrFNJuAUvfZuQnY7ra2uJpGr3T28BRyAmid30p58tw4toYnppZjZZEdjnHX0F/P
ynkEiCMnql7hDG5xtxiE2d5dEQA9Q/rkTMNdtOH2d9ig1ksBu2fasT0OQ9LEmreA
a6Wn1/hIS/1X3w7rB41J5HcCOisWbfG788cvFJh4ubhIW/H9jxnvKZVrr6+xvuWO
+Rqvnj1IVn++jH27YOB7TmuB7ssaFDnUeJPSLDJ0y4QoPgi30do++1bo/uYQu26S
Oo7sKRSpRZGQLDwqoYbm+KLAWB/Sqf3YEO2AKyXQtnkyQjyiHc93sJWENnj9DbM5
DdKYAwU621pDcwePQmmQFf+iTD+UrtqDiFOOPmZDxUlOjvxwxshESHAnXfC5Gcw/
zvnisx8bx4ZBLzmWHCAG/oLn9Duao7Lo43E3dWszdstXzds75LedmLxDr3xH5f7T
wBWzEIf4Uqfv0rJLL+K7qUsZ3r5gO/X8WI+VUsrR0wSyniguVIhROFP/2suh8WYA
xCI8S3fufIkaivPXiLHWw+jSHA2V5q3Q5bCn2ZMnePiEMkk27xiddQaAfzDxViUs
1G1FFL6Ljj9XNTEX7x6RmszwOWV7qlBpvkuIB8UCPtwLuGpEriD6oVvCjeXXH1Ap
AIOM9JAgTp24NW9prFIoZHtZcFAUFN+W0K7aowLF0t+RE9OJPoQaOfJ0bOTfZcGl
VL2Ssy83oT/mN3d5VvL3UufNe6xH5D0vnXKbSOvRplDgbi7p0xLzbgbxYMrhD0Be
69uTlQfaMQt2TJ0dDceoWXE+FPZX4v7If78HwbIjd2UpdGgOiMZ4IZ57jda094x4
0l5/iIUusKnY+DwhGx1RQZ05IUGvCMdVZGPp0o9HMb4ThMIjaaSg7QT3oQbJvXkx
+36bbuZyr9eGPv9S4h2xhgRHqRZjUlmFx/w/fJltkjtGYKvW5R2JX291AlIrrco/
YDe//0eSpRD5EXzbe96OUSJsUmntOzYJxfT7bhJhsptu2+blb2yMldeSo8zl1yml
RASMFZ3cZOwdEftAAIqKd8Sil4Hs+ovSm99cQvPaX5h54/NFAOxUNZDnItK5X2se
8rFexRbflzurHBU/M5nK39Pn1YYNe3X4IMp5XD1hJmsqyHS5cTMX92m9EppSFQUR
evwntjP2qcSBKFru8Smvk0wjzPFpzrjlYeLm8SkBTDYOOhbRzBJ8EwxBV+BdEVEi
pFOox95feZbdhUSX9x4Qo5Bxe6lXQmu15uZ505IlWj+AfwJs0qJ0xkoo3f+uq7jc
jRGWU9hAIguyAbG6f215d3YU91LmfBxXZJxgzgTJHRQhUQSwJBzPwbb/WfQG5W2k
ckDGkEahqCHsQvOf5/dOosnuFp0ikGlLON0vEaevj3gGZokI5wNX1WUAGCbu2K2y
RiuAHsDPFhF933gPHZZbk+MD8Bq0yAG1oTx0+cWiarsuuVC0PXMthRxLpaBWMAYt
a+mG9AxOXti6AE9sphZ6duuQ08W83xiXUgPCNcWL3lhnySxmELevduNU5mCQN5Rn
4DBP0PTmCtUeQYW88vrXuwNJvPHgv6Imvn/iJrl9M0a80ZLN2Ka6Y2Hj2q4wJBr6
ocZyGM5wnJMH2aRDDXx5ugcbifAJA25AA8S8g+6U5OvozOfZCNfhykO2Dm59CX0R
8zBSQJcMaG6TYzuMuw09iRRxp55t1dhc5BsWrJPQSzcIc/FhOwkbc+Ewiygqtgjk
68kr1FvgUgjxyqivru9pIr4BNWNKZFM7mSHTnM98qIk9ZxUuFjoJ8Ge9+emDmgP8
EAUDDrihM0hlb5XXThM41kQhtXbXqIZhDCXvQjMjz8UrFasp/0u93nUSlQEolsRu
vJ9pUutTjCqPFffYzcEV+nqoBh+7FdRos6aUqF7ZQWAvk1LRucVwBTa0hCPIh8Cm
bu/6sB3g6UiFJeR+oHIFKd3Svz6GuFu6CwkTg4g5dNSOsYeCCrvYRPcUK/PxTa4r
2GzPauygxZiivWI164aCzhJBeV1ng98ZVrzt+RykHh6xFGBt7+nJ69nu+Ahugb1b
FhtT0FCm3UYX0+Y9Cri86jEjMiCQu1HWM6mYaOgFY0+QgiLRzd/m+i3yF4U/w3Ia
WFT4JdchCWU4LCJLk4yQVc7JLrtvFL7m/HKk8MtttmDG9PZQtNEBlx1xc7GyjFU1
FM46ciiAHyIZbCHxUcc/4PN9OiO1HCa9alA24QJ8bPt3clqo9ufkYhWdURWwGxXP
GflmRUpWuD9DJbgXQL1nxHd+wvV2vmWIIESLW/WJIUPFHGVz0BODOFvOZ+3rm+qa
a03hZISnd158Vo+p+6fYlJcfCgg55TuOrCfFdpWUOHr4nhSWhRaXkfpuN13+DBcK
j9km4xbz6C8shBnBdE+dYcEjofNXDysjZX9kKOSZLMg+7dh202RTu+MJxPiBJuMk
AdDoyXPiRtVhSDnSoO08iBPVt58Jk50FgTRUaqypL+/qpqr6XHylD4PRbjMNiB3C
X3pr4cpAUvbohl6mP0XV/ZvtUDssFyCPyeyoRBnu0U7s2+QszFhFJoK+Jot++RiU
c6ZDwvoKEyiT3r49GnpEgtAfrAiUNXc/qA3SWYQ+S81N1Q72W6Mrf00Ifqosc9l5
uQUOwBNKHht+8ThDrVAG/5HKxcuZCBwevxBNUfH7oYy65nSA8Cw5WLNbNuf6AsjE
7utWZisKUPgZrzUuy9Vosc+J4OvUBnTH54XeII3T/PNokDtLRdQBrI21Xlst1wWz
V75aSOIXVI9OHZoEzZHOuGMEbDPiuy+o3Yompii6NE24Cayx+fCCUOqcI/18HiDi
w2VmI3yAou0Jed04bBt4jVdl+8dW2bbwuusA7cI9yrPk06UrMlgv8H5G+d1FvPav
BgrlcuUul/0CfhuWZpdT7xOI5Y/nJZt5ctkNaPjJYH3dO7LbI3MnNqGmmFaAwZDM
eAWp4vTKvNH2c2rRjnP+WP5BswsA+EDGaLbUEo5ofc3GD7919sRpmU164qql4zGN
4Fzw8BNUHhbec20qzaz6To7NBILiOB3YA93Us6Wd9aOzNnKpoJsUsmR2thuqztvF
mCjUROmOOCwQRdr3cIycXzymlsQrJ4cECTeuOyWpTX0jrQ+BZV03lGDbtXLkEi0D
3eqkj8noTS1amAGMtBLo/ozfui24CVLZASYozBSAmHiimF3SNygUfyLFTP5CsIft
58UjiPiSXIDniqLfu7/1uH7UXzj2HuPJeU8akL2OF8D3ABAHAatE52WSMxKz7s93
Vb2rJbwnfK1jiYyckqrFzJB/RrGlVsWfSLfNiISMJzc0X9feBg/XEPR5WT8sMTYL
Nm8hFC49L7yJgY/ZiRqJab7jaBqPwODWM7ghK+QqdONSlezY6ZA0b3t4Rcg3+N6v
agJZp9bfvUyBj7Ca8EM+rQYP6HSrRopfWTvwW7t7NN0SOfZe1Ju/v8mF4IyxBtuN
diz6E+0mws5cKOZIoO3xGl6YhMy5ZMbmxkVTECXNYwBg4xFC5YEKQxpObyBZZK+O
NTjmfpl1BTC4nonpTNHViI99X4kp9S+1I8yDX8XhcXPsAzwOeg0uwFqMAP/PEgLE
F8m6PbZS1BhHmmkR/ivjduiG/tfKKv3CcAG/v06mVDC4vyq4bWjcJPYi8lypJ68N
hBZGmnoF8+56W5Kswlki45qfLtWBQ8BZ1Ivi1ihu6eGN0CZEdfKVgIQwJWFo44DV
fRelyz7GmZXjgr2W/1XAXNxsxZ/UOic2MWNI4M6IIuw8aBVzdeHL012h9DGskz1h
U2/tmpKOBd9rJywRurvp2A+fdooWQDkCUR7OV7tbPbhgJSX8cTxOltsOlEzzKinp
+BjhHCDsMw8L6U2yC4rx2izd+6shLjcU5UYXfZikgCGTIVOWpQA+mCBFC1NCrfeV
tiGZsEcMlSDSpe9rIZ2JAW9zu85XkFP2/RN5tZ8catGHBhSKEmkyBRdkaMy4yO2p
QtCxzp3bhFcAAAhLqZZ7G2DtxFiBh8nf74wgdPjOQCCuRtgW4I/U9Is4cg8nIXHP
LWEXIlSrHBIoZpsiB5Py8P/GcgLn/8itKtmnwUIoswHfVRD8/q03jP9uQ3ooWEcx
UqHx42DMRBGYf0PEcCMqBYEw2O3Yynp+5EP9HCYbAWNOlR7jW/yRyQVCnEJRiN4F
Xga+DaEs3qEl95t6GcWS4at4onzy6qlcz7jAouMoaaDQBCnRuM9R/S+PgGS08XqP
vu80i0L0AU/S5rAFiMwaS9kS8XbRI7fyEBWxfDiq5wFe0zqWr7rQ1nItqjE9D5Iu
K3l2Ekp+zwlDGO+NaimT50k5+79bB2wLF/EltYv7kaZaVGjlBf7e3bJ+ctEll7wK
/TKOK9sBZhxJhcgiL+4AQkp886kuv/BCnqQAXXHFHfQy4Z059AyCCxRKSiPexUuV
asi56V8DmsgwAssx+waHfy4ol5BlDDMWriPQ1AWqAex6jPl7GQVLPXiOj/EaUtRa
3OahoERO0+3n1eJiGyHza2tCWuzIqgrJMQL3KRcz8SwNatOidebMf+bJQNzlW6AO
eCoOfk/KjcxEt1Y/EZmu/wlN/yGwisDujs40V5jst1/Y4z/+ozEXSefJMshj83eJ
BPtRNVApfsEBic6S8aPWLxEoWkfGExgtytlp2hT5Ws+ZQGpM3wJfwmr01OmHLA8A
yjbIKmB9HgKgSHS7dQuZ5fa+ejVrICPp59TLkXaJzRqzKsJwb//MxE/8HWpJ/7ac
7AaUKGwsNYGD5+caTO/Uv46J/Oo+FNYYYi/czPzLQACO3b8dcT+F/qlXCGwa/z6Q
hkxxdwaUG503LFE3ud/ENGqrguyMsyExjJvB9GnUPlA4oc6MIcPnq68zvdz8rj7O
RFotq7C9q1eMGTt/E+zAyQzRXvz1fwAu8U3gJlUPQEyb94UR/G8nKqOt9VJG35hd
/16OhQFAQcamUOVgjfwrbv/WarK/bQnKhoS8naVYlAgBeT/HpuldZYE0piygvkLn
VVHefv52s8LWS/C4Sp0w1vz86yB+VOM1nkU/9KfjkQkiJS0ZYfy5FWQMfST+y8Re
QhX/8A9Rks/IQYT7DS6F13z7sUmEb3N7pP+oexJozeCKKYOiKCGxEcaGFmHnipUN
L2nX18joE2on81bpIBtC0qY8jU+CQjufb5yiEj66QdyBq+R45O2nlzWKAkALULnw
/n2mp7qDOvh1DtQwUtne5q5AirON3SVr5Mh9bthUzDThrQ9FTUlz0MUbxtuJlFUj
8dhvoWgepnlf+l84T7a3YiaWCCN1yx3LcHTzNRQrpbPWxUQQTmARWixrXFuwfHXW
hE2vQZZCnnvob+t3QDZfx27duxHhtJddsYEs3gOSxf/ZAeU24hXfce7x4KfsFUhD
S9VYYe05nDPDKmS9gEcsfPuA1YCtzUJ0a63ssCjWlEOnejSkwIwCP+BXtU0QQMRC
YV3Or30UBHj4ngFfcEJYAQFN+YDgYwIaKXYcyLNFD/q3HFfjcXlYfwMHHo9UuCO0
Yl8Zt+VRNqyIw6pk9mPy1oifsky44cl/j/y6k1y5l5tEzTrXXX+5yFvZEwWB/I1G
R/dYsdrbAFjlt88sN6/N9a2z9QHih4Ti4yiU0kS+nZ1892KbXqrhUD0NyJZk8ioM
tV7IOkKgXbEh0O/q7QNIoOhf9/tdzWanEnA3bwplIMam2HeRxoodbzBBUNaHw66k
1D9sysJ/V/3CBWox2M0lC53Yg3Bj1mnzXJOamHhEs8cQH1ymfy1kXwRKSwJsrzlF
s+kssRmn6qLsuB1n9tA3qSHp7va3UMyrhtK9EoE62+SKsGk5w5j8qpQaopSA9DhO
Mhm/SVRDWKvQNO0TPxj+N9tmftxu6Eel/9zbsdZXHFJ6DuqmmHi46j0mUZg6ayi7
EZMLoCVv8HjdtKwzKBwm3v0wttRZNPwFe5m5YTwx1BlS1CI8qtXa72NOiHV36KK7
tP9S2siU2ZSysafF0XgWf5+/6eOtdhSEOEFeECiw0Vyd//fmDRzBrobGOr/dsgqZ
ifWdIPAMvIKZGBtYCJfRl8XlCr9HkesPaHzV5qc8L4cVTeSeqHQ9yb2nKUquDEKM
qhnqYzgUNLVKS3w4ZuJC4tZBjci/EVPYQdO3UDvs/8o7ZmRY/Ad2vJw8S7qBZ/8L
pw65JmoMvEyQNLNgFTo1bwSCCd0Hu70bF8ElDJy5iEkFE9CjS2dVMQUJeP/1ZNfd
DEevqBVwikG7l5Ekysu9vj8dAPOMmIC5dtahYynN1rvzlW20QAuLeZY6GeeL+8Ez
O8MtBIBTB9TFVDEZQPvkYKZNOtwTiFFi6FzKkv11XuQFo6gKDmW7BGPjrGfcqCAp
jWucVF+ExiH83++Zp/A4fgauzH6oUDHWN86/HYivfK8msb4ojWPnn4ucITK03YQp
x/hQZif0MDEv0+WBGqmXvX37g9h7hBZGN1VEb3vIE6Aig8UBB8SGtNL5WbEr4uVH
KXNkQa6Q1nobdMn4de29bRtJ7Hz0KIJwY7nbdBeU35nzFlnZ9s2OIe3cO6qmYSo4
3Q6N97mvHIyfCGzJlcWXxd2uNMFryACTwKWhOcu7WlpK356WogTwzex8+ZhbEBlU
axZT+k8jbsxFEgLfN6TJDuFRkMJWc/XYCXqNPnly4JHSiTOLCzJHu6tRDslCaU1h
ticuwBnYPkTFsMk3vS79wzjhcnPSpX+NJF28kkGl/mqrhX93T+WbomIc185GawaF
CF9U/2TQvyzeyx8rscfSJUEBP5Scjs919nKIhYLEbB/owvZI/Sa7Yh9iMip5hc2D
BCRON+tuZztwQ1MDCYvqiIB5CjxGEdTSdrhy+lpW13ZOMW45oHujwR37HnM99BPH
fhcO3Aut32lqvJetiMu3qkqJf2ATmu9h5tPsTgkwPthPmyhGjXHP3eYArUYNAg5W
8/4Dc0QZnC32Mi0m7KHD6KRLPfy5s46E9J+/tOf60jRuclKXey7LuO18PKjczQLl
WGP/1L1KPQLBlj1lzS/1eUOafRDkkaEGFnbDJHwT9cLtrZohucZRwFYugWue1zyj
L49h1OjwLWhgK0GBsRu+3R776rkeguIdWr33/eg5lxNeYpJ+tJtqvcfNhmd9MJyt
Uzz3etKk4o97o9FYswbJTASVfx1wBr9Iu9/sKqy6FBO6KEga6ZuqcVqdtcU7W9RN
+qu2auGFhzIsGSpPyMo2xp/Cni7Ha8UcG6ElNiYy7RLh12sHz2ZnquEMsqn6JFgq
B5h6MOGnRIl50TAlN6eIvFrWQ/ta+2IPbb97FtB6t3B1GgYyzu1/nQRGJjDjJD/8
1hPdQeWQOyRKqmoe/xyM12KhJVsxbBv1WUmp2tYp1rq7rfucsW2LDRc2kF230Nug
go9VplCa35ILlr34QCeZDxuhbavFmBATyiyqGinFAfPvb/G+blu0E8s++ZT3WJv3
hqV+Ot4dX2xlqDjzrDme/06uBcOR7M4ZReAlei8vX9mnuxv2Mxu1dNORKyD6FSY3
OVRx6ZmVejh6NUFtCMJL6HzBgpWfgHt/yiXz5gZfjIHuwFaVOqFdZgTvObsdYjET
hDcnbbZz7ffM5bBAyNV6z6lMVu+K4BhO51X/dYjx46eyX5TftCh9Cp1vUb/0EnkK
ya7+PTm5yQUEfhAoFqOYxZZMm9d7lHXz1gTGaYWqPUQJ9PHknayPCZxc8lQqxsd8
Hk0bi1l3ooy2FJJ1kbOe1uATT8wP6xmRTK6beuED6jmzvXEG8PYcYxklRuN0TrtF
tNa9LjbQ3QFVLANrbaj/vXe1cUT/gBWNnWCuc9GLmfcrzhOuPvkpmHxztz+KCgkb
YbNaqEva2gjkzAiQ/l8xQ6Ki9uPUa+TCFK6uA3g765f0swQdwpDsUJEzbxPp21ZC
qCYA2aMpMi/1/MPsOFcBePN7yoyCGp56oEsOEgHLaU5Z58u3/cnrWIwOveVuv5aN
4zFNGPmytYqNTm0kMFC/ktJsLLnI09ZKBL98m4xkevSV4Y1j+wbW0FlfhtyQa42R
icymrUF8rZ+5LLC4FgVUFmz41GO9eJHW/LP5plHrjpoz+ToKV/+DoQWz/HBDY7mT
OYZj/5+XJL9Q0Og8MleyCJclDghVFrQk6Nv3SypGQZ0Ch1eI9XociOyoBKoBFf8f
BdQslNPjPEM+RgjYaekJsQeNyJDaKZDD6adLFOVYNu9SEDNbRvJVRkqHdBpFa4Nl
AEXXNMz66PamRQ+0BBE3SpmLELRSXVEd0k6Q1IBqL3+6uIjXY8SqDDPMUg9Tekm8
AczzSYH09OGPCkN4J6/gnF0Fs2oUuJaFi3gEc00PS+hJD5DpK5d4d1NGg/IpzFPk
HkFaS1CLiiFCXedaJAuvJ9prksVmoMoEku2MlWzRA1L067wDKDJvggD1yXBy1lU5
WN0usSbMRpxNAVjBBLcGYnRxVyOTXgIRWQWSJ9d9L1ymoUjKyX/ZIh8xRetAFAak
+kcL8oCzyYVdp7I3Ve4vUO93IVkiE9yHk3Ya35Prq7sJr26t8WHo6eBJoCqi4ahR
dZHnbPxYiP71DPPAJhl9NjCmijb0GsMMJcHjsrSZoTAx/srMAXM2WKe8iO+7z+ou
hjdRhKY/8RKsIbCnwz7935XVbJ7AI+0OacTAVerQkFSns4grrBO+2Nj2UeaWC9K8
VJ39HO8Ih4kPUqNwUGcbP5WPzUOQaHGD49y2Yu9wyI7oZHcKua7M+nh1d08ZF3qN
21VMU33oxQhfWsesH91NHOckW2dh1DRxAZ1rhMForsah+IbxNeMYI0Y4278CaMOH
Dkhs2Rw5jB8W3HKQ9vxENN0gU2XLttRwETF1gUCJgpFRchYqiDhJxgcVHBExMG1v
fxAaIC4UFcBx8qaizTP7+avIe3NEdL83XhWydHDOQkvw87lZ9UTgjSQuY5GT8zuw
QAElmgcisHMuYhMkHygfEaSvCP/iAQx+Ag1d6jqvjKJGu0UK22p4pIvj4mNrXVI4
yBI9+rtkmxfk4ioL0C1TdafCX6LDB2QY6y00+5mJnmt+5oBHAJv5KlC83qB3sh38
yixC1QO+QiDZquG7Abm4PTns5M5d6zWra4a0GC7UjBgoiPNqId2OJiA1STpuxjct
N2E5t4Yux7FAJcNE/nBgKV5evmwRXfE28NQk4X1Giu+F4e9oQyeP92MNHf1vFiiM
bvoNYp9ZK0V6I3EwRB7CphNKutBLo33UMqRSo5pbV628OQiRUY0LxR8kEhqz+aXX
Cch+troDoAHVNOjhjsAzefZPBIOJPMPW2aDiQn7rRNWC6JAYXmb76uAq2c/Es1Hx
jA8ItOqLPcMy8xm8t6bw6mZ1pjtxr8xGRsxCftGR/Y+lEISK0YYyT5oWRXXzLvVa
UqzrNXOzCXDaaROuEeyIA3CSgNnojxUZUO8XEnGNpBDxMDRQqLJANat/oWlkjLko
nUDO0j2yq37VJ6+slt0CCi5vPZZnwANbVB4zGhA4LyCQNcp1/JoWmI4JK2ipLDXi
ENdezIWmI9ZbBsH6g+1Yj9Mzeh+xct8QsZ+pyEjM09OVlPjPHySkIcx46gw7rgBR
/frKwAkpd6y/XgZLRZd93MEJyNgniZfSeN10coIDKQ88aN7WL1eYI+zUwbRJ0vUK
W4MBUWzYXT7HvrfFR4kJ/H/78sbVjmvzjHcyA9EfMlW2IoQcXA9IeDhIaEmvARxe
7F3XvCXbJJji1oOKymjKsvQeRWkgc0W5oo/lczZApDpApzhuNaErA0jIrlv7AM9v
gXHCM9PwKmcOZJGX7lITIQaBJpgQBOBp9pHqZAbLBfTVHWfP5XPwfY0PZtqqEtZd
BDVoMj1gXnLeVK4cGrvBKnr3Kgv8z6liyQQ6oQAaYSPxxjnI6v84bS9rWN+aMZeC
Fhv89v9cFASpo5zUwH2mhLjuArCPXv3k2HUzFqnvPPV+mojx1SDhN1W3eamXbSSc
C6dK098QrOe9YMVvM5jRHFdg5SNQkpkriHrNhO+Q+hjZDqBTXXFCrUu/G7f1zYJq
DowNapRxMaf+p4lns8RPPkNCjDBdVgamwRjLnfqEbSPTJiArU2rnZUEOyFNWiyrX
Z+WIMDQFOrYDLwZI7jWJO9G5UJNaxAj7QCXVCTPNfMKQZbaEx/xg/6di2vAZ0w/L
oyWL91Zlas45EsNkVWYh9NwpNhLjM9A3C1P95z+YLML+jwBAPkx/ouHFbeS2SvhZ
slKtWR1Fwn5xbvpi/lN+Uhhtd2f105Tvd3VesBVoAFtUGujCMsg92BRIaPCXaJyg
z2/SoY+ee1RWGQfQ24ne/CYqqfAyc7jw+UmzTCXr/Nfgu5k3jqLVzhAdgUWVFYgq
RGrZU68SHlJkE7ptCkmSQT5gaUrIlahE/JDpJGUMpTVLFxVbWxGY7uEuBOKSiH2v
wUoBGi8Zwi6V6QTB3bD/6rQa6eW/C5Xz7pK8CJdRaocKIXbad/PLlcd0NOtor6eD
iCiQVkCHIDA1yswYCXfJVjQDzM17C9mLKuntReJCWECl4WoKzthwaPMBqrUqGoNz
sVFD9p0kBmT/NUXrs+VGSqs3Cg66ULuZ55jbYd7eMYdzvehPRHzhgHLJRwy4mc3S
MwoYV46npFSzf9u4ANdiTQ5vMMdhZ9iYomQUQuL7FhCQK1Vi4eSefh3p5UEOEnDD
S1eXNmyg+MCfd6G5qZnIcx6Q4EmJC0JHYpm+1JowqJ8pXfSELfb5Vk74B3nB7Yft
2203KY/u0+gpwd9dpvZJ6sT+O+G258utvSZBCsYRmScVP9O/GqWuphqblKtbcNmk
klFX38zxsSWYKiHaO1Ba+DDcs/gJzFOB4u7e70GHOkRpEveGbyrehyfQp31Kt+eC
FiaAQwOl4dcMU4YU4Pa9eIfB67BbdpUAVz5d7Gd4EW7Bg8f2nexh3+NAkJqlqwHR
1ykVERXErkDlLX2/3U5n8Zl8uzdBdx+l2ofe305ebuu9P8mMhhzVP6RVW2aCZmJP
LXqbI7ep8C7BtxaIKkSji/zCT6J9drEA0QXqlDdgmiP94xOlhv0szFEDyxf6mst5
IxhuFLXdwUHVn5rdLoYn+zDGGESUwVzgwCPupfyqJ3KlwUJ38gFNNmzG/F42Es9q
4rrZcsjgLxEk+hUxpLEVh1Sau7bGMbAVfR6rlQqic6oX+uuRfAWVpa6BXTT0JNyV
tnTdVbVJL8D08AFd3feQ+QoXHf6CV52YD6yD22AYeoWFE45cAVfG/ANqMFgpAsCk
vyOtd/Kz4cEd0In/JeGDohoiO+9aAZHtXL/PUf49QbebNFQRetSGUK70OeLEsmCc
Y2X63XsbgN2x5ibpliWaG2+r3UoifrnGDcukVuSfMKPL6QPvEJOWKhLggPuv94gI
TEQ3AKv4VUrAinVtqi1mXEiebpnGtPSynO2SVoYRW8W80xW4LylR3Z6GX++lbFeH
5fxOn58YWBlE1orEK4J+GqowrdMV4C6+jXc7VhjLs1AXh74m/MPTKhioAJBSJ9rO
P/WQ9MnfzKiaBbskD5yPqxhtgDef9+1iwf/+D9TBmXCX1i98DSl1jg+mMrnGT7IU
102QPTSFcmF66VBuEjPkcJphF0tXVIXYU5dDScYYxpHKciu1jF0VIk/9dH+nLPo2
CiuVx7xZu8i/g7qiScScFv3b2l0ciNJ7AuVdRbUCoFPpuTT/0L973Ox9Cog03xLP
YCW6L9GAMHBqpej9NsM/05jnXj9V3rt2hz12XDUP9R7b1tXq32et0lgOzOGAYoI0
+1zDC4uxMR3Do4tMOFJ7SgKwjU2rAqko5c2+iDJW+Btd219LdiTZFzG8t5IBAXXK
3NlKJ8IXI/Lqg1Bmzj089m3EB7edxJMGUW4cYk36xFBuADPAEVGTZv0x4i5Y4E1o
wk2Y9XpYELIZHwm5XMusNtV6Bemu5Mw3K2QN7O3gAulG3+rgEoqOqEQYz12Hhxsp
kVbH6ltIyaEh29mLaYjlxCt4OTiQovBDBtelbtfFeRF5bvwFZjswqt+e3duubk8D
pYy2xwh1NOx1zZFMzW6pAhczA+MNy87+dyZzaHwCqfmyVST1XPaEM6K/lOUalGrX
Bque6y9t1WhZ7JY79K8wGLDbNqRBm+tM+HzDm2OvEW6WC9QbaMTLZLTdHbx9y5re
qdur4uZynYNKwKcKf4+zmuDP5gOlKVcZd6a42fLMEZKCVbkk7uGrXFzRPjQV3zb5
JkbE33PBWZPxZvn5BR3JlrIoXfqe5G64hUJSOhRMcIzRHfhIUUd+7Pgz66g4uvjE
SKmDeHARgHGdkDX55JtCp4yxrtD6DMxWFlZq5d4xak6dNlamQLuH0YX2zXb25esh
NPSD0qTrqIWB5mzA4UPw9EeaIqNU2H7CZu40+u9j6Bp9xk79TPCDm7WyB0H+kkZl
PBBYdUZK1RQTAl+DR0AIXGR+HeYzU5RW/qimn5HuFCgSQhddgxCZ407v6/PALDUF
8tcirKhDH7Kf3yOlsuUUaHEE/wl2eSEe2qu4KP2oBx9AsAFBtq4n1cdE/w7CPge9
WSItxI15Lb12pIMRk6MpV+HU5Yp4EXii45hnlycFHxjvoS9XAA6z7FsMOzi+17rU
i+BSTtpaG0LRAEs62hBjU2dhU04ivGax60motY4zu6Jx0Xx/fwN/wiLeyLQMsrSC
tzKxZdUlZnwLcVSrX/MMhVGy8C1Elg+DxWYCnQUQ+S2bPq6Qz25EUVsHLGsvLfqt
SJFp+PFV+My1c8NPxrV+7zp7QF2vEezgFXt+fnomk14YXw0EPhk2YCNqw8FabyLB
PCphO+BlhTgsjXH6Qsk1bOvrCx47k9tJWGS81Ap69x/IjYk2vvIT8O2WR5v8sVlJ
iNZ6Unxc7DtBz/cVamCOfOMQoDGnAghbaN4R3f+IDPdNhJZezCQOMv4m2J5LC1Bs
wRYaM7r3Uc7tRZIKUO42JTGvgPuE2CHwKBXL5tPfqNYDR8mkWKjYNKP4/lx5Jywx
xPFnaEh8e+Djci/bljCbQ9fbm6YJkhdp29x1u/7rIJbFkl0OYQ5PjxfTRLfU/vOf
cmVI9s1Q/b2OiAUYDrDc19OViQM+EP1xD/HVSt1x138dJrb3612+WWc9EBOXN+M5
fgsyxGkT35qrYzGWH5i61tJ5VQbBQu93VFfGdpWHftvCCMFYtlOWncAAoXUfGnGj
jlCcEYOCI+zmPSSQNJ0pK657ugywMGBoZxm7T2VXN6cJTjFDRv2HBhsnxicZFtyU
p4Du+6ibIgWjALdteaUqPMGRhoWG0xz8Ymp3lCXsMUCZfE8RNh2NVAgiibIWTsRO
ZPp5FSJiU9iLGeqlsKXtKNw8olQUzYsccG/L49zgN48PR/qUg1+X7sqiOHDfOr+k
LECCzgGppCZg4FrV3yo9X/SzPowNyajwEo2X+19Sq0XuB8kxlB3qRy/Wlkg1t/LX
r1FsRcSzbDgzXdhEFK+/+aKmecRJoOMj7jNnN9Ee8bz6OolR2x+nXLtLe+CqOQq+
WLGeMlozepLKNPL6olh+R60j/4u20eaSz1ihhpq99thVBWaWNO+mk4KHbbwWYGCy
7xuNrL+cu5IX0nd0wxyrCRM4zH/tulKThg5WkLdWnAEM5jYX7f9B9OmvRvE1fR5k
4F+t1zp/dlaKDwPMCLwQV7q/FzGi1tBdocfqiE531DB2gUpVW1iAmtDWeCWeq8zw
exwrVEkVBguK0b8VSiAzsjepHNQdd7lI4rp8euKv328RPHloRDB62kWUlINdCfVJ
lV86+SC8zN3htXJ8wEy9mPxUexd9OeDJ8eQjL2RHIzdzoolhKLE/loGBjVq1y1DI
4BuikGzMgK5MAMUgXdQLjZu/PR4UfVtk1SCLNhDRsDIEcZMA2Ne95lNkTubNWXhw
xuHkuyvNfS031WZ2acW2RX7+rBnl2KkutChoR9sR0UV8TxkzveMQdyhgG3DcvVNz
HqLCB6ameNMG+nj748KJjGcrkmTgGuaUi7HAbvohxvwbU0lu/z/tDS4kHzl58lJr
Iy72NBXyljPbehrqzPkBznnAJw7ZE9qz0KKPuFzEE3eRIQdjNGvRgDcLePU8ySI9
0WUZJYmAJ4PMAwGvBXcxqKt43MxhO3itYc5rcIJeNxa6s3M6PvMO96VnhyEY7oPN
0akK3VtWVqElUuk91eeA6xGPKgDohVlno7mOYoHmruuw3if4SwTkGxUwBkjRjwAV
H6mbBPPc1D8cqeKpe2OJwpa7E6crL+qscltuv25YDSH68FqOHZCoRGsYa7OGbAUp
kBTKhjrzJOK8nhRVW5fiSJCRD3dKxHe9ApQzUuXLi8RmLBpC4LfRg33CxTWDjju6
pPTEpDNieQJTWhcXvcPqZEWN60O3WrOGqEX4AXwckIkC6hmooeqGvnBvn2zBJ2w1
yZ7Ag2DuD+KEvHfJAfje90lHHW+/Tij3D2ZdO8oC5++cKIDaapcAaQTkoZVg2hz2
CUSfEBNnutXu+LAAL7LZ1wFi+tVVbsJyqv9Aoh2mlD1o3cNuJbCtBg/W4KYXoo/v
XToEFpT03LeBDla9ThDGwQLm9fLW7TgZHkdAdNdax0UdbfxeGmLmA3Ur+Mr711V9
4imwk/mP5KOm42rTeAfL/S7/6FFafioJSecn5TzCD9tEBvqZKCc++3I97+gPtGU0
XkWTTQpWC7r4ssEe84685Z5u0TBj41d8bfh7upCg+eWm5uoNENQKuykKGpNFMJbw
pFNN2BmgoYkmRUwkxFwd0zP5hDXiVdey+Hs1xcxJ7p5Vvy8BrN1RrySSQT31m5tw
pwFQ86u+imSSV0ew94lLT67IZ9u2u+zmWQIfJTfrAUdfdYtch/3LHydGaW5TC4GA
MY6IRRpklcZcR+nJVo7yj3ux5H3HvOmFwjfhTR8N2tqsn1sDbSc/Hc+O2z1JQEmv
TgsN6uIUCG7/17FfOi19rEDoEcUF3X7eOdeR//EbjMxlLLl6CLMyb2qmMV/oLsX5
d8NtlFclBcawSLJHOBNcqqNkLcNucsBkSRmMtkb6zr590SyQ4QQepBPdejE/+lle
UJWARmp0PR9VeObnvWux3sFFuhM5nf2vs84RHZLxGb4oyr1DKNl2YS5/pLLy9FWP
Ja220CwEjK3Rw8mhf6O9KAvy4Y2lvUC/40KqvZE56/oCKqw8P9OdlmWC7fLn329S
nMKrVjaex3Di64dFgnD3t+KWRewCQ1atZdgcOYOKWlJhioY2loPwRQlpwkoDcqsB
bswH9ZdAQlsD2Yh05SjWifRrHEvVzPIcg+cKzOW+LwkRTyhP5R9rFr0qsDlIHazl
MTCFurJepFaeATxIAp5u5OJpPqr6jQ9kecFuhbUTtSl2XTa1d4AIOSGfASjankpa
N5tDEmtpGCIqysblcRdw8SUnbNRkZ42SKivXeh0/bLo+mEDHYy7JTmM8IiQyOoqQ
3naOiL1Ctigijx2XCKcGw5E1RlCMkHGByJ6R2rUrVewPMdFQ4/Lxihlr8olJwfiG
YWt7+fnh35vIqiBFhcGOehZFvmfOVkQLoj/denhA7DjUj6ntKs+x0Jl5qdRibTTl
4Qn65ArJzukTEZwRT8Jj/bheB9rnZds3o81CGz58uFLcuG9wcveTrB3NpehAvjDJ
A+Ym/enrQ8l+/a+aaeW1eBoLd5GJdBSGuA6mRjDyEiYFvW91hC7zFYofxP0s5caY
h33oEeQ9nXOa9PP/bnWArnSTejnNMkloTPiIJXdLt+gW4uJTQtRlrnVu4u5VEOmB
uCf6jYAd4935VL2AyQ8QNev8VBLjfwphxUNCaIaNlwuRd8gn0alMNTGrbybQSN2j
zAFZCorGYV3VvSH9DQz19dSj4p2I9vgDQwm6DHB4JMepgqRR2W3smdRad2SpqRO7
HthCwuWfPcYhbnQ1mByNGf4CYQIrvYaZapVgMbf+u/28CSbO508jEjjnWgg5hNFr
KFvAhi3FoanMBjlePFdu6jIPJ3QoW+x4mtLO5v6fRPEQ5oXZkizjSgVEyQXlJTle
G8K3r38Ej5bF8Q/w9iSHoZKCm1DbcziiR4mkSgZypKLkiyxfZQxqzf5RtL35YgGL
+mXwlGvV9GBmYW+MG0ehJrALQZcblA1DyGTsgskxde9+YI9tTXsQHAXi4Y9DaxJ6
Srri/W1zORPDq16H6OU4XDDPaQIOTgcg0UHGQxbeiI4Cn+7okbcMTU334t50oP/E
PhA8Sv+r5frAwsvinLkyoH9zUXdLbD0iYtbZXR+0FZvvMDD3A1YINN8goIMkm9/h
mgTH/CfiHRiC7+1nr5sWnwwayk5P6QMgy7W/gUA2UML/nXaCC43gMVxzuo6Laujs
frAVbjwtXteWsf5/7LJnqmRi9JCXWJEb0vM7XAYT0zLF/pUZwi2iywWA3lmuC24X
WNlAsbDjbg5k1NP8J41QtZx6OzqHwsWnclzysR12wnm59cyPubn6dHYGpsB5gsqL
IiSfLEhVbgn5XFCrval5TmoB+09pXh107SoSytFPwL/xhslMP70xQmlzi3bPDVps
sfiFs2K5t66ku0Oucj5KbAe7f6XTXi3tyMD5oM6U/XuZlausKHRv1Qmiwnd9fspV
C+Mf0Mvn3NfAgDrlAbsFhqKUsbOWBV+Y6/poNwKBK5GpA0vitnqAIaKnw7/ixB/+
G40TgZJ1Bnl+hIlL/Jo6eDLmagUz8wRYZuvWEHUNM2Xwi5qXnptzVfT83m5Uakjy
j8CtUdCtoeaT4m7d4BO5hHjoQypR7fdsa8DDg/GqtoBKsvsRyUuD2vybvVB0IJ++
GBcs8K4ZxwT40jHkNTXu/okFfKPU5O1zaBHYt5u4roeaODecT2xZKpb5ehxULkm7
t/Ks4/kMyvzkPJ3iwVvRfra9e2XQfyrT6aEI2OMP/TukcozwpDswjA7+g3y5zmrJ
t72nBMieIUyJy6vOTX7RsKTsWucWm5k5zwycKv7lynWvj0ypCHrt/yWuPFvDsDaw
6K8WXzMq6N1qDjJc+VuQhPUb38wJ9CV6nxdSNYj7e9uM+hFmGSjNB0+d421rL26p
xlDKgwn2EGDCs8XT7liuaay5wseVh9nFqvbAhy3oheHYhKeCQKlGD5fIEY1493oP
vjhnC6UoGM/oc5PKrWP6ehIfNWDK2Ko862058bZF+fK/PYnXvf/jQ+JaVOrz2LTz
PwD0cl8BcOCJjjyJwYkWcDOSX0v8Ti+x/Xgg5RGKvvh0PXpNdcN5m32tvsHO4R/U
sgAzxgIwuYC6DAk1NW94rWIKMPenLhMhHWs7no6B8I26yI3eQbeNlmVTXPf8uaPD
Ifb7pErO9XmaSCQymhIxn/c/ZY8niU5zv3d06dt2FdXYFvK4cKFFBdf8wdGQ00xy
tK8PEBc060Bp8nKA9WGAJNwNX5OqzyvtiIeqLiLZYsrGwEm/LU014o9rUHei5ztP
JXG8GuiHRlTrF4u0dVGfhjutAyjKtOLpfUwRObGRjFCMvTtgZ5yxie5+4xVd3oQD
h2I9td9Zei4cC9HOqMleEClUIe/4K+P8vvpmhUw0YsBW7UDwlqcDFUd6xOV8cGvf
7R4zcokwhnK0F94NSmOrjX/srjPovJbLA2Jehi+hcM1ConxXvGdIk98d/LnFcBCZ
4qfM7vsAiOxGR01sisOmObHD9Yd5BEGMF03OOa84tbOidHwbIwIf2bMjU3CKwxlL
STr76gcNaqj+G7NLh22ooWJ5VuJv266u1lKCFjh0nFs/3p4fvVmSRCIuRbxH6Gm6
xHEbq+DxroLV+1ZD1M2kAjVJkkB/f7hxEHyG3JpIkHakslCGLIUIk8dSBtswXxUU
hriXtuRWNQgBC+7tI9KxHVmiJEp16QFbHn66TvnILCTZEVaMIBagLk7O2tCoFiJT
342uxnmn6QpACYATX7H9EoBzNAzpYEc5OkfoyiSUOay0BeAqW+o5bQxFTj4diDRp
tnQWLfvvPYCGnH1jka6iJdkQ0MyM54EX1836r+ai53YG0+1qMfPA3ZLWdpmpvX+n
/uCz/uzUwfDw6M1GWzAKhABlHrMLbuksN489poNShb6C0WKQmIPATlEkfGs0MYfm
fPUxFZ6Xa62lz3mq30EvRWIMnwOwiX9dLOUvsPtu+ZF8Wo3pfLTXeScRuHoQPSsf
0y8ox0rM7hPS72ECJlvniFUT38LoeYaAop31x32G2zETq+Hmp2jXyBxruYV0LsKM
I70RXCxNry4kvwnJFPSWCNtsNC6iBwW0nX6S6XICrLP33x+sWXcr9reoGfyvXqCf
`pragma protect end_protected
