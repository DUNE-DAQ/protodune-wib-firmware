// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AlNWPORFUL65RRR4ExS9A/Lnd75Tx8EcDzMw6Wpi22zJqMW5JyN4Kmzf0kJwmu30
BYHlu8TcqJln/O/21xQB54sTqtK6M4c8IivjBOqEAvaIAEsDlrCYwl0n8iboG/ti
EPI02vVEQLOLgPHFJ5Q37Y2TWDRb9jbCvP0D2KNAVmg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11392)
8uR98D9heuuGY/e8A6WNWHkArKbaXAo98Y+1VwcmMKWslJPF7FoaGqv+ZNZ+d7as
yThYVcUb3kkiYNjCouycijLEPGIh3hTe6FHeZw6vRrcvmvMo15ImmhgKWInynSXe
t/K5piFjNAJ4sTlzI/bCN7g9MAMpB1AbNiqpH+zuKKahLGmyiLI3ilSlhf/zjZoR
WjGGaQN+9jn1LrtUVDBCeZj1xfoVIAbPNg3YdQgJOZzQFQ/6eLsSEGwmgHF4hNkx
9qo4so4xPot2adMpRg5cSoKghKhovCvpS/tMzB0MouTK+niDWEbm8YdpfJ94O1uo
7dRMzYxQI47F/mQe8XlG1T7/WE5ZpAqOagv6AlCYdyPY/6jlQpnz7s3hDjd3usWN
8Wu6pq6cvTWWt5mipD5pxKX0s1NMhpNqvlZdFD8WJ/U0ddOPxsKwzTudLlFagOD8
iQmCOvtSMQ56khHYD4sxLeYCuAd0lmuUoYTSZ655qCud3dZs8FZOT/Bt6Q0MuDvs
ih6AKA153rBRo1Il7O8arnXpE0G03CQndhfrDbHkJb2OfWyh+vOvBo0rYAWOXZL6
lqkgdN5TtV3BcQpIXukU3RFrdB8a1SQykcJJb8OLU9IHzFKWiJoKhkFSL0BJEFhA
OtC9K0qWSXT87VrWwkiLuT6kH0i2qFlHBQgDmYvG9/YYwmHnVp0qMIOdT5etKKR+
dAH0Q8B4CWC+gAhyieUw+x3duAPPfUd3TUorEeSpkWagtUJz3Mjej78OdKHYPfft
+dO3dQ/P8KrCanQ8aJGcUXHmocYLLnSnDNP86H6Os+nTPGSESSVnlTuYdjFciTmV
jMnKO1z7auRgSS6aC36dlF1gzX3GYWAg4V2/b/1ocXqWFUkk7i1mvZZBHWfZyQKb
8Cvf0YNErUJ5m0yxQkNgEQ2y9Ud4Mdy5wV2Kc0m8bFOBaDoamf1QcPYyAcIyUIRc
q/akBA4kubmngqbWg4PEkUuA0Dj8/Ya+FJl2FK64jtg/gq66FsdGL0t6VUyezaBu
rtCqYEE3TzpjLMoMPDcaf+zCjNw5oNs51dHxQpt9D24HIxiq2kUME5Ig1HCkqiV1
VHu7M+E4XaRdwTLdRv/MMzEEdJNbp5kBnwrUuUBCEx7IV4ifutjN1Q/af9MGjfov
eSKHPYTQRCA/9wnvEdYVoP/BdXGOzLvar4qhChWQcpSegFFOnow9xkNil0D4kpVR
xriNZFZ7KVuzEfBg2EUkaCmxHj1SupFLnWaY2xMMIZwLZEYW2Yc+dY09QJ6+DqzK
MThJ6Bq0xforN0clGdD/Y54xDDrN3641wY21hkdpnfGTUpew1TYYHP5bW2v9BIRC
ciHhjgoHmfBbmJ2ZhAZC/R1U5k9ZE761w4240Xa4364GCmhHnDbhNNM0F3cP0D8F
2sZQvz2nC+W/Ns5V7jQ3JeAFP0B1ciDqzHxelOumHLJvUWJV6w56GnnLoDH0iICd
tjgvgmdY+l0GEuq28Gyn0WIa+WZpgjCXXXsFyUJYbkbtDrdJmhbuBQFvjwq+nJP9
tA1esXAKIISL1l3G8Pr8uwb4Bge3G/POSi43VNwTrhOOxvfOWQgp3luzl5dJr5jD
/snc1KpOPJDdfkQMR2o/jeiDG9PkKZGpeGBi2jMGyhcEwC2A7TZprVOQ7pc4CWfP
ZoNLyPYODOWAdan1ttgYDjpVHhyp5s/JY3u+/6D7W0/uwGGl3QhUFvqLEUBrTcsd
qn22PHeBGNuGgQkJVqablEJJyEMyf8owt4YQqp4n410rAK5O8/iUsQaFDZ7nCDC8
rrk3a0SqH1mZZ1o034rIatQIBLP+bYJ6DCP+BSI5WNDYqd1SnlPBmhtVqTUpO+kK
S7ryu5LQAdL8m75d1fobT7mSutTQf/BhW+SBziqYMLJQJ1V6dLZvRDi9W9IHGwH7
HqaVNwjHSmycVZYiFIyvWiH9rUg8b3/gv8bc8QvV50g/Uefux4UUJ0JWhLrLgyCX
UnQxH+UQ868BW8D3cnYasGkViz6/4/ZA/1BYdk4WofpbgZzmd5WyMIgMD5+CgvxZ
kU+f0EYQT7TqJYfnfEpinRA6GaWp1tetFXjh6jTfQ391/KjnL1UoXmSJ1um/MPjE
k9/0EfkvN7oT+BcT9kVi7SysCqia+fBlVjwD+ajgFwM4jBikk1oG2urvhPw9WPC0
CyPaeq59a9X0t0CIz0fRSR6MGfj/1hZ36RBJKtEt5ec2xx4DFaASjE83ar7R/P8i
zwsNgfKQOPvGx63/ksR1vLIaW+wH7i5WnSVu3cCMk+/KoOUpT5K6p0bf6I8GKe5u
jKJsr2GRBFMvtCjtYFsWTcbM9tV9/YhOzTz+2W72EiE+s8s5psOO8PumClbyhc1C
inw7mvdDGRgOyAgZRIVUL5N7tykaS//B7M9lh7QbltfdmbVghj+eVs+8e4wtEhHY
4k7A/tW7GiUOZ3lo59OF6A0TBKDdGFiTdhMZo/FVZcHKNqRTH6aDPDYowKDe+U+U
84Ws5JgMSl5cSS3Mz3NDsEBMCXRBQd2W/f9I8HXvG0NtAlwob8MqAFNYZlg/7Bb5
BHLxVts4vj5GbFyJ7toGTvurUX8J1PnXYi8X3pYKwVK9vyXa0FzHI5ibiEIDkAOR
0OX+cLHzUDMp594Iumg0q44pxZCBTTD5WY/eUjG+z83NNG9a6Osv1AJBzUf1t0HS
+wLNFN1PpvnTiLlKySIjJ+sQyouaQoQN71p891D5yZzQWvJLFKAUroBSW88+Eamd
7veRyQscXzj5CawrCV4IupQ1mtVSURAY+2Z8dqR0q2i7jYVieymBQ35q30bk10zu
YoP1GHjO3onvgmyUQuIEAE3saBhXBgOJH6DAdluGVz7htR1f5Fuw40iTohOKKwW/
SXaEvpLJPQx2paR7uRsMSq+3cMDCZi9CLQP9hf/Xvc+fRgTOGEe0RLrHEbZgnq38
0tyYNXASwu/saf0f6ES0Mx/P0enxiRsSfs6r7Gwsb8EMRdwILADYbFmkLnwbB+Mx
E6U54qCWUgRXgqmkSLMsMm1UYIN/whe083UgKNElxElReYTn/Ztpx6kG2/FFrzn3
BlQxNlh8v5dnWwB1jjpUJHyev18M9S+E1aLTjHzOES5+7Ct+X4Ef8FnJtTGQ7Z/9
y0cLVtTPjua216tCC9Za5RhhLX1itUJKBBMLh5Ij1C6/sN5cCsKxSHIWbBHPGmNo
up/1rne/js/me8YEac+OnYTpOMwSTBcXRo/qUXIFpLIvmqyWeP0P/BFkD5eNwyyx
D7+s25tvAJsAMQb4UFt31UmJCuK+04KnORANg2eBVOg2WmsbqKTOXoxOq+PceSZj
FAPNe+wpcorpnskB30/bZ8sU69fbYjIj5FHxaviLEtyekfim+jGVJdK8oe86im6O
dZJlGro7G6oBxDyjtgd17FXzq4rA1Icw2bx87T7bNeknYln8AnPnRo9krcClddrN
3V3oX5BvFo3svCyxSqgjgXvL6cPhnYfRvngzbZsr3KCDBC+6GqmNH0gL656Tpr/0
QOFhMgfHz0UZcl5Q+IPJfZZFHt/89hI/C+Mf989pmDl+qgMR60H4NmDkPRHgfEiu
4sTOGbZC2XF8tnmkNxW0KEPNl6W0H8Wjeu8sJ1MIqllXM7jDUYk1qhh+tOioiPym
wggBfG3nZPOu5bFEdUiL4iBNeicik043qtOnwCIw9Os7PtcDeXuRB5ZBd8759xUY
X6gcR+VNVrJ0x1s8TYNpwjveGSLppoIn8fmNj6H85xan4w2ufeUfzXyGdf2ZXgDb
VjnBU2P3pQO2GIIJgMMO+/XjmgPeldazrzTQsmZllKWZwnULn+x5uelU4wPhG6HS
c3O1e/wTZwHAWy5OeoES+GapRzijXu8cOE3NFkG6GNfoX7ZgidKSfIH4BHZuIHjQ
bc892OPq5UOT/szPS0VN/kRBBq2vx10Q3cyR6xICDBe1K+QH7YGlMQg5CHFcJiAw
xMcDoRoiwixqs8T9pfxAMcnV9uTEJ+vQOHTAZWQDibOYgjEkCxCdSAnqMGJF1Hjj
pj0aIhFcikNg0IYc7SMWXK4fSCXz0uCVk91MVXoasNsyMqIIEcVQyDWs0sWhyl2G
PJD01bXYbf6DaLFjKO4T1/yApUUhBVQhoJuti226De9Ie1v+NqqgeYkKhdjCujfT
djVbA5NsKQ/mPIPXyeCuZ94+5Rczck5BJptu6ik1tDe8b/xGo/cyE0S/9T2Aw8iC
VI+oC4qs+wJWf/MWFiUEt/De7mdOlxiNA1PKBluo/MZDmmbjLSsAUxXj0J3Zn5fW
cANXdJsVMU6ucbsn3+rste4aZx/JmFW7EduW3dta1lDFEpwjFScSP3f36NHxT2f4
MNqz7CfhY49vWL7QK+ZVdPaRku5MFFeFZkrXqiWALGJw7h2yob33pIe481d/wWLG
bUNqQPPMigSudJgqnlbCq9RY+xhTxMZtTdzdE4T1hePEI3b7MlphgmZibWqEbDZS
i8+Cf1fcAFEuhX57IXRJv4P6HmE3wYWb9pBGUYQbM0IV7K3uOqa1TB4rR9Qj2pSF
2lAtks/63+sgs/oR4gtjfDRQrR800EjuhHvquWUrp9kG8916HTM/EPaY6WgiHQ0O
Pp5OjMnJ/9JuzOot5d+Xw6rCEhuiK32ZxmXDetH0+jmBP7sPTpKpaKhoiukX6fix
w06s7E3sW8vqRAeFWRsgvbSmDvT/vopPME3difMdmsXkB3ZoSnwQyv00nEipfhlF
cdP18Zy0vEzImsdfim4Gm1ntgMiz5HGfdcUE1FRXRh7XoltrJAWfRixC9lb7AqZO
tyJc2MaNPXU/ZFF0HTiFE8cStO/r5Rw9YkTCP5LOCm5enbwkqSsv9IIN6pZe+yyN
o2rVxm4NJWOxm2UmS3K35qtgMQ7zn1cyJepPsleKv40rajV+C2gno3VfvXDBhZY7
DxFlNj91Jy9aX42xOgd7wn6DC50GGI11mghhjsqzrkr+gs4PzA0zzmj1yY+Nfkq2
yQKUp9qGAbMn8MWQADT4uH2ykDZp5440DtqgYzxh+og6Rt2JX/n1o+OodTvNSRyU
ood5jt5ZL84nRneij8Nbpfl9qKPrVhg9HhaNv51z19LCOes+gSkO5Tz9dFyKkzct
JcIhWUVnoWLUnwtkW7/jq50wx1uc9G0oUIc4Pi/4afUdXiGwheLGhPUcpeTKBFXT
Oe0FLjT53Ad1qSbas7g+0VF+e60s7jji7B29nHRTW9bP6bJpLb5hc4aAwpIJFaKk
pSFBkLjYEf85eqORI5eQXySObba72dbY/4tPVOzppksRR12WZP6Q7rAlBIZZ+bHO
OJq14hr6h9OsORT27viM0B912uT2PXuqkiZWVVSfdLrd3PauNwXy9lMAIAUj68q7
zyMf5GWeW8uHwuEd7j+M+CFYkwVcf6HxgUgc73/OZtYw/sq3gdoyITtv2I3M7iiI
byUsdSL/vzikg7XedJzrZWO52H4TgMm/JI29Dxxdu8j5gGcgrDe/Ji1KRVZeA4My
Bi/9w3L9VeR8mEa0/dno28WugnFmDYUohP1gq4l2CNBX0wBUFlI/bfq543c0qTVb
akKh+YsHaqrjpWUMKFupnCxLVa16NNkrSUeEpG5+CqZVas6RPS7EPeAHky+90da3
mIt+FDW8bYEbUCZBtDZwHO+Z4ej/3ARjrNLt4hHX0SaLBl6gEzsEFXzhyN4Frp1j
WGHH3IoSjZBpbquC4roTdEmR9QnljXkIpXcBwI9TdibVKCJhkMHFDq26bZWe/sS6
iQErba5qwiD+MUUH6gDAw4pjvXrvEOzHkVP3ixGjYmbVb4VjkGGr3QPsDSbxsfp+
T1c/43z72xRe7v5y0lA2Xmvjs5xkoP/1IIkMU2kxR+JjKSw+M65EIamnALo3FTEr
QZwmjmdaJ/PzvkHNjl2dMBN4qh0jgGJ/rzDRpSMbBi0l9sIaflrRen7h/wgQb/wo
E6j7M1SzhFIljiVcyNAkMGiWV0pPFtNEV9+2yidR3VeoVz6v/TYudNmMouuiLlcT
Xrch+1LBr/gu4qeI50fBfPG10sKcaMciU01aQw9VuS8LYgQ2HPN8INb76CzJz5/n
38abzPvK7FT7EhhMaLQu4unvypeJ/kPKajpJCEvg9P73dNdKSsBUv3ns14BxOPgF
8myo2/v8u3Tfyy+FRG6+JFrMVlRIBykEfmuNfxO+dnU7mH3uL0YFuslyy6FqZG3g
QebCASjJF2ccxk1rV4aY6196Pt5WC7wZPheOq2x6vEupUjH2T+k/lA9d1P1BIp7J
9xQhSQjg1/QGes4EmWjkt/rh5TMbvIyA/wbJUZDG3o6zPzPkyVydLJpnZ8OKjSRQ
U9fj0X4PJlb4zvs45i2bNOi32EiGxE4ARg+zjJkjof18E+O5ucjD6CmfI49QZsUa
/AtbSBldMqFRF2Hh0big12ZIYMSHKbncsO5wd8PsP7ADrWNUABxsPBc0i2200uju
qkFhnoNJBATXu73Qb6dgl2JSfDeOY3lnRflE59g2QFz5KX3LSO9lSjFlZ8UbshLN
Y4KL8utD1P7QpKOcVclJSUXB3gSLqnY6k0TaQrx2rPUrXc2g0Ao1w5aYzQNlV+IZ
xtZp7Y1xO8RNq0VzyyRuBmhS5U+S6yCF1QC1KB+OXCYkgQks8R0UtUoO42GJhfZt
BpMDG8frTPdo56u24/QsIfOf2u0yXuSVtA9t1x0NQ7VzDxkejevRwwoaAzS9jVR9
h2xSZyZr6S3fbELcLBuXO5fhqiNBANt4IBqzFbl5oMdzncWgB23VrKBRpK2gw13Z
ASvar/QltMdoOUhWLQt7JACBuBuU19frHBFnviDcDp4MtHk4mZTulve4X9i6CZsA
OGXeUElqy2CQb/TNaO9+y/TONFYfdvnd5tmJ0BDAjJAXdWeK/MYtZ+CBcLEHTO5H
jZoMbhaxtxo0jzvcURfZCmfQRZwxJVOH7Y+49hATAs6Zl4rbTYC23lt+TCqKtGGq
tHuj5fpcaqXIAmOqNnfPdAg1FVXrArKe9FJlyorUkRzOHaUM3MnfJO9+mb1haAWp
sloAMBb8iREDKw88uQ913m+dH58CLy2Rj7+8WKgSVKK3+VI/njQ9tkkNsu8uRT5v
g9yOoYQhnaG1AHa0HcpMDpcPBEMs3cfzDZ9eY8396sl2cvkx7ylwVf0YPMnpwjIw
j1QOzas6QXOSQdkEXQRh3XCslUz6RU7Ocm5pL7vtuyzimAoMvIiUffSrtnY8RvBa
rmq0i2txwP8QjaTeQj80zSXI+tE6BUrvPQbN2a+UMV2Wd113zbBhe35jqONh8/8I
tmpZopWJsGKxZbSrFBgAxQp9rbGsxdtK+NuGIYZMEGCdM7pDhIQ1rnCLSZ4amiOF
6Nv1M68NJXlKpjTzFkeUTRT+AuUd2a+YJshILwbnYTXACQtSCC/rf6iIVkks++1C
/Sfu+7lMQi6ZREj4Sy2VH+lDbSDhxEPY+kHsAJVN7hyXOZpPCmXIjqrpRhnU0pY/
KEqnwZL2mtDosRVnovfL14amD1tYZOCtkKHOzup/XV5OtvYa9pmsnJ8/4nGYnZDF
sP7YR1l9Gj2Y+ywlf5g65QXWELW0VM0spWLlf0OQu6mYhI6WqfFGCnScM8K+i4aa
OuDuNwPZlxsu4VHKUTJTOJYwxdoCuCXidP+hsxlLui2H4/z3k8KPjJgAyt/wQdWX
J6gf0gk+yPvEF3tQnGJV969jozqtZVXu10klXUBZXuLtNchw1UEZCosdyhfayFxj
7GqIQHY03DX3/LLv5E+g/l2biXBfhMsEQaU8QD7M08OXoIsT49rrToDqvhDML0z7
hKwnKseb++ZlbKtjqPcaTJ0Qz9dj23NiB2EHzb17KvIn9Ly4Q/iLVxldpwQXSGfs
TeqY3JzOh+lk0/Ky89sTFhVuJxPvzNhb+R0WKBe505B/a/T8bIRUd6C6vLe78nEI
yBJKU1MPZXv/NZiQEBH0GzHDDURSnvUkYUw4AfyiMG6IhtVtBFkkixNckuZr5/zn
RdZs9oZ0bJ5yPr9+FPItgajMe3FhgP/lOFAvUgeI9BIJAZ70/tRev8VoCqKupFJB
OlAPt5Nn5KGXjJAqkiXvsvfNNL7VXO+GzoANSrXHnsSfRsKXP52/1om+xv6MZuHu
Q8t0VCrJS2Q9sbh4aaafl5JwE9AFseXEBNWTyHOe741WBawvj//5UwECno/SsFKs
tG9XEfrHNY+uo9k3XZ6DsBlcUN02TFn+GaRnnR5OtAoN5QZoJkv6vwrETTjLc0ag
dfs1AR0rayZMEtn7FL1DA3TvZHy2ejksEFsc05ZNdAjCx9+wxa0yt8DsfIyypqj2
tV35e1U5HofNPtIXJfGEDk20aWXRRTYfyApAf0O2+f6Xm/+PU7jO3+0k31SyTrsh
tEER2yZlwIao7/dDR4DSszz3JCGck052RA7UGJICe0/VfqTqCMgzKAlO2hQaryOi
OEDaP4eLnVg5bWE/3MHnSMe3RLawpLHh3s8gRXoskaKDGCu75VgBqgcmnroH7knI
26AS3asE87K7Ug6a5RfPxaItLuYxplOL/c61ZgJfBwx1jFG5oHeDsYGb2J8Qm3ge
xeOwKHi4HoDfMp0AhhSxYZahyr1JZBiy2ikJooT5zqdC3zt8VLddy3UWI/FaHLzI
m1uRr4PH9vvRUJ9yaAArHGUB+B1E/KzxElSmcxpqV5WnwpLQp3PyHVj6gvTVG3jy
7dRUVhTUVoTTfYpqAUrHHkdVJi27nIzI19sJOCz4G7IZThNNhUM/PT7u1uV0eO7i
dmKmP59ALoZcPTSlUb5aHj3pYW5G5Rb68fxw/HqeQo/Qpq1VifYHq01TwM5cinKp
tTGb3x47LRqYj64jtlPICYFy58cZsS7DH4G2EOpWs2k4W1hszPl8UViF4/WgJ5To
rot0uVm8U4ugtoN9aGJuO1/vRBl3MFKt/Ta/MhjP0mMXYTd+DlS/4csj1Wufu3xl
CWWttL6MJOInXHQ9O8TebLxCpZ/FjrXYb1VFS7vlTatwdXYDRGnmlf3mGpTAIWS3
iUvpCkMEfFWcRq2E3LkXNpwohR0Oa9KeBtz5ENC67l48dy1oWWuOuU7RTmNGmnUE
CvxU/TpQm5Qi3lLG1XmQekBc/GMMZi7I07cIh309SeAjlOMPqsD8SIIyYHJReLlj
vt+9hloj6/oIeSrrmGV/uwMZvkpXtbzHCoJ3lSVjd0ODZX+3WzFTcbkFPAmjFWeR
CpLDSp8QKFdCk3mclAoU8jisUeYF7YwuE+cRmIwPwCt5XcM1FT/9d2bb9+UcAOO7
wctCM08fYHBCQJzyVEIwV1kGvt4gBQ/VrKk2WjgmZ0HQSkDY3tDPpWKA6IuIr52A
26RIrNG+EkQgRAfeBvqplBofESM8R7orP+HcONTg95wCAHHeonf94S2aQ9QLHy9m
tFfzreutGElyIQj03hP+7aw+dgs+xd2D9JouwlLHA2yqOYy1uHNGLrqW36if7xuR
ZBobZdvHZPVcnQT2XGTqunkYpdWTRZcYupJykiaXAuSm9abptyfwy6Z9L9pSwXOK
IkDagFpw2ASWKGfQduIWcoIvLdCWEhmPhaoKqzugHC+Iv2GOPe+0eO4sL24YPuU6
G2Ly69hCtpXtj7PiJPaZdK5w4LO78WnCste6VWqUWLMIV8cMtWD/QCR553lTc0TA
GKAp3k6aF8+TUH1cxRzzveKG61AxRJG+mimGE2KVQTQN6kyM3eYUhr72hXdrVpGq
7Dm5cNXJWwwj/lGyt3S5BSFvALDXdwVJM8UJo2u9MO53EIfpHzwH8nx6SL28kiMD
G1K0pEKyLb/FITEHR8lOdSEny4A3G/UwXKKfW8YUkbHaxvpqNpSP73TXfJblft8A
f4AR/fzN0+kk0M7ld5sQ4J1QeytQrOo9efiMkKxjP4xaE/gh+VRIR2WZU8ZyUt9c
1djDZXHEXDS6MExJLYeypmW7JYYThHpkWIMKUZkkxlGjuGgxwpilD8xhzMkbAsrW
YWpTU+aZiGZW2RHcuaodOOEq/wf7Cmckwe5LeqULvNzayzBvWwPuu14GtiFui4dG
ucJLePRDBlC5aLPMnidZPmoPNXaxB48Yg7CFJLcUbG4XqgNaUuqXIN+spCDpblnJ
JRxayTA7Aib5tbPF/MhsKnceftwUd+94XuVtino0YBJOE12cJNoILWWSPUxbf1Jl
JzTaPELgQi5Y3i8qXeUehaiB9mRFDGQ+xD/w6HNYjt1HmVyaAQ4ap2SvNuwfTth9
3gMlXO4ElrCg2z0TIEGMzhI+3ZMzoefSCdrIBx83ZDs4V8q+YRWhcp380xSo9Kwz
4Dd5/i6RR+2TAmSpriW3yxE0KJHU8yZbnJhp9w7no5wMuU3a3HLsRsExcSqYj8dS
IHQYGQVK7v1FzaPyxsI4OfM4Jy+16kmk5AsRw0AmMB9tRFrTpVLzDW6BtzvIGUEy
p81IDqlR/H5N48dtpHimYyxbA0xRWSmbqACIGjIwrxP2lhcFYO00vPv1ygHGQt3W
ywVUey9wjLvBimNTgBVEXuvWDU60u8d3wTAziKsa4vcjp4j/Aq111SAVVAJDnn8w
IaaLTI+16SWJIAkHtk3wXGg+I8MbX3MYrlJHZORrcMsjcStrQCb147ElCu2oJBbl
aOifXLmziwgNjGmJ75r+l1qPpTHuCCz/GW6VE6Eb9xe/5j9jCfc9MUisw4F9yZCW
TShOO713tjEyLnEgPMnG3rssftegqsZBFITGX6NSkf1oA8xXuNgYDUjW7iQ8hKCz
zETvDFuiMPmHoDDZ/0GH8nkfyq/3wxjB0q3bhawmHJlzCjlSPPV8mk2G4akzBpCY
cP2GNO8855hSGXo3M2eN2SmXVEVBfp1o9FtX9+N+NKmmcGzkOTs6T80AW/awjcot
k0RRwFyo9jjtkUpKQ9Y7Ehs4awf64swYIaE9063F4tajzdY3qa0STEEzzxO4NDdS
1Y7/EkO3GYjQGg/Osm+F/tx9RSYjjwMUU4TgnZuiW+SYKrirDm2El7PQ1JPsoGzG
KAXrIkrhMJ86eSgqrl7/6LCQIx4Y951rGTaMMY+oGUJSm6DC3aoCBbUlqBuWhZQd
lMw/5zUWRESs75B6fKvi2osNV3ol98Kgtlzj60+G6a0B4OOO++FIgL4L52HJCJ4v
6AEQ3jdcwlxoyhBRAigWQnlYItEc7Yi24OZuFfT1+KPZcrBJwdO4ciJ4D52WX0N/
+msq8mUzhqTB04JjZy+Z6whonTT6t9B2mgLfL+lguOSG+yolCSmMxeonqVpKvNYM
MkJQgnxRTiz41RyvomDfVqIKD2F7mj9bbCMyrD5sJQk8Gud21e/p+E/cYJoQOsYa
fIdTw2GuiRvmXXldeiu1yD6H+Gxh5pnk5u7x5CbCpoAy+Ia0VTJlMobWXFTCE6My
kjbC7DQk63s1yRvMbGqln+A3ikPdo0qwauWWks7XjmxHV1NResvWAk8JWsnty08I
40DJd4Ouk+Qqyev8MFZi1si9vH6seqr+Qf4+GCTLTR+aFdz5xh5GyW+03MQO6HPX
ekph79kBB2vk9s4HZknTrhKzuxIp5thN35nEa/w7tJVcPYcZpdRQ8K9EBHOn42wY
sFR+ZwaRTKEb0ylkwV0DsNlKxt7uH5gra70Zs03jAkrfA/dTxKjcgwP52wIxv4Cv
Dt1nD1jRUIHhARJcgXf3wFQUthgSTqxf1y1LRSL+v7Avi0U6EBCMaRNfunO9K09n
E298hmXlp/qW39ingfJmHaMDCeAMaBYmr0ke5AkA3i+n55xQO0V4KerR9Xkjr0G+
SycIM/Y227h/zl0bOpSPMVNxHZPShxP+7XyB0njHRuoFHgw+Lgm6uEGph0GIgFDd
XoJSwlS85+1YcKqFaPNjj5PKK51JyFCYnftOXXQmN0+AIEHCmjIlilVZAb9sY5+8
MdPh+K27N1BIO6pcHitZVtFdfUWdZtlo94ynHOiDIdXCUvHeNB4GKnFXxewSkYWi
+52bknIc0fKtbTxg9z0IeDt6IMfeD98MCQi05dGzI3NCGkLJR9ZnLMQWfe3OAJs1
EcrV0c9eN9koNy5OWFoAktj/UMCHVAs1XkgQF2uyXAewvDmJ518M6b2DeUFbHovF
04KVoLWFZ0SLQEavDyANPjg7Ru62UQaqjeXTbHbTd3rrhLeeeuFfYPCGQJmqiwo6
iM6iqrI7QarEcxt5nBvGTEyQ4bEORRNFI9vkLyWL0/e/lssSX7717B9BXeHsiYmv
dk5OYvAnNop9o29W4ZLCbtO0TUOmSOoRVPGy297oAe32Cglzr9yHqPBQcaGuRYjf
Xp+2VRulhqRYXn9aWwLBhzE1niJnMbh5qrWR7EUdxwIHgCNsjsFx0kXeFckLIU4Q
D7OtHzbW/wTCwzr7kMX4AMX7pa8G/soi/qWE5xTtYqoJIsMAVXdPUg4ijcsy55QF
usOrlyfwMnZTkHgXcmCtAP+Lfs5GLth291oiRY0t15ExhRA6s9wAV6yqdkRy8jPe
FOnbF+I6QnPhfPVnd+iNOqzl59vnpD9sjQ0oIVTwXnSa5mSlGHqkpslBrslmA50f
DjlJo1N4qVFyNgODBXzgQJCzIuNThBJ1Ffpb9p2H4Zggc4Vjh3ZPLONde0N4lSTH
yyVDPvxLONABFM5+UtaevEkG8ufuGuQsEb8j6YZItC72Dk+B2gaC4ZF52r090zk0
xi37uRnuYYx8Y6Ye5ZrCldvK63pramgHz+1sTMXo5TqJkVvjcqUyhs04hfjXgxFK
4xOYmf87CtK5bvyO8mmx0dAjrGDFEK5+8V31GMdnjNpjibvdIOob4JCDueRC3zVS
ZNOEe80FlZLcl8UNms1o+6VNd94NZW7R7wzfYh8d52Bpjzurfio6OCNeQuVi9o7s
G3WN9KBLfZvYsgwWxVpZcN0orRe3UQt4pNuK3g8knXs6SKWJBBPPzzaXopzdtwZF
ZooDi4Q8MLyb0z9owbIpnI8eE1fV+htnOoX4wlAxJxbmWs9dbLW/fV9jFWu0QHV8
bUDCLvm04XDV0s7w/1Yr0YdxNiB4XXpZlvkPD87Q4zO4SpvWsXkd0Fn4NFZZWy3l
bhfZLsHqGAxAx/xHkVWQYn5e9nHQlJwDYKDm/EuhVhF5554xChjCMJWltwrlRBqw
704MO9S4SHZ/8+RkID6pqhdp4u5L5B2lCJnOYfJ5a5iFh3A4otSH163/REFHz7vR
BP3KurzLzxTddkHJWVT+2N/H9ZjihWangVf/rQVK5la2SL+zPNj8UG6IlVQEFp08
CebZnG09BoARVJckKk+7AbQiV2s7+6keq+VleiZGUy1HZ6bP6WRP52xfAbEcG9i7
HpugKs8y4JQMhqtQup37vYSN/FG4Iv1agOPqbBqfNFFEo8YXDJR0cE9dWFK7O+8J
RA1dHxYNVsIVpJVuLl6Rkpo1/BKKzgNrcnT6bTK/P2fql4l3sNUs2FSmQmGva4Gb
8edufjcBgz/n8Pr7/GUF8J3mk/a20X4GwKKUj6GqxpUgL2IVu+ooY3diyV14t8gw
Bhbp299P6+Duv6w8ZninXWcBDNfT5+4sXnUmERGORAY7D0i/p7c6LaJw5n3uD2Xl
ZgVOQRXLtpv8lmOoV70mdyrqcm+UnjYTASXl0EbkipW1vW+EtM3g96DOi7tAD8UA
ocjuWIYvXUXkWmMa4QuWS5rx1fr1WJbkbzSSe4mvBHxxd1vDX1Aq/Vg+2FIRwrau
7DcfC1VZ8hmMZ7qJCthm/Dj/4dcfJu8vdi1EsE63q8F4n1yspNtxSVIyGEFlcjoP
w3wNpXrhJUZfBRK0t8IhpneI3e3r34fU0Vr6Rzs9OxIOQefWY3OAWNW+2DYC+oJA
0bt/qZDO+K6tiL9a7SUfeysGGYXCH5sojp3EWawGCsH8DBHyxZIRL6GDAclJqWJz
lZj4yB502k1ZGvK70pKELX6nVWkDXyhcCN2JpjO9PLP01COmgh/8Vpey+5gMv91C
zflazmzdzkZQ0gs1/ALxkG2MLC2FZaEOFmFzzdoIKwYxiEislGdxEs8b7XZeqZOe
LTwA/hoPfJH8oNJrEWZ/49VB6VP3PwmpX7dpkExrjeYlVhYTG4RSM0kQMXp24l9M
pKdcPL12PyH9e/vJ15StospJ2T1VAZKkMf2ruZiXXuH5VnU4p8KP3DoxWpuH9084
1D78h+K+/AdqexWQhiMl4HDvYKwAvvbH1wCPKF8lCzkdb4wU27K3J6qnZmkIrmbr
VqFNzbiDv7TmowH1W0uA9mwAdjwiMvXXU3IxFpocid8dGtX1DBro4K5QSXtBa6QZ
VwGNHc/K/TrFG3deeGD2h6WWWSzo+3G25/zBjarcbK1ZvuqiqqL24+9zdBPLgcPK
lK4/ffXm4A3xry+wo/jqiBdG7IlTga8q5ZXpfRF+Fo64Gr5MJazMfIC7v4/oN0Fg
TLdqjGKS+hHCL89baxOL7hQqCq3kM6OvvC/5MU3IpI072M8HPGqrEEsIRILjf8lw
ZDJN6cwz4HoxT9Nktv09ijjPjUkyQn3SUjiot/DEz304dfm59PXzko3Qs5cszNus
Gqc8j+TikpJ12bX7C20fm/OhflfCxQYWzrflI8Ad6S8L8mcTehE0qMsHtr88RIkZ
/3WphidN/rYbWyvvFHCeRljRtW2vCU9NMQsTDIDbMYy5L2WiCyZpx0B6qqMTviXJ
EK21HNwMXHp/cBvT1gwwR23TBLEVBjw+X00PXYoMXeiINs/4+lLyk8BiAYMaPqQ5
0dfz5zF9heoEC3x1KZyf/QIk9u31/VzbrCDqAYlY0RB3H1XXZpjyvlqi0iaRi/WA
OgsbSG/5kVjWycNa4H9rT8qmWoWvIalr8Xbd0kT8ETlk8c3YU5lqxa3owGjBoe+5
X94/ZLQRAApGEAu81/3ZWJJS9epQw9JGl81lRwdc6RL31+IF/G8FIKBe4Iky38Lt
bJ1fQIAoy8lCA/v3hAK5YqwVDUXPyB30rZaWpt4ebNMGomRKbW5e3zVXVo1S/UFX
BcAjFyuVhFplkPvbSs7Qtn2Mk+WC3jLGcIbjsm00rd9mLLgnYaSLeVAO1BzwXHZS
Y/fD+ufk51m10N8DmFgWaRzXB82spTIaEObSZopiP+begk8n+TQyrwvD+BqBTuxW
2cNoSzbrGS4q9zmg0ay6WCfbHll+MxMV9lUAzB8VskVBYhD04AR611jvYbUFRG2U
cKILf6E2jikdqCslHb8oIA==
`pragma protect end_protected
