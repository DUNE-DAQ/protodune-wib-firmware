-- megafunction wizard: %Triple-Speed Ethernet v13.1%
-- GENERATION: XML
-- tse_rgmii.vhd

-- Generated using ACDS version 13.1 182 at 2014.06.26.16:52:06

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tse_rgmii is
	port (
		clk           : in  std_logic                     := '0';             -- control_port_clock_connection.clk
		reset         : in  std_logic                     := '0';             --              reset_connection.reset
		address       : in  std_logic_vector(7 downto 0)  := (others => '0'); --                  control_port.address
		readdata      : out std_logic_vector(31 downto 0);                    --                              .readdata
		read          : in  std_logic                     := '0';             --                              .read
		writedata     : in  std_logic_vector(31 downto 0) := (others => '0'); --                              .writedata
		write         : in  std_logic                     := '0';             --                              .write
		waitrequest   : out std_logic;                                        --                              .waitrequest
		tx_clk        : in  std_logic                     := '0';             --   pcs_mac_tx_clock_connection.clk
		rx_clk        : in  std_logic                     := '0';             --   pcs_mac_rx_clock_connection.clk
		set_10        : in  std_logic                     := '0';             --         mac_status_connection.set_10
		set_1000      : in  std_logic                     := '0';             --                              .set_1000
		eth_mode      : out std_logic;                                        --                              .eth_mode
		ena_10        : out std_logic;                                        --                              .ena_10
		rgmii_in      : in  std_logic_vector(3 downto 0)  := (others => '0'); --          mac_rgmii_connection.rgmii_in
		rgmii_out     : out std_logic_vector(3 downto 0);                     --                              .rgmii_out
		rx_control    : in  std_logic                     := '0';             --                              .rx_control
		tx_control    : out std_logic;                                        --                              .tx_control
		ff_rx_clk     : in  std_logic                     := '0';             --      receive_clock_connection.clk
		ff_tx_clk     : in  std_logic                     := '0';             --     transmit_clock_connection.clk
		ff_rx_data    : out std_logic_vector(7 downto 0);                     --                       receive.data
		ff_rx_eop     : out std_logic;                                        --                              .endofpacket
		rx_err        : out std_logic_vector(5 downto 0);                     --                              .error
		ff_rx_rdy     : in  std_logic                     := '0';             --                              .ready
		ff_rx_sop     : out std_logic;                                        --                              .startofpacket
		ff_rx_dval    : out std_logic;                                        --                              .valid
		ff_tx_data    : in  std_logic_vector(7 downto 0)  := (others => '0'); --                      transmit.data
		ff_tx_eop     : in  std_logic                     := '0';             --                              .endofpacket
		ff_tx_err     : in  std_logic                     := '0';             --                              .error
		ff_tx_rdy     : out std_logic;                                        --                              .ready
		ff_tx_sop     : in  std_logic                     := '0';             --                              .startofpacket
		ff_tx_wren    : in  std_logic                     := '0';             --                              .valid
		ff_tx_crc_fwd : in  std_logic                     := '0';             --           mac_misc_connection.ff_tx_crc_fwd
		ff_tx_septy   : out std_logic;                                        --                              .ff_tx_septy
		tx_ff_uflow   : out std_logic;                                        --                              .tx_ff_uflow
		ff_tx_a_full  : out std_logic;                                        --                              .ff_tx_a_full
		ff_tx_a_empty : out std_logic;                                        --                              .ff_tx_a_empty
		rx_err_stat   : out std_logic_vector(17 downto 0);                    --                              .rx_err_stat
		rx_frm_type   : out std_logic_vector(3 downto 0);                     --                              .rx_frm_type
		ff_rx_dsav    : out std_logic;                                        --                              .ff_rx_dsav
		ff_rx_a_full  : out std_logic;                                        --                              .ff_rx_a_full
		ff_rx_a_empty : out std_logic                                         --                              .ff_rx_a_empty
	);
end entity tse_rgmii;

architecture rtl of tse_rgmii is
	component tse_rgmii_0002 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			address       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			read          : in  std_logic                     := 'X';             -- read
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			write         : in  std_logic                     := 'X';             -- write
			waitrequest   : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			rgmii_in      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rgmii_in
			rgmii_out     : out std_logic_vector(3 downto 0);                     -- rgmii_out
			rx_control    : in  std_logic                     := 'X';             -- rx_control
			tx_control    : out std_logic;                                        -- tx_control
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(7 downto 0);                     -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component tse_rgmii_0002;

begin

	tse_rgmii_inst : component tse_rgmii_0002
		port map (
			clk           => clk,           -- control_port_clock_connection.clk
			reset         => reset,         --              reset_connection.reset
			address       => address,       --                  control_port.address
			readdata      => readdata,      --                              .readdata
			read          => read,          --                              .read
			writedata     => writedata,     --                              .writedata
			write         => write,         --                              .write
			waitrequest   => waitrequest,   --                              .waitrequest
			tx_clk        => tx_clk,        --   pcs_mac_tx_clock_connection.clk
			rx_clk        => rx_clk,        --   pcs_mac_rx_clock_connection.clk
			set_10        => set_10,        --         mac_status_connection.set_10
			set_1000      => set_1000,      --                              .set_1000
			eth_mode      => eth_mode,      --                              .eth_mode
			ena_10        => ena_10,        --                              .ena_10
			rgmii_in      => rgmii_in,      --          mac_rgmii_connection.rgmii_in
			rgmii_out     => rgmii_out,     --                              .rgmii_out
			rx_control    => rx_control,    --                              .rx_control
			tx_control    => tx_control,    --                              .tx_control
			ff_rx_clk     => ff_rx_clk,     --      receive_clock_connection.clk
			ff_tx_clk     => ff_tx_clk,     --     transmit_clock_connection.clk
			ff_rx_data    => ff_rx_data,    --                       receive.data
			ff_rx_eop     => ff_rx_eop,     --                              .endofpacket
			rx_err        => rx_err,        --                              .error
			ff_rx_rdy     => ff_rx_rdy,     --                              .ready
			ff_rx_sop     => ff_rx_sop,     --                              .startofpacket
			ff_rx_dval    => ff_rx_dval,    --                              .valid
			ff_tx_data    => ff_tx_data,    --                      transmit.data
			ff_tx_eop     => ff_tx_eop,     --                              .endofpacket
			ff_tx_err     => ff_tx_err,     --                              .error
			ff_tx_rdy     => ff_tx_rdy,     --                              .ready
			ff_tx_sop     => ff_tx_sop,     --                              .startofpacket
			ff_tx_wren    => ff_tx_wren,    --                              .valid
			ff_tx_crc_fwd => ff_tx_crc_fwd, --           mac_misc_connection.ff_tx_crc_fwd
			ff_tx_septy   => ff_tx_septy,   --                              .ff_tx_septy
			tx_ff_uflow   => tx_ff_uflow,   --                              .tx_ff_uflow
			ff_tx_a_full  => ff_tx_a_full,  --                              .ff_tx_a_full
			ff_tx_a_empty => ff_tx_a_empty, --                              .ff_tx_a_empty
			rx_err_stat   => rx_err_stat,   --                              .rx_err_stat
			rx_frm_type   => rx_frm_type,   --                              .rx_frm_type
			ff_rx_dsav    => ff_rx_dsav,    --                              .ff_rx_dsav
			ff_rx_a_full  => ff_rx_a_full,  --                              .ff_rx_a_full
			ff_rx_a_empty => ff_rx_a_empty  --                              .ff_rx_a_empty
		);

end architecture rtl; -- of tse_rgmii
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2014 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_eth_tse" version="13.1" >
-- Retrieval info: 	<generic name="deviceFamilyName" value="Arria V" />
-- Retrieval info: 	<generic name="core_variation" value="MAC_ONLY" />
-- Retrieval info: 	<generic name="ifGMII" value="RGMII" />
-- Retrieval info: 	<generic name="enable_use_internal_fifo" value="true" />
-- Retrieval info: 	<generic name="max_channels" value="1" />
-- Retrieval info: 	<generic name="use_misc_ports" value="true" />
-- Retrieval info: 	<generic name="transceiver_type" value="NONE" />
-- Retrieval info: 	<generic name="enable_hd_logic" value="false" />
-- Retrieval info: 	<generic name="enable_gmii_loopback" value="false" />
-- Retrieval info: 	<generic name="enable_sup_addr" value="true" />
-- Retrieval info: 	<generic name="stat_cnt_ena" value="true" />
-- Retrieval info: 	<generic name="ext_stat_cnt_ena" value="false" />
-- Retrieval info: 	<generic name="ena_hash" value="false" />
-- Retrieval info: 	<generic name="enable_shift16" value="false" />
-- Retrieval info: 	<generic name="enable_mac_flow_ctrl" value="false" />
-- Retrieval info: 	<generic name="enable_mac_vlan" value="false" />
-- Retrieval info: 	<generic name="enable_magic_detect" value="false" />
-- Retrieval info: 	<generic name="useMDIO" value="false" />
-- Retrieval info: 	<generic name="mdio_clk_div" value="40" />
-- Retrieval info: 	<generic name="enable_ena" value="8" />
-- Retrieval info: 	<generic name="eg_addr" value="12" />
-- Retrieval info: 	<generic name="ing_addr" value="12" />
-- Retrieval info: 	<generic name="phy_identifier" value="0" />
-- Retrieval info: 	<generic name="enable_sgmii" value="false" />
-- Retrieval info: 	<generic name="export_pwrdn" value="false" />
-- Retrieval info: 	<generic name="enable_alt_reconfig" value="false" />
-- Retrieval info: 	<generic name="starting_channel_number" value="0" />
-- Retrieval info: 	<generic name="phyip_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="phyip_en_synce_support" value="false" />
-- Retrieval info: 	<generic name="phyip_pma_bonding_mode" value="x1" />
-- Retrieval info: 	<generic name="nf_phyip_rcfg_enable" value="false" />
-- Retrieval info: 	<generic name="enable_timestamping" value="false" />
-- Retrieval info: 	<generic name="enable_ptp_1step" value="false" />
-- Retrieval info: 	<generic name="tstamp_fp_width" value="4" />
-- Retrieval info: 	<generic name="AUTO_DEVICE" value="Unknown" />
-- Retrieval info: </instance>
-- IPFS_FILES : tse_rgmii.vho
-- RELATED_FILES: tse_rgmii.vhd, tse_rgmii_0002.v, altera_eth_tse_mac.v, altera_tse_clk_cntl.v, altera_tse_crc328checker.v, altera_tse_crc328generator.v, altera_tse_crc32ctl8.v, altera_tse_crc32galois8.v, altera_tse_gmii_io.v, altera_tse_lb_read_cntl.v, altera_tse_lb_wrt_cntl.v, altera_tse_hashing.v, altera_tse_host_control.v, altera_tse_host_control_small.v, altera_tse_mac_control.v, altera_tse_register_map.v, altera_tse_register_map_small.v, altera_tse_rx_counter_cntl.v, altera_tse_shared_mac_control.v, altera_tse_shared_register_map.v, altera_tse_tx_counter_cntl.v, altera_tse_lfsr_10.v, altera_tse_loopback_ff.v, altera_tse_altshifttaps.v, altera_tse_fifoless_mac_rx.v, altera_tse_mac_rx.v, altera_tse_fifoless_mac_tx.v, altera_tse_mac_tx.v, altera_tse_magic_detection.v, altera_tse_mdio.v, altera_tse_mdio_clk_gen.v, altera_tse_mdio_cntl.v, altera_tse_top_mdio.v, altera_tse_mii_rx_if.v, altera_tse_mii_tx_if.v, altera_tse_pipeline_base.v, altera_tse_pipeline_stage.sv, altera_tse_dpram_16x32.v, altera_tse_dpram_8x32.v, altera_tse_quad_16x32.v, altera_tse_quad_8x32.v, altera_tse_fifoless_retransmit_cntl.v, altera_tse_retransmit_cntl.v, altera_tse_rgmii_in1.v, altera_tse_rgmii_in4.v, altera_tse_nf_rgmii_module.v, altera_tse_rgmii_module.v, altera_tse_rgmii_out1.v, altera_tse_rgmii_out4.v, altera_tse_rx_ff.v, altera_tse_rx_min_ff.v, altera_tse_rx_ff_cntrl.v, altera_tse_rx_ff_cntrl_32.v, altera_tse_rx_ff_cntrl_32_shift16.v, altera_tse_rx_ff_length.v, altera_tse_rx_stat_extract.v, altera_tse_timing_adapter32.v, altera_tse_timing_adapter8.v, altera_tse_timing_adapter_fifo32.v, altera_tse_timing_adapter_fifo8.v, altera_tse_top_1geth.v, altera_tse_top_fifoless_1geth.v, altera_tse_top_w_fifo.v, altera_tse_top_w_fifo_10_100_1000.v, altera_tse_top_wo_fifo.v, altera_tse_top_wo_fifo_10_100_1000.v, altera_tse_top_gen_host.v, altera_tse_tx_ff.v, altera_tse_tx_min_ff.v, altera_tse_tx_ff_cntrl.v, altera_tse_tx_ff_cntrl_32.v, altera_tse_tx_ff_cntrl_32_shift16.v, altera_tse_tx_ff_length.v, altera_tse_tx_ff_read_cntl.v, altera_tse_tx_stat_extract.v, altera_tse_false_path_marker.v, altera_tse_reset_synchronizer.v, altera_tse_clock_crosser.v, altera_tse_a_fifo_13.v, altera_tse_a_fifo_24.v, altera_tse_a_fifo_34.v, altera_tse_a_fifo_opt_1246.v, altera_tse_a_fifo_opt_14_44.v, altera_tse_a_fifo_opt_36_10.v, altera_tse_gray_cnt.v, altera_tse_sdpm_altsyncram.v, altera_tse_altsyncram_dpm_fifo.v, altera_tse_bin_cnt.v, altera_tse_ph_calculator.sv, altera_tse_sdpm_gen.v, altera_tse_dc_fifo.v
