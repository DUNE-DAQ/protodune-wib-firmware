// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
enLxGUhFk5YaZFdL+QkqBo4XePscOVJxmYVkPG2/CMAtjQ3do9O/lbdbeEkz27sS
UodrcwN9tJK5qtrFm3mUWl3HMp6S/t5Ut5aoBQmVzxqVKvoo6bOuhu+hRNT+cMn1
1sWclQroPfLT/XV7qfYMnv8igMOskYvoVwd0pInTRAs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34480)
/ekCmqyu7QM/FgkhBi/3D8xB0KNCrv2gBkVT1b/h84MsQfF56sYVD/XL1eHOw0KG
yRgeAo7XVLUzC+qQDZZqxqAnhOgXObn2k9SIpDtddUb0eWn8/kn8EjSv2Gq6yXVm
UY73ar6dLvlDH6jM636lu7jzBKS13TIPe822W/zFbu1Q/AbL1pOtv9AmsL/E3rw8
rKl4ur+GCJcf7h4midyfEaxoogWdWSAdFcZtQw6935FILzdnegHfCtjiMBH8sYV+
t3XTYO/sYFvIA4mRf6Qkh+iMd9Me3bqwGodITheCd9VpPcC+VUzT+Xk+f8X7Js+H
dZ6XwQOPu8aUiuOwiup/pFHPDaJYFyZbIg3JW9FFZUeyOvLMHQR8qIbj7n9rdV9A
SlQ1hasvMz7iTXCuPFvABoZMoQ6LxHS3/n5/5zZO+zcSZwtfkJK+OHKsscZlSmIf
KTez+vmT5Tt/QRv8xNbECO+fLTIr27wMqL6TvRjrZCSedjcqWzf8frksBhjzIln4
zt6R0TFY0w8ShX+g5bhqbzj9DfmLkcJhwawq77z3aFt8YP2YrZx8mrlRP1Qx+rwn
Sl5IMaGYOJHcRILcpkCtiz278p9UdOt92sN8hDp6dlPu3FYzJsPdiieSNLPA/sfT
GFR/IKCIFbBUu5WWqvzKNX97D3MoBbRqyFD349h8+aZ3lYBxOyiYIcwwutJFXeIC
K0o2rsJjZwwvsWMydczKhMbyocYQRUC6aEljf3u4n1aT8t4FithQU5jUVJVQPXPZ
93BC9L53wG/acc6oDYAaOrYNVvCFo2j7rTI8ukI2hdzKZsuzGUtugFXnydsvNyU7
mzdahxnjSSVDmGd0wbDABrR5F3VuV/Vm2ARXxb2CQ0HVoCI8wEXqzcA9oPHXuBd5
4wOGCD/M5Nqxp2oUHOi5q5kXsqeSRE2a8HN7RjzK8pdUYB2UL1K+hp9RZAgjHYW5
u8w6pQgOm8PnD1xeq+2cX97WpI1WmSlf3jAy1omslGNpJV8nINAsiiap/eO9VBz7
OrHsDzo27vBc59mDcvE+SLrYvfPPco55Ic8hJ1FhvOVO+l5lhWuqHo2eeHD4diIJ
6kWFlbRfHjaqMlFWwR5gjqTui1TFI4CyrS1zuecwBorwMi3b62mzMS2Smmpju+V0
tO1NJu1RcBmAZ9H9RpUXK5CJi40DCsTjF0sPALOAOcyovwYcsT264HGZOwFKmgB0
R4FeFskfN6FBBqvXt24iATS6ocr5ReKPT+OMmapBLRh9gBP96RE8/TRfS1s4fVBX
x0trQKWpU0RNk6PlfhFhySGR7FfJPcOzcT+llb9odzRjuDsTzINMrEs8eM91Bu2V
beLZTMFXuGmQmRvei4kWM5G50v3ObVRSmqixWnX/HcTwYHRwQjYMJXTjh92nnmdV
xuc7/vS3//Jg/pUbg5Vtf1iPMmQdjuVOQsFMIZ3BfqxPE3QtrkSgQ5F7+1KviYtu
7Dk+MmDXH+nBkAtWIZoHO8uU78AeuL1iPGB+Nnx/GIEm/Zq01l+ekRp7uRPKU0YB
y055yPUsvxOidtgTUNRF45g0q7UyOuYvzr8JHUTEr7H4GHlDq6R6NCLfjuwF3HgP
tJLA2z4b2S6hgLvqOaPGCpYjhBsl6oyYba7CP1o1fjDBunK9g8dzLt9dAw3DFHyY
QeyY6IzP+WOjuqa++GK/CxomejEMcFF+ynaLzP7EjgIW/rfUTrasrmPh8TzYdpLP
bmWaywnUQTm5YYK9nQrDpgqL8TEx0dRwBbZIuba3X0ZtxzacpH+smVScIdP7cg3i
7robuqCMtEuW2ApBGaVFY2dBPDvDimKBs+7VIAiEhM11cknIMS1GJ3A9KEupI8vt
Xp4IqUz22MPJ2uOz1XVeoWtY7HGZy0vvzjFmrvylPzViHoLaKI7V/FBy6OVz0W4C
caYV01uw0b0AEFZrqjG1ItpSV4HEVBJS8ZtWrsrhMG2e6tzkRDHLRf7yLotMEdEz
APjKZqlBAN97iNWAfYEjo8pt+VgOCDzKMySAs6CcO6Zg7yLVFFiu4MbyhoeOaZYa
JOeorn8TIqwS8WS8vMpLJXRhu6+knTnGDv3jNNq84hVPuVxGLzMcd12AiTwzuJ4y
G2unnwx/pXEdYoxHAA7jq8IEQ+yYvOL9HCvJsjAGYW0VlzfhKUNslU4uNYNZG2r2
bc3o6t7jDNBUqNAFrReHVnoCt0pfjMZ+n6z7YE0eYA6bOh5EfqHqCAKqfeiZia7g
coQ3Sub8e8Armn5j7meqVp6oi2FgrD5CZTQib+bXf1Y1k7MfJcQnB1ch7/zlvdeo
Uue+aDKBuU6sQ29QhD8pzJIzKvCrxIriUb5aZzN6Pf4hdjTD+L4pZX6emXHU5bSw
1/BKzvQ7Ud6PnaBzQaxr+IzjP/PJW/rk17VcV57IIBPL/by3fInnmXolM+8pb0U1
EFOcOcMzuJYF/jypltDYio9XXsECpB9N99NfzXCYAaJY5d2P4jpg0NTiBahRyyS2
ylbV309IPqAFrGs1s/mydYvYU0z85Nv48jgy0L3+ewhpIY1n9fSL57lqknX44Vgv
A7YSfwu1Rhq7YjcCRFpWOwENim7b8HT60z8UGIFcUArPqBohbjT0W7f26EGyjTly
OOT/WUKHN/yal8rmFkMEDMwsOTKmcPT/nx1Xb8H6sE3q9dFQozqyQNhXD5iVPMQQ
fAXBWPKuugBNpDBXiZGhu0AyKgUrWZ4ftlS6jWjWq9B69Q40N8Ce3tjDD/fvufxt
DSqKzW9GG00X+SkhzJaKqOw7IrShmlVOwvZKjGT7ZMSGPmh7oUs0Jyr/TCzPPEP1
79r3tQE3+Q77TJe8zPsm3VHMcMoTWi8+P+Ogk7c7Q2BbIsFMQhT6WRPG/xp7jtDu
gpSTZwN8wKx8PxLhYfDgKfuQ8QVgMtO/78rspERcbW+3KXUqBYLztbXVeOyGCmxr
WoDuJDWVnrafhgaBTxeYQwk23P3Dqpq750ZUdPc3Ew7mdwGQDkBAdDU/QLY+2dcQ
6UAEXgVC7iiPR3mMJbiD7pW0YJnI4Pz7felgGXUkfuhUYfIHNevqJqyMrROK9uE5
7Wed8FE7YqmUKEmINHjDDouniyzaIWffUWxPaG6M+qFVEntNa98/oJUfiZTJrTlo
qdON34MfHDv0zzIFXgI5yK0W23C/QLnqE65PgDREuPjmWo+MFn9ydg/60b7ECjrS
PRk8NIpJ7nwhSZuwGR+HoHLH9uZXUT2V5xLT26zLOv8I2AxgJ7SZk9CXE6myc05h
A3VViULoSFTM20gtz9Sezn8ECmmrtfFoxDJwE5BmdjcI165KKiO8aKjmsc89AFVi
F9d7mmqY968zW2ALS53TiuAOgdI6dZg5pmfwLQvc6jzG2peEbkc2ODIDNnHr0lSQ
wGyDqKiN9ge1oYdFzgbsNHGe+vdH8UUmA0qT2vX+w842MHz+BUN2NVskZ7RdfAu8
656nyq1ynquu6klQluqKdXTirKmnZgzpsGpR+g2knnuDScU2P44GEwJlM2xun3gu
wV+kDZauYq2SauROxDopCI6ZVBonM1eWESmStucJtFy+ssotqFA1iKn08BECTe1z
waPlh0UD1xQG2rHDE5aO64+sPfls/Pbtu33RLYnkuPHKHta5l8SEclqcuHMrqst0
d0SI/v1CGWjwbi06YUhoTBQloUVpDUQUTrQuPVmuJevpGD4b6Rs5g6/7gZl15z3g
G4P/FIIK2V0kg9KihpZO1sLlA/DqlTuCScSyyNkklwNE/XsWI7WN2hBJZELYykJU
yuPcnblpsGtPtmnprMmqiMONK3khmJA7+ExllgAcb9VNhgaA/0rTaM6nxcgWpg6T
P9HdHYIY+cWO+5QzUP78ydD39dPGULWYwpV1leF6UelBRYqQtPtI/ONgXt56dgRi
x9U457t36R/9Of68fBK/FYQJd/fzI3NI/p3+f10Js5t65jW05y+785nbpb7Ad2rA
Gjtun/6hiAC01VIIYJtY0AtAUNpG1rlzvhA8pQcVVyhcIp5lY/Wbs8sSUY7KMSqx
n+nAmBxDGD4WY1qJOQZrbYNFD+jiv04HSkDaYqScUlqPV3PQDgVvdBWzB4LtTr4i
9048mkJ5AFUTBvWaskkkdIST2IgQXdgzyQ2/KeiWVEWh7QEJ7uOgcenyOFfLuvtm
iSTdayJXIIcBlWqm/6wFcTHSXqSkeZ1su1lCBD4Um7kG9HJ57hNJmfDdU5m3Sdb2
U8r7fQo2V4dqocbnTktib+RJlf8NFpNR5Vtrvgsek313QAfmr7ecmchx+x5K+7om
bUes+cOU8LqZjMhhqt0pnIb4HkzbP3u/Y97P63nSA9Mkxsdx86kzJacFen612C69
DGdcTZSiLYVu4ItdtGx0Bi3BNX9sO4qJnZzpW0RS+nwVK988BdWXcE4KH9Q9M2Ai
Rv7HWhQWVklD4jmKpW1j6Vhca7V3VFh3IesqeRzFSLFC5in9ah8qlChekTG0Vvmb
wau2nl6hufgW9mcRYh9XxZrvhfTZP6xiS2d/7w9chBM2LYPn7x6x6ogruh7G1bSz
hmdzBz2UO3iZJpInQyoYhFUx0ri7HYpBBOW4jOCRF2dz1KQe0/Oq6gY22C2bKBdq
KjVeAMg+U8yBqK5aVsXtpOwtuQ11U7VtPS+G6W2WTXkAoNp4D5iOnBGohMD/XKLF
yDJPSJC8/KALvf1nytfZXI4Q0EmDjZqeJoNuzoEclKN8OmqYjAHg63400dbgCW6Y
CEUnAuRs6gmT82LdcEZEdWH6bZdIkhBwht38EP/uPb76Owuy6zJjUrak9D9wfCOl
l/uNuLeIuLPobn2coRe++tFupjfWe0o1qJFQTYn8rMriUmysQo/09fyDk2NhrLtL
b3pWXjBUNyarf0QeLEQeXK8CwP4Je5q1WBq5xUDrn8EK29lzORyctYp8xYuECPgu
iy9pMjix+mtrSPRo+X9REEoVLWjLtezB8+0eH8Q3vW3gs+43ELBJnfFNybDJay/1
HtxenZGlQbn3Lv68hQdaZu3PwPdN5DaP1yYJm0sdNA8mpHNWzaZfPlafaIudR1Su
8lxHyVG1RWGm6QRyqqW70uHamxyUMI8gM3r5aBr3Y3gGh3pjXuA7De6WQAhqs0uC
LSRcHTije79/G31u2MfZtXIGDW1ZIDbTg40pguTDuliLcX+fX86JLmVkxwO6PxVa
rE/RMHMj14jWS+WKQQBeY4Wu2EpjujSQoJvBQeX6dofWzA/xP7ZNrgr7whCD/Sf0
DDmldjwqFWG9+CqBomB5Rotqreao1PjVDm1qOpYsJGvO7xnBpHIeb6x/7Wmxyc4O
/+VKxQirBTTzRwr0QN1Cj12bOMxOobPvHlXRSHlan9ysv6LKrcBWKZEjqQx0l2Dp
tE+F2t5Ad8USZcJNx+dlPqIh4dmStPVM5c2hm5JtKnIhmVucEVPd8VMkCyl+29hF
IX90NHG5vL0tPb6DLqoEazhnVV1Jtl9MUd5Dr3tX9RdkJy+bzg4mG30Cxn7XIkhZ
ep1S1zW4/VeMAk3fxhz5h4Tx8rZkkTP7HSK2XneLoagmuZOVea5xw9ot0kxXuGcV
BK8xK/B2w4EddeyODMnq30zvyvZDQLaeLU3TNGykagk7hC/Da3EnP4k+3KaMTyct
gxreA58hPKXDAAayHgaUrcshWYUcwnxlWYB2uaN7iudYGNSkoysmaJCB6E7SwhJj
oP2sHvq17KNvuNnJgS7aaU4HF8PZq1VsH2aAaLfgpQd3FBJMxWoQdWWaN5CV7g5g
aFIZgmowoZ9QyQdSZIg02Zqvn6jWxzH251UNZOzddJcjc0FXdLRNon5mpgFeBRJ+
u3NClo/kE1b1NZ62xeVkh/vP+2Kx69louP5v06t85Ale/HRJkfpgX3NlFuqb2d37
68qAmeNL18N38AxgPHSr/IyON4AIpb6IaNElRxk6zGEdy2R87Tl95ctZuVhZPQmG
J9JYqkrHQhT9+aGcoGpEVxEOVdJR2Hve7Vqq7p+udtTul4fNCQtg1wCUnei8rs2A
Dk88J1c+K8nqXlmoeXkxLOHBEhL6Wj6NvhbD04vf6aeaiRmz5JtNwcPLJf+qPJTA
CRElyaWjqLozRP0xpsD5AnttFoIP71v1TnbivCL+oiOyjJE8eGBzI43V12QD2n/t
BgMWMkCVsLVpZNogbxqM7ovozK+MG7qVw8csbQGzP/oPGvx6fkkjIF8wK9tdKaJW
EGuRvmVPUmTVTznJU54yTWsJsf4y9qkVkAvfPo+l9rtvJtxqNk3V3pCd7LNjWelg
ZbdtsytnEZB6XRqdpMvLX8XNPfVLClD6DxL7hd89u/2d9OsQxvVMC0nOLtguPK+C
8Wdo1mgOn9pAiygWqT82ip4CrEcQcu5afbT+Tt4II1VaDL1ER2oQ/F4/kfWibtu/
7dVlhQ1/apV/uZAJ8OQoNHCgNMU8Rm5hYdDX34j7ml7h5khb8f/lo8Q3L9MgK564
S2jvv26bP3XQLcSHiIcuj7jKC12va4ZgaYpB5DvWKlE5ovmwju+hdOoUP0fM+Q66
IytnKvgiMZu6dw6e8NOGJfXV7ie3yhbMmR15lSk+hwlKDz00WOGaQxWB7wgoQBgE
7+OJh2mIVefzwtxgeXiXBqpdhuvcr7fC1IQmOdp0GWxfJAR2XFfOUqJufrvn/3X4
7MOpBg9eTDTspznQdxNBHIx7xIA6SUBC7rS5AIooXmWjaJ4E1B0kWq32SbSOHZeu
sX8znqBIbWnzbo+z/CGU4sguXHSnjDM1dcpMsGPSTo4zI6GBtR3hETTLwk3Iq65D
jNH/iwPA327L0xQFflAuvArvqI6kp0hS2m6SQDrijYi+RQKSOfA7z0ujV+SCMK/o
7EKghCucnBp4FgtglipEZ2rdkKUuwHRFRi9/LcOMbDHyjtzo9jWTTkYPqA9sqpzy
WHww+Qo1RXDdIs8M+IfSAwBO5jK4uvv5rBH2bDy2TGua4ptdykL1fVMibCH+ie9F
azkj80eRyWB2niYUdYmUHNOwaQMlfpJs//L7yAWDrO6ra7GhETlpBpZmPT5HNyon
3tsfOv1pWR6G95wH9Lf5duhAwHqQCnlw554+/SQEVOOJoXOhwb150QEMNCj7GGYF
8PX/3STVHkdxXAh74Y+DbOmtKSmeQpq3CxVQ08F8WZsDucOijieoy7B9SgaZfRZd
L2GQf3NIOZknJGlnFGvf3MsnMl+NLImN9F61wC4ig88t9nhHwtHj/aowBcq4acDD
OHqBW4fA9tzLhG9ZaoNFzJH+CZ1xyE+3TNdBXb6XqaIqOmEMzLPP292cB0hv9MIA
/+NQ3ldydP6zWTDes/nTr9a1VNWHPmLujVlnKvT939b4q4AcbEszS7nUmZ9zRt+0
Ml/jU5otJnFLzlb63xP7rupnI2eEK/Ky757TDvZ7280+ZpKi5EoTlPKu8mr8t8T6
9LAo/IMiZsyMtxYyOJ/Y74to7GFVGBRy9+GNS0M3DR/vvnxD5vClLZqj/tKfb305
E65FruF+rNPKHeVcUiZkbnC6uwVCKAlxkSHghwjvUvyy0A2OI6bPW2GsBDdNP0kq
6nJ+ZGBNyO6+m0SPvtaaId3Isw4GyeVQcGFNLega+IqlkmB+GNuzE1DJ8gZe8Ml5
1PaHPwfObA8MWqHG5Dd0smPJh7RXDiyPZPkOMjT3S22qEcaSUzkkpM/ykvmnqwud
JMKHi8X8PtOaj+toVkDKv+dwergiPPHGweg8hUnfmPJCinqotxqehH7sGVNafeza
7roWq2boYrzBq+HAtapGW1npilKulGgLwKzPq3LMWiLh3ChaIqNWZeXDjGbSqCP+
h05EJNLaX8jCyQtvM1QaZYuLu+EdzYQk1qUoLgmI06YwBNi37/nM7zYZg+rcG2XJ
2Ev7vthGhlEtFTfcsdWkb8kfvNiljo4YtsbZTLcG83L0Ka97GnugsV66CkmAcX3K
2LSVzNnKuN6+rZC5jmwbb5BQ6y1oMpRgMAPCAQyoxewIBrC87Ky4g0dHh2OxzujR
f1vJu24BpbgRO1X0iPapIhNCs7QGwu1lper5ncBqZyI78Qr8vcfOC0himlXKboJ7
m833LEtPX6q87eaAlCrZJ4t/gx6uqdFdISCMTyEFaof95JEPvEKk4V5x2indShID
cKDMxhoo8l2QG5dOhgRFCOweO1Oy8XpNI2vis4hUdZ+TcVPGcTykNO///4jC2lqA
VIlYO09k0g0wsGs1yZoWbqkLD+xAx/WF+v15OO+PZa3xPwr0/jVPqiB6RJgr3RZ2
QMbdM/2bLwYXa7ksEgYjyltiwERohT2vLvzBpqtEltMLjlp4H/uLJtHN0DLS9+rf
PF974H2x6zEc2e0qpwjWZBx05SHAxmw9/tDQAAJ+DApfZQ4v4+RTwM7KbBweKpHA
vNhHZhmnp5iEvhOfxGPl1v1o/NVtkcsHh9DpyWcq0QKT9nu8lQw8BjYRDBxxNJ4D
71Gd2/qJNKlONb5biDZCmlk2CED8+rn4Adjg98Ad3QeapNVE+HALTGKY7Mc6VKPT
H2VH0CYwJ2+vGza2HItciIHPMzgyXt0yOAQkiDQv6kgdvCEDmyC9LYwmoBFiF2AM
4qjt5YtO9hALUSgWFAmZd+8jqBs91MDRem7+pqElIN23TCg+1ZHpLLaLr3yUWUNG
ZsaI13VndjQW9/CHC9p4U/v3lwEvm+TjmMH4vP4nAABhTGqSDXyV2BNNCagB3E1G
WIbfcMV5l1zg0vfK/xLrLRfnO/rjy0hTLbDpGbcjSguTudbzO6CXZkruMzfPWQ9f
IK45kdYUMCD3prP+SPpI58fb0PBPftWGqq6rPRJSppqzGxyO2ZH1wKMPSovU4NfI
swQvQzRzlatp6gDyugvqWqY4rWm7OcsSyHjrHyaaNz4CZXY5AuEf5AScyAqkbX2d
WkyXAizycjZXSFCGiP5xivnc+tOKpsz+UzccKgcfBXHJc6RZaRZH4sKnDf2Ok4ld
G/wbCfBY3fcaqV38MKk3axVFHBzvuvQLtfLnfQbKIfCcjWeTj6os29PyZWKaZFqQ
ET+MHtdaLj2KZr5ap8+HjTCoVoEoE0Gd+xA3BZlVpHx8EOgU6jxEEnHn/dRASsc1
6rtByUljPe+egprYz4KwrbxxeiSH1MT7npCCVPKCw6IYhSqH7UCLCXS0Y7rFVxtZ
t0YNFlFoiA/O+3Ni3tWn3fVvAQL+VdfZK1TbysbU3VzR0dp/A26VmlYOfLQ1A5N8
SR54kKTytNDsqbNaoOh2ql/PnPvCpEOK0P+mOpwARbhBwQIZB8X+KLZOZA8YV9wH
78L+9f8BxABllpXZX7N0Wgdw+YqUWNFvt9CQVr0Qv3gmfNYKLr0cHxhzkz0+tlvx
dbfE1HbNqLUamkiEHyTtQLzPbaCWctdVWi/n7m54NXKaD8NvEBQ7sdxJa4uidEOw
g0TN/Yky4eAALRYhiJxOGd15/5DyyBkOGzKOLCtZkWdzKvFhW20G5SJEpW89ROcY
BzBNch+6KxSj643l1FBJkhzj9sDRCCu/scI6uOCVcVue/Ziag120+4PUYFLWoCg6
VKCVjj0ApeT+X3MFIUrU5ky4XMbg0rl9Aw2lQOKqMCr7smN/f8xDt4czqU7ASaAY
95SYk2Xmt8dXBrGuuKChnsdOAkn0sG/XvW6R1ewSDemqsCdEF/eEBA5VSmoHrLQK
002l+MerJBGVMr9gEZIVKBu7DikdXqdCBdPCGyBtqOt/PD23ulu/evsXYxj/WmyH
iXTptPVNCTGnfOw9vL19Djqm9FrI47hOYYILXeQpLtKKU5B25p33TRXKKscsPVzu
bDX0zCCjyvhqfKql6dstKtn2xYgxtv0BvIQi6rG9xlM4IS8OaIwCZgrx8X01jd/m
tvYcVoubsDi1yE/hyVNA63PkZU8ENQcFbYWtHlBeu/61XmqHFgTi8rUd/AwI7ooT
FylFQMl3bVl/lB2DDiHhRGOGCGZZCftKHlPLAAEmgWa4MJ56Mf7GwmU5Fb9yr+bF
nGrvQ/ausAriJdrQZtxDtDDrAhm0LUPPuujdvDMKfUnyk2tyhLhoD64cWAfp4c6u
GKw11s4lANPEVyIeOxgb87upVeq/q60zTqaDceb9A0H/O3ScJyqbs9HPHvNGs7D8
dk819mBPUy5JWFHiz096RRRHLKpyij+d2yaArlHtrAe0ma4BshjGxRxkn2Vs0ZkC
6R0p4QnqhNenJW3CMB7Acwm+VY25lqlDW2KGTwwwPpEA+u/CKPCANbJ3OjCnj1DS
0VDGTrGQkzb2aGvqxCKphoPrH/iNGm/Ys6MeLPo5In2+5/fDveSAIU9z4+KrnXd9
E6BhPR9PzExp1SN6u0s+OVsx2XETjwSmXTC3Y9I6Fe5gm4z9Z1xkxjILQVemfqHR
ScjnAACUgWvwlMju/vy1wj+eBwMNNDB2Hw0RxFv1kSyjhytdioiDSDqUoOcrNmmV
O79z86So4KljFygX2neSt0MwzHNZSRXn+qqgW2kEwRnAK67aGsWdIO69k0xVpqNg
OURHBjh6xihE3Lw87Wp03oVtrBJiJzhvo6KjNnl6FU7uPHrJebjgNGnTipke8Cpb
3d43KXLraDutI0J4dgz1vf1C1Uout3w8TgZ0MgIhB46LflGy2RZTT691Ne/Xy986
3WFcPFmdsRPqiwJmo8XamfEn/2AHAZCd6PJReveDw3rXh33MjEGHJb74nt/Yn/WN
UrTVMbzRxhc7Fjr/olnD4Q87ap/qLnjWao1oOOUJr1no/uuKTKqWd1b3RCYX4RWO
vr0XqsiyWrrrc1C4W6EOwGm/HLu2YQy0BdxNcfSeysF8XHAa8GYITsXCWkASF0Ee
sUT7oXTusxn3V/TzSkfpF5h605YmwRqRH6PZU2JMLnOUEuOfewjhTMdViLzpkJYT
oDVRPz/wFALbMfyN5rHT0Ajk7HDgYNwT4pdkards2nvjUawK2A2J1H1hxBswHXp6
p5hNoKVO/w/cL+wRaYRmZzEi4In2TXd7jOgNb1lVXsp4KomFGIDOHnOLajTC5u5a
ISqpkqUH/QshKlMjh/ZiZD66PKgxmOAQ3NPAbdRRS6qm7ydSU2ZMxh2V6eJb5J+M
+CzIDNFrVS36JorOjEmFHnCXSZm+liw268AurbOP0FmhCZwB6qIrc1JpckOhrB+D
4ZK87udtSjhOacoB8TgzhMUDv6stZAC9pfLhFTOMZ4RPwH57zqJzDvhsrkkLxJqg
wdBXG2/hobjxC8Yt9MJPKSg1mcnNHcojLFycHr2BJbLowwaM1pYrPBeWCymZBGN+
l2Mw0Rc+Ek/vIfGuUAsfPVOhNI/vAny4MEtmbtq9rRO+GmeRxbdCHWP5Juf6ec3P
W7jiYjClImQNl3ik7930tg4nhh+/EGyuqHW6VylZx/Gpyn37B49G3Cmd56bABgJ6
PgMYQ1XOxKP/1Q9063uncse93gXoTDqSrP7QsXUnwcntt6HU+H+PfZZVZlAhyGyb
UCkYhO3Y/RvX7uCt3NrIDbGCzxKyriquDvaRp9ZKiZdbX7P2zf4LorpGdPPRyZH1
zqSmTq/L4+e/e3MHkZ497tdkH4zX3GI8h26FDaSPuQ0eAk6iud5I3kLBPHE32l2d
Wim7AQvsr/a68PuVkCC33qb/ol8PJRzwi5z3Ash/0+plyrBCCc1NTCGGJPlXGla5
YzEzvfFViF0zWcYUduUVpBo+cgKIw+u5HV5h1Z5pVQFyz8/YDgsgXeYX991m4CBF
knyxixBhknoR3R2ZACePnCUgdJleY5vzky+9jHzjqHLqaD4/JHk398vIIeoOtIfo
j0chWBFVvWaQoBWat5LEHiWPyo6e6TyBF+ha4hyiUdW+yoo6AQAywneisy6tJk3e
JXQJx9a/zhucntuVHTqqENZkRfwP6SwjKcMcI4TPJKbSXc34QlMBYoTAyb6OEVOD
ynVhLjLKpPe8fuWRMpBxRw5usCs5BESblGs+ulgftc+atz3qejYq48bqhH3ZuRUK
FmcPKc2OioRjqJf+wwl0ngd4fCIhlcWqkKs+aVom0EhLm2jYWxvMOUl+RM5iXcur
2zK02seyh+zLnnZSMJIf/1QKPVJjg+bxATPSpntD7jvI22K/6O5j/Ecjq4iSZN5X
2H1wsrv2RfnT6xSOs1Of8U53npZh1OuUmWB6BP2ebYqRESGqEGQOKcRW3Zuh9w46
qZyKpTKh5FqWYtNfDF+3KsRjcGS6TAPeFJOO40mvR37E6fXtJaz9RTgIeTW/BNfp
gy3p0IEMn9Axga2wJ5osCfJ0btbyYzxyL/Ocx86zhwUqZ8FREP8dBRHKQNsnW+pd
LoNZA9KhPfTkEBbHprKCefktY0cxiFcTU5/MqA0dhwsHdmB4022WMDM/dl3Ol7r8
FwDZgbzNPfhfX6SMD0BQrvtETlZsh6ezb3gaKcFEBst9nSsNGJ4uUfCNd5C84WDa
ypFdi4ogXUZlhNY1uUbL3tlQh727yYJeGLSSAu+lwZ87NrGw7DzbyH0kDU3UTZei
0zawlSofZCrDlsve2Qi91Fs6jWQritzmxWNThf/G4qQTGjyiv1ynCyLJGbrqVON8
SsvZjadBO0QFWxhS7EHdTYp1DSs+ap3LVQVd0JbcXoinB3VnZ3QXiFr7Kpa7gpeF
gIwsZx3YpbMTFG59o/25NbvrgVfAwlC+0OVQqUq2etbm5r/fh49olskppmYUpbkP
kjy+muxcnPnEBwzgPCSpFvV63KIYN9UGtk3zCLcpopcXMpLic2P13bqomOO/0JoI
T3OtOU4CE/QlAOMrK52uOiCnwO0ocgid225nkPcTzPEnx1H1U5Vapenbx83c0Hfm
CKRa/PZlMK/PaZCw3GCRNVecymq1X3k37eUqYW4T0XwxN7xW6dOp5HqQDnHv+amP
3Sr2sxX/3hudMdxnCggX3VvxAGgOaNZTE2+ml7uMmgn+wULQNF3fOh0c8tgDp2Nz
ZO6kiMYQg/50Pyh5CC1HqP/RUOc8tOZX0fyaqTrYwmRYN2NNwlHlzdfgCQRe2W93
Zg8Vb3Aj94FeWNY+Ah8jGgCIuO2A9pZ+Ae4xXJzg65DOZbC2e/4JKluTmFQHrCVX
spqghBXmggHCv2IRLZkg+xBWjSbMKCR53bza8Kogif5iar81iwueIs/+bzqmfpdA
k62KWbfEYyI48uYYji/EyjLP8bysHuNnKCttKSYdRUDepcH2QTcNOuMeeHZiP0zf
ffQLgFn8W78PU0i/pm1Na0pCQvLjdYLup1UBtuQclnE/a5rxTPgVgRJTi7LEV6z2
w16ir3oeu9uEiBZcuAd9EXn89l+5dWs0f4dOENT5v1jDtNuNLa0pxCy3fPbkEsNd
wWGCzIO/5MkWDMWZW6avQFNT76rkVgnR8yIybs34iIL4T/Qj5lyqG+yYfCvXxvWt
J0f9V85LwHNrwwbjebleR3IR4NRUTdUQcNl8LkGFBeYiqYLJjtNFcJjeUlwIQF0L
hNvB9U46TOmxHjRbQqlUEFmh2tUZYD0G5Mpq+9n+XXczdte0MzKEH4Bo7/H3CAho
WnF716LxLgxrjeHFAE8x56fkGO8jL4A2EPIWE9WsCxOqT8oNegXjBkrOgeI0JOD2
4YgUzqfUPuiivSXSLd1oMc2k2tW8F7KUPBkKYE3NztRPOiras6Ga/gyRtWsZSLoq
PraAWzd1ouN7fZY1sqIgTkPZBzHqssqhLiMS7df9T7iITio72QaAvHvuzkOB7n/o
ytPlUUj48LK6KibnLvX8xMzGZvvygB43u5JZEM2lrTumokyGSaTT6e2GJDo2D44K
NvqPvrLTKlEddXBW4zTHP1gqtfS36/IEWdx+mGeGvZj+4g7QBQCfMy3SzA8aLogj
k/M+q9LG/bor3EJmLqoWAZ/2jsR89BJCB+9TIYTXUI2vqPSeLumyA4aDggInPj2+
sm3PFzXxNw8BcKy09penlWQFvV8cnpq9QFJPAyB9Ow+ZE/T5WORizTG07mqcRO1X
+A+DJAROQ3/dJEkQRh/HPzF/+4qI56zAF9JWnOJgOJbU+iXAf4BbdBVZz06bSVXO
RgKZKCoGqLwljnyb78ctBHbbOCPexxBl/NZfjhUDW/brNGp6SYmeYsnA3hJzwIx2
CKY4rS/DZEGEO5F4O4NZ/+n2x3HAsxI0wJKgywg3X5q/Se8pSZOJdKxvZqKw/et7
DLrfJS56KuRRSdIgDAaYyiYKW80+47Tyqh320ws/BrZM68yBL6c/terwwynHVMKx
rdHocfADADp7M264xtzjGp8jIpoaaYsow41No1RxlFYrlk+TJk6GMJ352UelFia/
gaYoy3TBVy/T5KhZsaCOHvPy9D5NDjJ9k9rRByF/HDxDI7BM7rRaU2fmM74Emm61
TcpOa0/6eJnXyX0g14fh507lSi9/nSdNANhHqXntaQ9nvP8sjgDwHc5oXpGbxvHs
+3VuYFTzx+iNOntITM7qbnFXtaxHaaRQkYIhECrpIy3k5eLU6GxB4Q1eu4RMDPWm
MOsBCbpnJFo1JxixAnC1mxlb6OYFx8czghQ1J9p4y761isF7+VtiS0s9IGQOb3QP
HX9IfT+98FYDkjWq06xxkMZ/lOzFFNNUPzcBeGqIpx3eelZUHPBoIyhoRiXxAlg5
G9IdQbwpZsTT9tGxSYsQSOV/B8KcpbzVYG6C4VdUIc4NJ7Hl8fPM70zqsGaMlDA3
MRjA7mjohbgSh6xnl8JnDPy8yglJvPWc7KM9VbmDnUZr0BwNTdEBzB2uaztIuW8f
oWVcuCeDUsUnG3yAUTGUL6IQFOK38VkfhctBWfEPDz/Mmyrp5+MPR+HySdQuDVVI
vwgGq6mnd5ixx2+Zz/Ru7i/+qK6OlITLk92FlZ3dwW9ah8HINmnfivpH5XI53OU3
lVk8CPL0e22QU/RatVIyucAvH8zcIbPCLqT1nfw47WE0ibsCQYbzFUyfzD1m+lRu
riz4QKqUJr/qdy8K9pLGR9c96hz9plp68x9t9dL7r6cE4gc+hyMManzBQ5YnaQM1
8tgrfHgTb1HN7uk3clcx7s/2ijS52LZT23BvoBDGmOksvYVKv/aQ1F8irtgiJd24
FuLezC4MZN7ohzbL8DN9vf8c69wWUXOtUP7oW8lqwS0zt+BnfUSk/isMfTvL/Kpv
v2ra9PtzqBculL7OpCB3AEGK0UNFQUrbis+Fv+UAZjdbD6oYe8+NCiISoqK+AZr+
mWld+UNQ+pbVvH3rt6SCs8BDOHRPhoR0toOHacI0ug0yx0XcBtdRgKlj2bT1UXXe
0xUd6/FcbZ6RzsllAIYyK8p3tk+DStssDOQlHzQxZcFu3GlhydttHwcBL9ms5LTI
FvwCz9LojyHbSU6u4Wi2qoA0FMFzD94EezOOAX1pQPcJhgq+6luPJCoqTGnn9zdX
/YYuqkoDXMKDUOAPNDI0C2VaDChPjtKcYM3y6xXcWbo08bul9t8WE8UAFCHcmyry
N4/X/am8txxueW35FpIXpxuW4FqzoqwuvzuR6A7dxkXuDvgSJBXmGuOuJd6yJGuB
+6X1NP1zg4zTJG9bPG4wOi+yG93DfWod7Yk16k/4Zzt4ByB4lWiiI+igecjoHfkA
bN/zdMxVKslTjplchBa6vIUDecUHnhfYfjjIL9VjkVX41G7rnZQh1S/qrvM0Gw4f
u0eGPJXJik6LrtGKwl/k1aBmnxWOdQmencqbmWJys2J8Rrtop1MA9ApVURFp9+ut
d2EwtdxcFO4iMp3tYUfFk0Zk3+z64kGwpmhej5qAP0R6AM55pjXjX21id65Ipcn9
P/oEuBWuiI9gsXgaDKwPJfXvEoOjf2xGfkJa9EbrYCoMnf5vHr0IAfxhp1RQey3s
hMOuMnb0dG9VbLY3j4c08Vk7i8PA1ErSZwdFNGBeFahQDKXhJao7mZurEf67HaAV
ZBm2XTrfanOeL/2HkY8mbK8dpOzof3ve+941Ujm/9dcqia3qcHGT7HHwl7kHIUq4
dkztIwiFxson11ARLGx00Z/g8DSyhhLzPPCdypxbxWHNgCeGbucWDpabjMs7ySYj
/uDwGdgvDGNZFlDRr9Px6DGz6wXBUSnnUMAYPJeFIU7Z2sfxK5ihD8aVaGcDkq2l
rlQYSki5J7P6GFV2Mb2+YRoys20fkEPkEdEmj8rNGduYk1VKfW1wIGJKOSCJmchH
OBFgCXWcWI+aG00rBHh/lExBruQ3hiIdwER/TsFlKQXMgJZ9X7M5QoVFAKznCpp6
09h03ldwkg8K3QeNq4y4MODLEAZ/08C0qY5Q3lzX5WouV/pymyWpxbOkmGGk7Oa2
Vgq/rowmEZycQRP5APvCtd99wSdZeFP7iRDljich1Gep0OBCjO2gZRKHGZGF1NuF
Wkc97wQ5BVaqrJH4kLE1PDdZEzFCETSuC098X0Shql+6A9yaaG23kMcxWehF5ydn
8xeeOWPXKD1nom3DNUD00pK2y7VQE1FIIMszPi6zW8FJPvZURZaKMlnkHciDVZds
vgxYWjk5imb63eOTj8H0uyPBuwhWM9KDjICX10IAPYQ763g7gwKCIZl1Ks9F2rEI
gH/QV9OHYrOIEanYDYTfsL6qAckSgu6Rr+WQVqEyDrUVA+HT8dGJ5UTrRwHzkV5b
U65713fqybxftoMQzoiCzp5Z+xAsHCb1w32JR92z6gpZVViJ6f12nQzM88hwngox
w/4O1jcFjIojPQBlsq8M0zeLnsDmjS/S5OY5XXK1x5TPrm/nypkZu4RuugfqAOGK
HzEnrv3RG+hiYSJHo+N9Sdbx369I0A0ZNPZjyEdGYHHy+VKxqDosX2h4TuaUCgjf
h/1yoTWzKrYjiFvMXZ5deMBSDOGVaNuNXXQ89N5XTIRjpB97vDLjIjjoh9Ls9DQ5
TF0vQt8X0dvt0gs8r4Y/jARW3etUPnIDK2RCR4XrgdSZeGpIoH+wA9KyQXyQfnQi
tQobag18khAU4EQL/f3yNfgukA2lvV66EyZKXFlDP3ORMDrjMBg+sYniJnzXBKUM
PdMoDWM7TU+3PnpxocibFgYlFMkKTLW2Td0lBiM6WXnnNgR663CLdcIhZcZXh+f1
y7sejbfzp1rni0CDEdy5KwTlXouQZzgWADsUod0PnmLNh5FR4Bb/DjvzIFbihdgU
SOnWDRpNodQVZ2RtsOoRIosHhHpkcZZvsjMxO5EBZ9kTUc6TjxwuHUAqllarlLru
yXbGVvoawCiSiVfHSXaW/JjBc3LsDDja9P12wlmSGXKKXhdIzvzX72nioUsJ67Z6
wd8iV6LLOrfF9fJ/kny0iwWTBHVQ0fsbXuu9N8YeNzRtl3E1gdbonGtn+BUmvroo
DwIfd+1YIh2ljnQMMmc39twvAsY2rNc5PSfEYrH9nNpE0xiZtrfTqKJ2qEFlyTsT
ktzvHjegiJE6tfWQOrCroRM+UFlDZBqvchAUvXtJ1S0KHmVegn/r0ZnOlUTMQ+6C
JYHctUlUxfowNxlHKlznw5ZvIgwsHNzSekgg4Yn7b/uasj7jFviAAruNt+ieWRFi
naikxeYwF0Umub1C284CvhdsLPfvN7lXbutJitpSiQY8XVTyu95KRJjNkj9pf2Bo
UGRvYyUP1yGgxQsfKISxMHwFCSkosSsstHmzr8ptbepQxMewBKDcTLMLsxNjt4va
CY++4lu5SHmNFfpSpEoAK9z5i+Wey6neV7T3VGhfvfK/FdLZoJAwMnHcnTMtlj3+
9+DTAB3Bz5XCv0R9EF4rGan3k3nfKzwU18UKCy8QWudDkXDCp9Rm+16a0koDEuGn
+mFSl4GU4Dq1z56rAvGncwgty+iNXMb0s2lZcGssB+IuV2N3mT+is5ofXrYu13ut
p54nnlyODcjTqshE9EqMbtarknJ/CoDg6HiAmbr7pibFHn/aAYlKttarWk74PMg0
ZRKHAZP2+AzQgcaJgiSAZACWQIXKiX6UetcG/4e5Kz7s3yfSkZtKqyCBwFzvAcnu
Xj+Mm2GGqDKkAHfuLwh0wHVmUlxWAE8XwVHVY+Vdp27KLZYgHRzoo6VwYSJrWku3
SGWnbPHmlqM+jDzBkGkU+2u9oVv++YT+wrbsHLpeYxSkuTVCM2bsuzBLxzuLVNyH
nr9qxz41OUnwo1yZtdoKYAXhH+s14IvpQVH8QiTz2cAkX9kCkvlZ4ooj9eyVUD+V
yd+4Mre/b1z1gzGOM+y6tyEtCUgvFMOO72H+wgHPwVbtX/6+IF/dcRlbAvq7JwcM
CHm5dHfXEaI2ibked9gkkI5TjXPw31INtwr3wjTtLXO2n6R0gLuRohqBUUrv8sgO
hV0Gh73DeML74zZdSpaS2zjPvxl5NTP93t+SaIkPrm0Jc8PUKKB9PRkX9NaYiVy1
1QNYMMC5s6zJ+8JPz2U/Qt9/BAlTcXzzgvMMBgSHNzMNr8wkj4/EbApXBzyurxRp
sqa3XxYu7LCPChpPI1plgo/C+HH091Mxci1FZeU34TRCEDI0EGOTryfahpjg4kBn
akRhGdNRG8CKK3sz5C3ijf+OdByNc0/0ROFL9lqxL0GbPrMimTvx35aliFJyJpzm
EPJTmuMKkoa2jEhhei8ovuvOOwAU8d8UiZU5Kilxsp794wBFCzefLZFYuBvhUvMg
E9SGNrX4Dch5M1uuHiyVsmOu5Rfk/Wea1uObgdTD6iANut9gS1JjV6c08zUVrqFx
6alLYyv5xa9IyjnLYbrshOyByJ5HvX8iGLTVoVwx1uaHM/XmlE7388Md5+XvFyp8
0/V38PyoJUzKU1xpeN+H3PHEHCN5+bi0iayjFrpL4JI4FEehqqjwm5TxmDSSQDBI
NZx7rlMSPC82j5pDke2Iefzusd1Ndg1MlacW+kxORJj2ASWKJ13OqwP0ra0WCE8x
TWsblofCn+nGHD7PJZdluLJaR3Sa9+7m0UdJICovrOcbuzOFY+TXWhuiSl4ZJhQ1
ZUdShtteZoa7SaKJr7PSdIkvVGIVMXLNzl1zclUUy/SiVfpm2WIDVWXI6ouxO8UV
02soMNHjr7N/rRgQXQMq8YjjrjfFl6hOtDdEYiKVL9Aay+JimKzuS9ru715tG3mS
/uOmzbxuGUa8N4lEMbavxNbGGPjr9g5NQk70Q9FT9N36+aZXbp4UvpQm3iLC9y4x
wXtZs2JacqcgdeXr86bEcWKagCgcSIez/zcBMhu+7hxeOSmZ/D8DjSJL6b8d+gtP
vT6g7U85eFhBa4BZqLujiz480PEk1TNPY41IZC+y7F2/ZkTK6w8RWy6me9kPvpQM
qpzpKis5lq9PBsxO6JmQiKY2maa/s0luq3uxv8f/+xC7JNtKOWn/gNYr3eECIS+n
GbrzBwdAsSuqWXaPajY7esIk6/2LqEkE5NZO5Xqp3iWSITXiXFpbtMkfRrdsRzf5
f+DyvNQ8tlEYFQTqVRswVZfnjI5v79X9sUK+YSrVdfItMdGcjKtKSeQ3r/hmqJ1q
1sNbzMmAwJ4oy0SJXJqRGrFtwPhQpRBCsSmgs8Tr7WWHOdHhan53RqA+h1Kxj7Oj
aEKvg+A6poKCLi4TrvLTK0rpeI3s6gcxpksUFBLHn2747eRyVqX8VkkDKVdIYq63
81mqYbc8SG7O7mQ6T0QQf+f1DZTr5FBWKq4je7mU+PCO47Wh9XysSGX5jQQupMeA
DSz3xmAnH91X9KpbVRo/u26x+wrT8vQUPkU+39qVoS4STGDj5P3NPk1hJ9TRXVIF
UcKHysvtuPSKox/UDQoHu7+tw/JV0ysMj9vBOioZpkJivcJBS/T7Nyv8m9QVtX3y
OMfdmsfzl29kA8/O1egURTadCNp6ZNF178n2ThoXT5UY4knErfe3rJqDD9mZUEPF
rbKxMLn3rwPLmVsO/gPeZIzGNS8ed3kFpgIIgP4itzEUxFktqJRz78fjKzo3eKi1
wzGh3CvPzyLU7xojh4LmDuOjhmqjqsplm9rCEiqjQnpgVlLcZw8ztEL6crznImHF
g5mQesyjYZ2CaA/VfpityUnJnzpqdpIUSvph6tTPMtpG6NKEhnO98ehqQLGP5mEM
Dt8xFDskbDEhDvbT0lEfiDGwpQ29wr7Rp7FN5v2ABexBEgR9yGoA7P1YVGqauMbE
/qHWVaEEQCTIYnXBDxm9gexDQnUwO+oDChTkCNLRNLi0QyIH1AQSNoZFxYklilDB
l/mxaW/oNsMgqTTX8WEt1q6I7NIeaLrWeoznrRX9U+fCi43fkKKytoUs5O3z0/cp
sjEain6hLXoGDBO4ahtP1C6pp/n+FLLSUCMsXRIs6YxDs1MOYzhFIbQ0gsZ9VAT9
hZDlYPjNzIPmM0gEZaeRbRvHSyI4FhqMla3JTdQ3RO/6FKoOrTtdkEzvthHrKwQ9
1aBDTJN/7cRU1woU2oSeaY5MB5rjhyPraz+Ce5BWQknU/3XHWwPyHX2/Gn/ifyiI
Dm0dmAjvAgX91PRTBfXkgBYsBaQLPHlpFxRamR0q656ewn9M3TefSXxCWF9CaIxR
GxVJdT02amVkCKvaCm5tHm7lZKn6QOcEgk7gU+D8oXeoZIS58+zbkcmeKAP0aKL5
4YlgJzAIn5c93Hp5wM70nzHkK9mdzB+3QAaFyOtLkCNqeJUg9OsqRQ1e3+YS6XqE
htKxAxNLOrsM8pyrU+mmJYxxV+0cOosROL5ttIcy2OZbYcOUjx2Awar4T+4x2Ark
PCzmyMCQ5Dd60gt1dYtX8AWS1mBy4RG8ezxEc6V5WultQl6TGgUTbqjD77dbo559
xuhJTWstf1CLVNyR2G1Lzaqi1lIOKwqs58eEa7l6JR4fW9rIuPdcDq4KstyapFCG
i0r5oNTArgDezlWqjlYtUsTW1GH4w47LFdsl9EJJQYLsdcPQK6UiJfCC30aeyWht
cUS/2GxMa5ZgLod6eR6FHp8hFLl6sG4T7XfmjoQJsJsZPdGuSV2b/4DAK6QeGLqA
bybzjLDusVGpOBKVSnvW1Sw//V0jqWpO67/ltkztYwk3kMxwew5+mQ+Rw5LZ5tKl
q25EXfSd2BQDAb8Qre0dilXQCjMDr3YnQCaLDu1P+rt0bun7u+OMDt6R0rBcudm3
xOx4ft5blbmF/eEa3Pb4nhPFIijnvUXSqOguRTJQYbyN2yGf4LSwpzsESyPphexj
EESA3fDXxulWF3/meZl705S89p4twhiiV8ZsHhle5VEgGLTtC0lcH2UxwuJUuwCv
9ZrUIr/AuD4PhrNIuCOPq88l9XvOFV/rftVKLmsa2/5mIZQXGJxtpbVlr7L7DnTU
f4syJDayO7HhbV71yOzwMIFimZD1gRA3ijIYieLgoDrEwYR/bz865/oi7fEQNoOv
sX2UiiR6OrTNCBi4cq8E83JOOboA+UBvOrAliWt58p70n8F+PON8Sz8lEbyPzOF8
xDjlkohHzjXJLCKHSBj4T5CFgFiS/T+6a4QvUAtiX7QNlMQfuhR6YJIuafiV64fO
rKXR05lNegXJGH4iLBZ1Oze89a7ctk8WyrV11Aly2BKpPyNT20mx5hk35CIL7ntE
Dpzm4g7LwJYuXs07/R1Y2c1qkIsBcE/fJ8JQ+GgqNslZX2JOfxKpVya85ewt3IXJ
ePofMS8ygwk8Qx/nzVRysW7Acbzd6ouXMYVUTzfNtj+zcnK4Eglxp1kDtjiefZjM
SsbxXLwmrckNMRAxnhEOS1g+9XrgtzPxehafk7eun6QWO3rXA4pEPE+S1YRoDjRx
HmF87d8cVmihdaiYMHQDyQVQHFEtScTaBnwxoRfpKibNTTJ/QeLPBbDxAZWjvo6O
ZEjmge6G3BU05KJiaYEq7nGbVwAXhDZF+Pu17O7OdPIBAiZxzw+NS5LQKvQCPk3B
SwKOahJV1h9lRS+c/AMnj9M7Ksc3RRh1jjGhvUXRgAxRZBFIqNLzjljXqtHKcJYK
5TAey4qII2P4Zx0FnYktPXNZYKn5MvQxrs9mgxCdsKZ6YYelq0/sBtD3MukyzxIp
cZ4zz/fdsyEVroQA1rNd6DC/ojdHk25+JAHQRM1cvyxgDvxQrb4ngEX/WkfQ4e/E
2JliAT9BzekhBM1e/eu+RzyMi7rBewyyDyC8AxILk8trpCIjelXsE6Fv2BueEB5q
1vZQLIeo/jcnlrNNkZ2uVeDI6SM1OkBqBSNLTZHW2mxg2pdNGD1ixlCUMYqoveIi
BOxJL1s2Qn0g217SzYu7GeG2u1zCummkTpT6osgp1rHt85tVOpCmuuE8tDFe6/Vj
ENYrz0N0n2H+2Dg/hCbv/zMLHBuk4AyzBYJHDkwPHPPNy0+I0Ng6O6adOzaB29lS
NH81oei8Guwsapb7WoamImP3ArJ0U3/mVmz888C1eOOd//WX4D3kOU/ErWfSeTQb
NXtFRzPbCUUE6InvrzU12XEdQJoyrOv8io7Ni1J8Jn6etgHsKBs4U/wctso9qpFf
Y73aTazYNRU7/XFuu/AYn3mfMDLdgxOYUZ3hxGrAbHUMuw4BX4PY6pK77J1llQLL
Gt2kuLUmnq5W7qGdV7DVU4M3rI3NFU6o2qEK+K6dFBbYS1TGt+/d7DWRBS2RUvGg
rIlJeSObPE0wFDqFIObxn3/UIIWvn1uVJScGR7HEGLyHdoq2cy8r9Rs89Flkwsg0
IkxNYmcMLcJ+li2wkeWctMUq/kfgL/ZwI0brnCeLEXejjhzL1T4rIsRapNR+OoJC
qvKB8OOMmskalc5lB9zM5mqnBO4tRNm0HTW3mhFo80L3JrKmNpYb3GOZqgWxSI8G
AUShV8LbaQ8Ofrv2tybAajPxGFRHfZ8n1PJnR0JfWZW6fUAiCSyH04GTFwevEbfy
1ySRFkwj/BnMghldaMKd36XNO+yMzCNS/fqo9OXXmcspUNv/CPlq0C/gyKi1GJRm
HeSHOMX9zaLRSVSuY1ButfcI8p9nn0Z1VN1pzPTcfls0/bvsvwWqCzfwGLns6cl/
coGHOIynOKbQE5d6PTCs5MZkIcceD0rKKipF11tEeWk6ZgGHIS2yXjF2rWQ4YBt4
mtDrsTcfcnrHzSf7QAWx9OXVJHCqQ05Ny/4hCtYRW5tihIJ0gGcxjk5d22tjqin/
CuCGr9Fo6vhdUcR9f89N7boimm1wJg5FYm2BelvOLDG8aETlHpHAhOQe2wXbCz75
9uo3cvF1Ks8LC0vo6zp8C5uRnwyXj7oQnpP7WUl2YjztrJ4L5mJ/gE2QTfMt6Vic
TK0ubRNV8wLMY+WDuz9KORqf5Mk0tjcLuhekO7w/InG4JlZo4S1qRL9BEyqoibf3
8851wzd9gDcu45zz1Q73X/P3/SwdN5lpBK8soMOzxueUEmYojpDYmw3BIQL1Bav3
+a4FLic5yq8CRSiIFcviU6A5J64FNjzO1DD8koRKxmzSCKEU7pm50BYGrnXrwMIu
Xb9uRuN6KUqbfDe/rv5D8aU1UcHkoNW7SqV2w581ufLFoSp8DbP5KgHtk4q2NJsR
5y1r9BMB65i1dxx1jwl0oUSbkrJHjNFOl6bMUSVSDu7WkmnF670Uq2BHnfWygQlZ
RQ78jRHcXHEUI6ghg94WS4n6Y7giuzHxxpW7z3o6JT0A0dnojs50ecWJCCbskL3O
N1U9CX3ckC6I0Y5MJO/t4cMoLCzpl4zfWuXfJSnY0U++BBTn2komubHtTWp04zzF
89/b7KBQVdHLBg2QNl0JEHz0Bb3tsQGIalUwtoWFqgIT1IT7LP/UiyFLg1LrjSD2
StCg4WKW+ssCujbEpNmF86qBAaFv7umFfqcEPDIjF850HnBCns12Xu+TPPt4f8EW
Iu7ktoXphBZGw6vOZb4Oh6qZG/UoWZ2uR7HGNGAaKWGmQuWZ/JOE+vNwDRTsfovF
R+WCTjnoM1MmOxrIYfEqnT6oSSxhd2xCZLii1eqWMwiwX3YGnHviMLnYir1QkT1u
7kQ49oH3Jw5ivu5ckRWW4A+Ik1f7cx+ErUMaIZWdcWqdG3YyshS/hpZLLKCjsAKR
1kJay2RgbFQBKuqGBE9c+cssLk15tN0DAt74m5AhTBlQigqOsFy8oQbGzeOSg95g
fzj/HQ0AQzbnYaHUvw5Phf2cNgBHj49kjVHKvpUbqXPT0JRp7Xrj6g1pGu2mRVkx
4qJR2fNyGV3pAeGhKclcvCHTI2RoUFa0bMQWDM1v/Xkv7bizRkEVZsbAjEYKl0bD
OwZkovV8gbgYxzOJvaTqXmJitFLaFDX7bgEJrqLuWKhlI/hjx2JKcbX9MwXSos6N
0Jn6ID3iOb9KYGqi5kbt95a6RiUNgKN9a4JUWKqqpdR4Iy7hs79tOJguVOd8P3HP
bAR0fv+AfhFMLc+b76+iC7WMXYWn6xtHKedZOojKyMBUIC/MQX2yyJw07M3nPdRh
5lB794r3cfM17qOCz8iIwkWqtbg/mtryxenOavaU7m8Y4f8G1aeQyzzuaj7SCu1A
KZiyOiqWsLR5QxZJwhdAb2D++ndYKN20fAa8IaRjyiW5ayG8gAQdKpzGdaYe4By2
Jgb3ifE9YIPNedTOtDw3FjrX0orWdnopOCi4nAil6bSAl+wBU5K/7ZKFwk/OdSAt
fHf55vCQHpNOejNo/1VKxDlxZIvx5ClaJ1P209imkZpda9hONwxJt4G2txjfC3V4
azA97cuHf4OsRZGFoEEYqxZaMbj1rqQ9rph7Eq7PZWX3Z29ji0qOY8TZDjj3nygp
wqWIP3QFpUIFFbWzimCx9cn7D6YZy882lZYf8TNxKYSTc/8uhRxg/+vTyrwlSyaE
YAeXeUY3m7OnqKpgo7aF8oA4+yay+3ADODkcOBwT10x5Fapl0VlzYLD8JT5PcOGM
BGsVMKDoFxgJq0y30SJLSWpfl+o0uezYgYtsD4XUBHaS88Ba+mDmK/DV9HUEf0bd
dWqxpep4VQWki+8bOT4mbByI970GBgzk7DATb33dZJzgCwpOy3UTuhoTHAK+Ljgx
CFIru2EY6CM6GLJNwq7zTjbx/pZYoT4ggUxasVDeQM0i5v4m4lfgNO0XBtipiVRD
UvlbhTCMHxIbSaOwZcR/RQyiFo08rVLJAqAlsSQNALhXwnc7vygI/NWsXYlY2ACF
lD4pytv1rZee34FXnkivMcM1eveoi6UweLHdniMY5GSiVXSADwETIcAz1kd+oltx
hdg6pKaoh0o9sUO+83vIpC4ccjyWTMwxzW8Q3Z1xTMcojpi+h5YciebTjG7C7XzR
giwD3A7JlTCXU2fa1+/RvZZylD2cANLVUWejUE5V1TPpifjiH5od0TIjtMlwb6E6
07JqmvdfBS7Nl5t2S/QiRY6mP+jKS032EWTWK2zi3pU7j8TDQ96iG9yFIYy69Jtc
RAHodaPmL1HHaQKTz4viSviRThmMlzY64yb2viHV3ezr44Je+3dXAEGc62BooBtH
SWg2rXFgKMVZBuwigyKxQwEALrZPQ+CgaElXs017OtRpxGzl+HN06MDIpBD/mhKr
WP2JRyAhLduqWG2gwPo8X37+ERdCCzipu8xTDZF2O36thqy6C1qwbXUy1G+6WnXM
l8IGLsE1aBUMOIxGHKY6/UlF9JW6jbELMfMX00gQUOeqs3YXJUswdTZhR9tb3i5V
CTKVlsW81VQW+q4Xo/+RHV14JDfOv2w1SK3P5Q9kEetCefheK9fzK9aOvbbQd7QT
xlBLETGqP9BUhok5lu+ooH56Hx59dTQpSxTeB3KbSWo3vuWVnc4EMzA1ZIexm81E
j0FIo6PNmp0X2f11mIpqHsT/FqD9W30OIqUHAWp4MXwzlKHaa8wwB1iEjJvUxxIt
eivS3X+YZ3xPSrfcPvqg8m4yxy9XasPF3rb8MfWOq1j2BgA+CgACJazThMIWF/B3
vA7ifIpAx/TJZmVOZmYHpC5zCxJE4H2Py8WGU9K9mBYT1v0FS3SCTHUAWdOfSSQs
2wS6nrj0Nvl3u2B0oX1pcHlN6rEbBu20KMA6xYAFNy6dM8cPBYFqkJmZjE1xuQAq
O+WnyAuxjJwzccitg976l1jVLeFG9rVwhgHhUSk9A7QLCjfqT3UA327iGabFWwzo
k0Ma64261/pdQc26jVmThGLifO8eI5hNPXPFNPWSGNTp62fTl2tUgB44+Hx/zAXE
JBZb+I8JVfn3ILRmmS5JhCMBAmKeQ4agKOKJALSoor9inbTJlQVtudd1UjcSUB0M
O9V6aS5qmtRheSdqCulKO8idFOuVOoUcxMRPWB391pBY6dMQCjzf6OX49G/RVTqS
0Xo78xu+FadBbuJNej/eSJPH/hZXrKyoymR9y7kcnctC57vyGWSyOTpLGaVs+55P
USKZFmMB80WAmgKrJhMQrzn8QSQr5a7tAx9qu8q1LTldfU/Jeq19zvLgpK0rHL0E
24zL/qaxhc2R1LLCmsuHyDKvKp2LUA3GV/6LspIOlRKK4X9PSKqyf2COeH+5TscG
wa3jX4YEbMfGu59a6uY2v3sAmpPvq7kdD52bFuvXTIk6foVep0EtKSglP5YnqTXL
UH1nwWRCzg95K1BALvjrs3tnsf+rI7uHr4fmptxQQ4ogKvAN3tVJsfbI20CIoH/c
FiMzy7PxjO8SwA5ZNKKTMbnSD9d2g3KXnc9zTAW8ll1Nmzxqp5yKj8gCbtus4d8d
zdR6p1XL0qLKqSxoxk8NUH/M7zxK29SNnHFiEajfdNZKzQq/9Mi00iVkzlTRlolV
5gVc8sWnUuoCBPXpmvzr3TBHNptFuj/xc7uB86tYeE+zygIchQsmz70vKd1oRuGs
AN/5RIdcMrn1lFQtiqtnTM4Tna1ThsHu86YF3lplKKHcr7uqzH+HYDiBBDDtTbxd
lf6oVKMbwEVoZfqV8k5e6m4m4sMLqLqM7BT3QJuZSwZHZu6abPXLvdh8zf+NPxJf
D+vmNsLfy5jZPvP/LgrzMkNpATxjdcRMEXMuiFTjJFIMi8BQv5a8qAmsAvH4IhJd
mvpLbDl4DDy7v1UQCSULWDd7pyzVylttE3gcjfjxtQoDlEaBVvOy7ebqs3QxFz1v
xkQLDJy8swZNua/1m7j/YTJnPNzRdD1hDxoP9hJsaNU+8JGHay3z6r0mxjBXC9sH
TT62FqNGrGUhHL2u/orcri1f7kBnBPluwjyynx06MikqEv/w8TIk/H5J8Z+26S6o
9dkMB86phlh9m5HABrOjPjPR65BEP3cIdX35uTsBAoOYRWeHbAxRXG15nvzqxL3+
pglo/Rtm1YpLcidzktcgHrN8IqGCi4EfHiJ5NNuOg1xl7mZPgdWLzkbHF6kA0/cM
O34AC5ZBW1cGqzBiddROUfM9dqEGEIDGBehR5dnoL/h05zWuHo8YwooBqDMz8pDG
ejlvb+F7GezDSZgY1sdzf4ZAO91HhfKXw0Fu1Di40sDJbCNDbEGW4DtxLxXpQ5kl
qK8ecrh8lXHIFAhTltyRfU82vYaIiUdObxPfPGArRY0IpsoiAsNQ4auhk3h3wgd5
3iB/VfIeH5wNV7jMTUmWTLtnJNDkGeolNFaJJo+nIi3NGxlm5GL3VQ0k4rmGpmmk
pkuy5lDH+9YvIcrF1nu/0WxH/5rWMAmen/uq2fE1rR9Gwg4aId0pMjHh+nioBis1
OA00zr/kSpI6gK2GwQ43taeJbxCOkPNpkatoDrmv35Ahf8onZ+I6GX18gsuTD3PQ
/+wHaoGSL3SSOh6JeHOVKoEvGmEpMOPsDIwVax0sUNPHmdA0Ndx3HnVwFIaZ4vsH
RirzGxFz7s6Xj5HaA0/7M2Kz8BMAmjaPgxRByj+hxeSm43VrgQG8vRsSguKJGKnk
9dX7uZnJLL0Di9cxqb2rMVVOZeFMy+4l3OpzDQS/TmLl4kMwrrlfoMeJfvb+s+v4
MQnORyeuXYKuOfkbYWI5t/Ht6L7NOLMZh/5vhrUW/t26vIHHJUWwYcslRaJuSD7r
oFl3mpVy2qwCmMsmcJ46Hyf2u9sa9lbFOB5sNAt1gwUQAUqwSSd9urg+6Fcikh3y
uVqdwMjtLjl7sa5UzMjTi8y5nojOvf/H1MojT6p84qEOZXrPWQQivNnW5UFOAqMn
uhkftcml3t6Ow+hLHPf1cXlQvkROeKsJFSn1HuSIN1opt4VZm+aqjTwAdOosA/iQ
Jevctx0YDtSj+CnEoASm4fC6PRbjKiBoF5OzaZm0duvKd9F3crzBgCME4LDXE/jv
+DvLoIwKVcl+Z4d1cp9fYDdBKDMUb8a2crgc0RjIYlj9YjZvvM0mxQmtP2tFUeaN
mgWDG0TziI7vp26QCyGcBI95KvTsB7RMolfMXeG8YVDi+DrNheQ9QSfiZc2Inf4c
weiRJxcUjY1GS8mlIrWDTIyChW5Q4A3s/32O45jwpHx5mr9XopYprIX15y+x0IPe
dXEv3D+Wp76QzixZ0dRiO8h81oNqUtT8Ba1sLCarQ3vrJn0cEJglELO3KY7bQ5bU
SbPv+btGlEbDoCL1suaZnWS9eAJhIjMF7aba9iR1Z9qVGwECxPH7iEaNlwWyy5lo
5WsboLgC2GL3XgXi6Nn4U9whpfNlJn+vpkeKRViQS2339gPymj2QTi2sp8f8JoOH
xOxtNui/axVmVjX4oJrWwAxjQKyWlCud4fUQN4KS7mhk3uf2DnlSz3GUs67tJWjm
aGZm/B8rhAFTcnK/uY4MtSL0PTalGLVM0QOlMdYGHk5K/D4Pnq4isybarQY+DRYx
w+MCBWnai5EL9WBHRaChM6p1ED0JZBMI3akG93ZqUxEBhWKON/jeOAyhhU3D1QY/
F6EJU9zX8vvw2PaIhFTFu4rAGeCaSehMV0seV3qyPBNC6b/7ZJqjFH1COJub7Gwq
vuwjXItFrtZ+L7O8s5Z185TTFParfjR5rZUAxJ9V3lFx9NH4LIoSS2La8nMXK1o/
Fdu0GBSabdide268OFoRh4rh3O2szirzxN41nwcDcWf+RfSLyLzQsxsPXOXneXbD
zJ6pZm0pEkfL+nM4+Tl8xqTMtv5kUvH58gY80ECfnO1PCYqV6Oc1PrzSzVMXkIF4
zNLlCKOtKLAzdhlsI0w4xtqs+s4GzoszGfa0XItPoWEWRAR/DLS/Is6hF3L4mpB/
6jcdu+4thYMXd94zwg5nY0MGec9EBiXfrx8FGLicomIGM70IUntVBhUcY3ORla7I
U9hqtYbFnAmZRzl3okLCaGbODkOAVUNZnOqwkSGRgdHyGaEykPQNtuhSeulXBgjy
ilcZHhZZMDFp6vaZ/usvx4zSAYkobOURL6lhCF/wLSn/Bmyltedy2ew03wescI98
NqcK9hPNRCJf46rp/N98NZkFvnKSNUWkzzgJvrPYP4lg4q85N1n0LWxO8HKKvlOw
crk8ZHihHF2yddwKBsNkasclGskQWvqMiAe0fzrb85LN5b9FkGDVdZplQHQbQRuN
bDi5CBXhdpYJ4sDCmpZIdrchDyRu9N5xk2U3YKuweWD0n7AZNEh4UvbQIXxOEzbh
O0Ma08W4okySpJFrM4NxgVOEsHPctIvhr/UJJU3dAzAWGZB2XV7SI39jc6o2jNiY
XgArzMmhwEG6AB6nGLZhSRUbZWe+kkYq0RMBZyL7kP18M4Grr/b2BGJ6hO8NxuC8
BWD3RDUhAAAsJH8gcqqj7TK6wOZ2PtytVah5p0ltlam6Mf2pzrewXqr61qjlRm+w
wf5HDc0u9SShszKmy4al2XC0EaYIap4TpmrF5USTYKvUHT3iYEQPaeS3vzXrBDsX
jayxqt3us9suulCmbRZrrxNDBif5wxNjINgkasUQ6kcbsVKPYa6W0VmPOsZPlqpA
Ws2eNXAuVnhYhMhnBeG5IhPcCuEoCNLlYvf4YT5xsoRjtZnGS1jpcWRyZTbVzWhT
SaE5ITXsQHLBZk9cPiBrKRfbDYSRVlFm7glKY+3R5sJz9B6uK15wsPs4294KqGBu
4v5VaZq+juLxUfKU1uMAZQU/GJRo2ggRvI3zFvWGJptxeE7iy6zEX5n60ujC5MJD
vqL6QaVIZ8XvHkhMjqn8KSAyMfRUd/Uxe+HCW1hWI+MdtIxG5VdPvKKDIYCq+SEY
tlkSErm24tORfBTBwN629y2oDDHWVn8qqWUD61D43Vn2kF4FQe6GOZr0a2HDo+0p
MvkiRHySvGV/CYSWqQqSB/6HQPNOjP6ZYSbDNTTDZkMz3piBvzct0pxwiKgtnxA+
G6dDeNzwAyrFiqdeoQWebP93qJEH5HWhl1Cys8yxyiq8m8l0G2jR72bjiyzYyi9f
Yh8Qg0IjHvV6BY92TgnZJzkgqJO9/7fs430u6ldQsNQltU3DeFKTq5RgaKDNSyZF
8Y/3jLEs39UazJ0FInxJhpo8OOoRZwULAmKuJx0v5HnJWdaN/gj47NB+LnXHeCZq
wWLiO39CnED7K2gpq0llR8m7wmFXLkPVj9gfVX2fk7rCQBgKlgFT4ps1iNjHfa7l
qJgcY/9zCKY7n2SRnMvkAqj5VGAKgPzKjQ3XSXC4Dz7Py6IdjgGAyqt41dGWPDFx
YN7cymxtCmWT3WiZ/p7TnT8oMmoBoJ1l04iAGWOV9sF6h4z5eeAR7EmRetxifjlb
6tbKboxG1fvUoLH0CbyDIw5guKI+e4pfUccP/ZF+fC6RTo7y4NabfQ0FSRVZTKSO
nYAr/HzzyVysY3tgVGZkVMbhM+XNwXur6dEf7139l4/f+vsXDBfcYFfQR+XIZI79
6Lgg3K0gQct+7VEA2VXfBwmrXz+Qs2GSp9akz0Nw2OpchbawPGEck358iL/fNbgR
yyadcwF57TwWwszb+z3n8wYuaGczJJMqwQnhsbhu5Cb/Vq0KmqVCJoAhk+1gFJaZ
JeHbWixanNdYQFJ41H+jCp+hnPBaCNIBgAsaDgZ1BUTNpHZkB2xD35tdZ0zHbr/y
1/fo76UARXGGlJYxrRkWuE39OlC4A6CUASo5pG07XjJBK9p0WC/L7bxLFFEPDS/E
KM4YavzND7UBMmfHfA01jadYOWjEntC2rLbqbh9/TdbNfnXaGHjNLCChReWEe2Yk
ACsVJYSI3Urga/L8DOTvug7YCOlwPoC4MQLS6G3ZnH+nTiBj8USxG3xmSiqeA+cG
tevCki/IuJvS9KcarIjIDUYxpMbUdCeRd9gPtgP2mWdu594AfBfbpCj7xLE4Hp4P
MpgUP07/OziPdb3YKmC5s2xaxR9vBfakX8WGtdFgJqllYgxNtziIP9TnLuKORlK6
2sjS0nil8LtosoggMYlVXToWwMh9JRXFNZ+ep+nSSQA2T7CAG2I03ZyfelC2azDV
vg/Y1xCC70YV2Jnp+S93tJvHIeT+5Dgy0n3kpIl87lX+lBPiT2EqVvaWWkZhT4HT
rEcc/clldXth4DXEWEmQdjoWakq3GMHGl4tOkv0GqPnIFujKqyFLfohxJH+zszaZ
+MdkWfSVibPTYw1e3tKSiShlvm1u8EGiy4VtZB1uSFywAhdiIIIJPZ4Ax2/qoPGi
Hk256cOJDQTDY4FRIzyBWL9zRuCJwDHCnAltnfaHL+bH1nYTlK5npCPSmIxaiENx
Gs0AYSSpPLQiESgK7VIvZUk6OzGmBC8oEdUhsGh/twPujZGcAzGkS9gcv7Av+8y3
PhEeVo0T08yKekmjDspilMLSXLVSQm3VWYOHNrYEOQU/4MC5DnlpZNdDmcg2Z0ZW
01JBEXaMvTcSgRvoIA9OlflcOH/ZN7VwPGuq/kSvE1ndUgmab9s6SFp9kShberWG
k3WyZWkP94gZUoaqCua3tWWE4yw2zgQpaZzICQbOLcFLWXPGZNB4fiwj1EXfhQ5n
H2Z710LyP0HyW5OAGvWwsKvkVpb64vcnXrFPeft6bqLpNItD7lvMT3UM+sh1Pys+
+hsYFmyAgUIKR96Pi5DI0Xywesvp46DIys2lPucEOTL11MiBmff5Y2KZxCTAtMrw
U5R3T8sjyckvH/NgxnHypTMkqxzdq/68VhfXP6YGaVziuoAcBUGw09lsNOYCuVCH
ACNCz/+JshuEfcSVLTsOwH86NnqjQynCnAYhXv2dHKfr0AqEuSHJcOkKa8EUXLIH
bLBsoekw4S5tTZSxMsxSAY5nWl0oKo3LEgLUttMSgLAt2XRiMWSMlce8e2v/edmt
W1mI4jue6Au4bfzVSTmXy5qYeVlOi0oH+m+1Qdlup1V5aRkGKWGy/Y3TDQYkFqPL
NiZI+IORxBQyOZsCIqcmEUniVBfjVEsQDRkIZTzmcRKjirW1hDMVVjzHwLP1sK55
tmU3uXapwB9oGxZIYusQXljC++dBqjL2yNNPOYvyEJJKY0wbwIYfwMTW1gwmaMgc
ikbnfEpMss/Pr2zO4ckZ7jG1FyjHKzDY4AUoSW6csBJgqPwedYxu2cqUeH5QKcig
qhGnuUrdPu1u7V6CHR0Q6SOds4vFlMbKBYiMmh6j6IYyXqZCIc+ZTRyTjtlCmNdA
WEl4ZBEVxx070LQtIA5Z6sWI4cO6MpM0rGtkXBkMmALuFhDV5kJXNTfDSUTm5oFR
9fPmBREQtIlHsHoEiv2N/i+lLqwq8f7gKXAl1tkDzxWam3UnAwJk4GRzQrSnbeKd
bF/kCtPBl3NpasRZxu39cb55hXKHrQcNayu5tlRAYfgQqd8u1srtZ/37bhK6TSNh
frVMI+eAl9ltHTk5m9NOVUfGsovzWUxo87klB3zy7rIEviTXzdVqm0BJg+G1I/NS
N2QxiUElw/7mxFFMhwxuj4GedVy57RmTLQI1YUZxSQ0sHo7XbnuzrG/RrkjqTr/z
+CLU7NBWwfERsmJCgn958xzUZmtPtyTl9GU35eSL7Zh8a+yfQPLuE+/ySVwemqW9
LtEL3V/Vf+uTS9EpxFE1oupGqzdYwzIUE59FBolijIEdUj56paddkykdTlx+ToKw
5MMIhYakhUeS1CgRgyEfasDkyjyScf3Jh/stqbhALWy0M1fN+i/erUu8+cloARwi
J1FHIbqg2XT55NcBvPrYczEj7nfEhXbLVQ024a7qZhQrMVD0SOZ+R5nGhhrsBDWS
Pp0H+nhFrVCzjIYtgBgU2TZ/yZwENvlu3vw6dsXbOsaUKtPx0Bic2MC+B7jOQKTR
qTW0iQsh1YY/jOnT13XSF8gmLlK46rxtEmsnqTCerEKueJEZsYOp8TG44Y7cMAeM
idaY9PuWBwnZjzeDKUEm1HMilJVQl3aeDq+UJ2ihQIp0glDpX8RCo5IsNEQ25gK3
MR4I8Hx5J0L+J+5PPNpHYjhFbtDfnhgpsKLHpRHoKQZlv/wRkCpVM+tLBpNnY8nk
Q7s/9xVehQq9YSx+UEr7tYo5zRfL3i/EvMRDrs5Vx92C2YzXuG/ck2fWr/ktU5pA
vX4SrAnhB5B9qXvmk5crFuWuk4tqxEeiQlzGlrHunON17kyAAzGz8k2IhtzOFGMT
tUSjvUc4r/lobv+2DX2Y+HxD7qq6Zi4r3VO7gjwpE1St+Hyu2wYBhZobeD0jv03Q
PB0uyosgZ5VQjUdHFHPh9Ws0etrdBAEwJbs6SylqUQQCELUFPG1fdRIwRoTFKn/y
m+vdcoNMcd4bYM8Wt3hA7Mx+f7DyOeDBMR1rKrgpBy0KgsjfBM36HY4iU2wJUlhC
hmvmWH+5h21JbC098kvDGFANqRRHF5Vx6LN9j2P769rhK8cgbC0WC0tT5biySLji
EPlKaeAtejV+G0WHQI/DgxIWpmqtMlNUKNAnuE51wV5i7Em+Vdwa+kT/5Nvw/orR
LpoIUtpWqnAFz5Isa+9Smost1OtUKeIe+7PrTflSkPMdMy82+/2j+kFlmtmYgr+j
I8W5cGrB/vSNuiAKZTxr6vpSuZC3wGGG2lJYPlbLqjWZoaezKWAISpMpeKToUJuY
RDLnarZ/2BqmCdA309UrVsaY6G7hepagShVU+mQjf5obEm1+Ntn7iZEJW8ZWpI7a
5HJD4joeoXjldLo+iCM8w6nSeI1xzU9BORCiiocFWTBmr5RzK1Iewfx5fJE7I/61
W+fcqFsave7zKcVgY77eL4T5MW6yCH+HGPjuO1sPpKKQh5+Cvb7FG7A3GepWEdOs
GmsNCQQTJOakn/pJ9SDrvPV0osq8vNG4zroodAGCHgPMhXxPEb76xEGj0S+JU+u1
93rEziypACv6YMwcxuKbeV97U6Qxi56iRV8MZUjUe/lNBfQo/qKTx+DBLagfOA+P
ILN3/HMGqgXnHGIVwKwxCHxpK3Hqu+QfAHNZ6szBZqJ2+uY7Pc3bizBik8M8GAfZ
BfueWj8c5bZC8OaPFqK+KhsxTAKNXrLxaFOMD+dOdSWyyJg5mltX7VXVfxsIIk2L
nubDVygm/DxmHDQkl2O/vYrTgICT6e0ibVM+CKpsQGknvEnFPuluBkoq0JbIbqzm
gNq5Po4xJqz3rSq8lsMQfAb+KHmWt6ZypV+MLfjVYaaIr2213sZf1sAi5Sh+UW87
cHxhcGSlKnSbNIQ8WnoEaT2dDyCBIQBoX2FdO5yRiZ5mP/1Lc/UPgeFbUIOkuWja
OcCSiQNOCfONA596M5CSdpyWi07R/ce8fKGWcKO/3w6hzC1rgtcGr961Q9kevkge
XlGL5/vyPnaRMeqgUsRVYcZXlmbDs2b8yBmyC2J1CDo5N0OXJYUOfreUfRUY0ybq
mtbimv3ETLe14nzZ3aBT46LwD+kVwVVjAPyUDUKWWFLKeoaUnSDs+7ay6tKR5S1Z
1/X+UI2SYtZ2tJ/w+KRG+HFftoyFyXeL+Y8yaYa8h8v1lVJBfUdJNh9wXczz6QcZ
M074yPNvF/UESz3+69wx9hL7q0c/BLKdk5yAg+VGVP4MF4JIHtigw8cr2S0X6sx9
p5ZhYh9hHslym1vsN4BXmgdLX0MDVpnqKzOIl2xyqYanXrSlcy7FOukym314jHKU
+GKqpSR4jIZf9DYdHqUgjVrRl3Q3B4BHVAjnylngBnbf8YDO42Scd9SXmWr+g73f
CdXetE6+MqR68rmZhuXWSWmYnjrS6w6bF0GYJXPzSpCybifzfveJO2evo5URvXKx
20et9pnVBueW6PivB06oJUqlHMg3yZ46ebGqzmNqpacZhEf+HCv7zlykPA9SLnT4
r8gt5FgzV7g2a4Ekrt8UaFRD0qxjMjpxh97+I126OB7Adfb1tfCgPk22c9nH7VEe
FPpWJ4vkuLtRMwTcq+/I6XpiwCtG5Rxsr0LaPr9H5zFqAJV+NqrFx4tUSD6kYZXj
gPTXUB0mCDubtRGUqO4JSlHav8mdklQ6TDvatJJ0BeOBWmkIK7Jx5cjDtuEJmNp6
6HBcMGYzEIJCBgDKBURRKYJSBW+7FErQiL8FHQtDW4f5XxQ7iLARqfn7YxSNiXU1
EE3C5RvtqQeEL+bo53vbNhv9sZGxy2/vrcEodU4yOxst3DXZ0WmmygFSNXJKP/BH
qngWGP5i+L7G+W+tz+261SuRoQ/FFGZgebUymryuLNKxBCXkjhY0JAnwaBGc2It6
1UPQRJG5PSSx8yqfAugO+iJLbE74bBbR+TRFAZOW26oJbLBikBJMyzyfDfcRPEvt
PzRH1HjaWJBTn2rpE/qxdJkCN9WnaXgc4frL1PSH3cH52QrFvcELayegnutqC11K
I2yOiexIajlmYtcPOSShKthssBdxOChEDdY1an2+e8rjqN2R98BvHg3wecpZyvsQ
D9sg4hm0oOluzSotG1ULIKKMZT/QBe3Gcb5LXNxoEyt7V5bZif7oWualS+XSm7u6
QJgQegSx11YmPWssC2bUUiljjONiYPS6uKUvnOXub4DTOP65Sj9ZiAgQMNDeivwy
ix4ImkXzUzIAJClv+yiAo7ETSer7690XmEqVP/55mgTXtCNQfxn5ebqbtH2y0bDU
7P32zofsawQpwHrxKBZvRsneiJ2rGDn1gYqq1t0p6IKHqx7YJBlkFZCZ6ZTcKTcT
9QKEU0+8aoJ6Zpvl6cl6KbMtu5rCSuoz8+aRy+MPu5IJlHSQsSIvPniUjt1QNcKx
9rBkgCTzuYMONCOwuRxIEuaadANjXn/OKsPWW1Ffo9A9sVPGuXYnJS6omourVU3t
9z0HAfHiEFV34gj7gZQsSZiD5Uw0J6vLTfLzXTUbx7QWj0dw0b6dulO6gTsd+Md5
buvBMwQgey2XgcNQwBHWGNPTUh0MTU7BQ52s17TH23TrfbAOdGzIw3b76RJ3zmkQ
iKUa/olfCdxE+BdDWdmf2CES5tX2JKVaMMA/7htgTDgSCq4Fd8ZKFbFM/xeYCXd+
VGWRvc1IZi0EOHKBrlzzGzOVUzytN1E2SdVdLpOXClGWH6IPkX2sSYJznHb+4GOF
gar5VzBIzctN7TzBNK5kVtBO8VoXwgn9SZ5Q3PKqIf55DzAU53jMadqacZ0VaBV9
61HNrE9ThFBVeN+nd7Pp1WoF7oXM4LPgprBUR2i7cV4//IqYEQbCwEifbyG0n7/3
wpQZD29fIHMpbO+Uz0Yz15eKX5mM8Gts8R6npwll2W0Xvz+AvS0iXTy5yq0uWUBm
V8yGY344cQ6rZImxW76VVaEoT9Pn4UMKtOOK7fJOKth2ihMXfEk1mEzVRB/9uayJ
o0VJYoOL2m8DhPlRsu1jKZ6O758rqL9eXV9lKOMfRzxm74PtIKCy0kYKfE7Cd9Oh
ujyI+r5NZDeSg3AgB6UbBrcR1dKhJ18UPH3RLd+IpOj/DC0oTWGl1Wyqqg4vjhFV
ud1MFdiykKkMKeX8ECn27S8ogrxEAk0SJR4KZpzeSmJ8J3JKuVXCJHNdo2ZU1Wj4
EcDPVY6xFAJk6/lkl0VeF6zHFibeeHrFE/suWXDeOGsZBXpvECZN0EXn8nf6BTMQ
wHN97eSd/55bxESDUBQKX/YKPaS5bB6vUTsjTSxT87sh+XmqNv2aQYE5CyYtiBr9
JL8TsnQF872Ewuk7GXBjdm1zMzlTyu5yaqD59zNPAfZLUuuVy40PTvE5jLWvgjtT
yaEhjYxM30HDsdMl8Sqp52wLuISCmTo6+Gu667V3GfXvNPLHaYMvEyIDw26D4+5v
4LqtXM+BCit9v507+yklTnIO1/jCJ4ILiJCdTMCnFPD6R3Kb/EPutib139m51KBh
TC9tg2vW4UG/1cu7RBBS3fTtlVpv/Cxt7tKVGQRuUb1KgifJqcCrtC4tCxHhSmRK
kbcA+QLSU3VCeyLFrl+5PFVo6aR6YXYn61yKuZUKgcbZ4qSEE8t0rowlpM4KRSQ3
OakIRJV80IB3ypwzxgJH+SqyfA5onMR/P4qGcO0+QRRgUZeThBgX9Y1QMgnfJ3A4
yX8hBrwNH5A8fh/MV4KH81h9x2c1Apfm8GhCtP2US9GwoknmyzQuGIR/gS/ifVkd
Xy9wWslaQCyFuRURB+uKaTdkSDixS94c+I1R15lK9QgZe5lk87LAtOP1qB6jYCRo
BXqVvuPE22h0wfeCrCzgOsS9Qq5Ikkwv2vC+Zz0U2RgaLQNWabl/P99Io+f5JtrJ
abFwYolOba8f6bSYjpw+8WgiOQL8bUhp7bqJG1lvno2v7/woNgC24tfupuF+PIN5
2iqeL5X1IyaRGNcm5+w8Nfn4WQky5jjRutHfWmxFpq3vLdnsRm5VV356bWcXsHgA
uEW7T6eraG6JhDdN9GPDD3OFHols0I5dNwDlZYLfERAJDGakVh2XqH2R9Mo/OTna
VyeSgM4Wf3mrTp9LARmLd6Kg4kL6lH3emtDw3wPswrKxIUUUDWKjDysGNtL7sCK0
UZFgcyr6lmlFFO4/KGCOFRPrr41aOWeSvTRd1ogBs+D9g/Jx9F198MvKm4AMZibx
G6RZYZa4/D4bhiL7gH7L0gNvgqofxpJp+jJapoQhnbZRJ+V9qgbmQ9j4eqrbzRVS
P/XLWwmrBOnseqshq9uyzjr3Pbg0f16x798Wsdqa6QprpNXs5NoSVw8Bgq5Mfz3q
Bf+pWP45/tnhlch7s+u3QSY8PGJ2bJz/Zx88BMpbdTHZxdajy70DsHxRit2Ca3BQ
eZnplCJm5qDBc2xstLAxS3n+wqJoqheqH0gAyCN2GcfraeBF6kcoEQjWJ9NwiEMs
ibR2rBnOqXyfldug3qJfbpcOq0t0mbPj2rw6HHwfusUdbzz07mkktNevssRJjgrB
/YHtGo4alQFYd3lyBldzubktJDIEdtAnuNrRXjf2JTE6pdvzE+7zmhB4Z66+uzMt
jnN6HhRFJGnI5wtCnEyLAEZVuXMjWABG8LJVzoGkabY1/qMTfeF8zjO5rfx3WhEf
akbStpxOMLrfni7dezVg4yYZhY5s71by0jt1hVQbwa1t4tSDRsp2nJkQ/2XV2jv0
n5DmFckewhFeTgLqspYtGQAA5INkJMv3N3Bx1O7FWOBLzjKqDvi3+umcynekNUrn
FH8H4xfVB1iX4LNi1CoxS7WuBmMkhFBZwJwlG71Hgq4FkFoC3AWxZ5kbA0ZUoFrq
0+Doy5/G0Id8idol700rE9fv3Bt4WGDMZT3FCMgTF5Jm2UMVvNgY/ML7nudlX5Sd
Mm9YW/DBrmvlTgar0NKT43QvS1lIcZPhxiyyqSDbHJugIy8/SFkHM+FbfxEVBFLV
mOPdZGkvnuhWSOweikboiR2m1t7VN4ib8Zga+tWQoelHnVC9rN1MDaFMC65Bj21h
/G1OqsVlAbDlp2TzH0qlPRkCPi6zbZpDbCu0azEgCAdH5K4YjPpjAYXK635DqfqI
2GRhyYRj+izzQ5abL9jCW2ljTpls4eUfmXNg7UJQ85t3Nuxp8FQxKvP4EuZPS8yC
kP3m1klgSRHDUPifClfnWXbQAUuARXY27GVoA3IpXTRS6G0B4F3N0dLrhA13dytr
c34McNc9PNtTXjhd3QKWoLamLr03R9zmNhGrIw1ShSQXgcrv9sa4RxvbQKbNacJ1
MKkHJvQoi+2M1aSTWkJKr8yoeZfc+A8sMWgXhDGNru3cI2KAkr3LdHvzin2XdeZZ
sfGhn17tdC2FvfpLOy3iS37f7CbA7/cE1xPmc2DpSpDt4YKIX78TXvlCbx3F16Xh
G+hNmYRQ6MwXsBGEmPlVLz2haaEGqtUYXFfe3DKWLc97qfR9oBGcEF93hu4WGl08
1AHlctdIiJ8ixIbHvfIgm3ojWBvQoff53iH25RnnpXeh5KRpASQiot7yjQMed0wL
QFIR9t+NrTIqYeYxEgbwvibEvL+pHcOla2sYFIp3OxF1M/Jdn2HJWJYAr76tiSeb
HtoUA1JGD5dYyZ9xg/c7khjQGO4VPRY54TqYmZ/fw/F0hZPw49wYOezvU3U/BWSf
2hg9ajGGwEuzhbE6LW8x6Yf9krGU6k5bA8L9JoGxTt5mE7uoIiPCtRmCt2sU1C0b
CZf0/vLQP5KgrBh9ybkA73Dvip121YnnZaT5+KNYfwyrNKMMW7JRo2XKj/lBd3or
TU4JTzQyzeO8sZspptZTWnkyPK6+M4+B0WJsn5sdbuXSAqZIfSlvGdhrkohrSjb4
tYENiPStyTt3ngMwIwzeeG/nIZ/oqxRpmpXr7p6T2+cVPi5Jb6LtsoILs4OA5ije
LGAJhh5+pemt4FqmDJUXtfIfGXgd6aSI24hVG+tcHqslE/T/9aCCoZ2MmxzRvFEJ
fnWdnUjjqpR7saRUK4uKcHsQ8W7BLJn3BIg6T3IY73ttj/Mo5dww2ddZtIsoRTV3
AnNjmDy9o5qHfiI1/r3u3d6Stjnw6iNfS1Pi+mOeAVJ0Xv2nKsOXpPffOQK1zSNj
q7tRb8qPfOciNqMCvO5JS5Oj85LVTZLld+8h6zakxK1dxGrAPwV5JB633mP0GTkg
C5uiQRBekuQfD2yc9jI9X0ks1CZn90ry0zWWvRjzXMHILkHVmQckk6qmiR8UIyF+
vNCxGV8rmgO2YA+Oxof8VuMfCGfASXYV6kBhP5ChGJgAI0x+e+JoD62+yn8CFQIS
hXHiwSDsOWDfyHJlZOEpkIgN+JK/MkzXF0K+npvdNzGlt5nkMsZs9Ejk/Etjbsyh
1oG2cTYobqruRCTB6ZqyF4UBkUJbSxxMl4nliGpbzyaz34A14fYum9M8zuYXemmR
djWBOYnGtqpKQPx1QaqSq0H/MTgzEGMTtysr5N/SQT1zus4fOFsoFfW7PEJa0FdC
NUaT0a7s5z8S1/RYQHPa12IwLAZh6YMtu7TOend6SAzhxhrbIsIyyO8EC4kogJt6
ThnLUgxgjOpsI41mCazrNKcftCyRtojWtPhoBVcGwHYAVnl+9MvWhrYXwxGj3WA2
TsBqVUbwKI8RX4GXbM42RFO7m1OIDsUi1V3vyPKtmmRyvKMePgTH39juG54QLKwi
byqRAcGa7PloySr61FYuO/vWNzNf5HcE4bolpYm4Hu58SeXC0HDWPBk1+8X0/Kc8
VmRKvBwBGT6K9n8J9Iju8udrnEF5DdtmP3q4FBssmMEkYZ3lDI/2l+BfbejASUwJ
TMWO1P5qa4hL5UrHsXWdnRWP5HocL7/1HfeG8WL5L4D3I4Yw/G4TLZesCCx9uKz/
RYb7q9Xq21C35Bl2INAVWbXJHEm/TYup5gQ3cddpk0XNVnIRi2y/32+Z/HAW4sFA
hszJDMQA4DGYBXYnz80hLQdqmkfRmSdxVlJJuw/BkbcDhU+lSB8C9idJ8kE8CUgp
SZXndg9id/1wiUjF5TvsURO2XACVX6xrGvCR1RMqAr+57SOcpfUBOf4WbvX2xGTt
Y7/IfxnRzh2xza2frLP1wYScanEbAvGjrO10f8XYKDX2hQUcSeM05Ao8mDVWhnCw
sKFA68TAZsR/vn/Fb47LDL6E+C1dMnIxzEH0s8A54Tc8PLaJ0bQ2rbaZncm+g3S5
YxOOanu5McwciEGESJx/DZFx0M2Otb0gAQU5+3fPrzV/JlEQJXS4EGDsLLG7GJUX
dUh423BptQmEt7xGg6Spq2ES1/YrgQGLhl+ImPOdMMpM7KoxUe9aQu2PYGdZ+q/K
+bZYwP6eq6ANdHBMJUAPntiBXcu4Al97BnimsA7IM7ULxrYZqsoWCNxkrBWzV2t/
NVIvK+2QEFj9uXYciCkhc2Zuslbo3Y0EBBev3ISGk1cyd2MTVh+8oBlDbV+UEvto
trzsFe9MVK2ilhd7Wqwiw85lFbJ1xppiJx7Wytwja5NASKnyXdLjpsb76euX3AG9
yga430tfDQE7mBVD20K+xkYsGjGqlQsrVvrww7T/Ln8TQ4ma3uQfSq7o4b5GASRy
jgaRySbWUw9j17t6cGrp9ZAQLx6aNyE5qN8egUqH1W4KMo7RuMnbtGDlN3AK63nu
NMH2bdbl3bakns2ODw6cKX8b5kYva2uXcPbpqpZwakL2YWCUxsZ9KEAcMz1vTOgg
JZK5Ld2qF4Pu/SKcPkgdQZL4BOFMsUXLbfjNYqMXd2S95LaQm0liDXGVircD2tkS
XMscR8DHWCvnkXsgDyf2afD+1BsyZR5Zhp2c2QS2Gz0TdswolHhqlpHsOGaENslc
u80vTDx65zydjXh6Y1M5rQS7mj0rrbkTQtnYDHNeOfPVqLxZ9h9DS2E67k4bfi6W
LXE3qVu6vpODi0ORd5AtihV4T3Iawg+XHBDuUS4+MQS35j1e17xY9fIABsR4R0Z3
IlMZx8yqLEGg0bIVH4BRe0H8oQgc/f/yM2xl88PFNZ3gPH07upMglTfDYnQtRLBw
bnWIYTyqmfCSImHOAMRZmT13Qm6BiXYRaoqUCzOmB0eEKDcVdgT0VQ3MG76qW/02
Gwf1R7YqLP6YTeK12DDtHvRbl+Sdzj2Q+ZzP1tIkZQ3Hj9rSjl58cG1mOe5CYoyU
jNZqEqp0knUyXQ8/1EXvTQa8hrytZFIT5t5tRK8VFfIJiUKz5kzkGogELSQ3dVUT
Ype0Zcy5DpTkOsLahtmiqJupZdeeQBR0CUT8rNvkBcZdp57nZAnBhNS7AhdUiEYt
SYdpGBhq+HZIbQDn9StyVTITLKQSWwo2sNdNuBdweEagZMUIqqth/xENsHfEhqvV
jWw84irkQahGFrhAY44h0O+oLwk7Dbav9F+QkM5ul5J5fQ2DRMa8Z8MxF6ap1xw6
NRwJMPbY6CbUDBPjP/yY0SCvXzHaGxBTxOi6wy2xWilQyL8g/Aic8VSiZfEZAY94
4zFHFnNZ0pgm9yDcgvFFNJ6LnelEOV7OXKcH4N/afrHbvEGdIZ0r/lwkNhQadWXM
rfEuhBMejEziCtmJkvOoRrB9+BzFLZbMOk9FL1kq4MV+ghnUTALbR+PO3pPihSg7
UysKFNzYsG+cHEee+glQTvisZTM/hYfRgd+waLWxj7liPKvPClOXjFH0Xi12i6u+
BUpO+wIf2K0zcXi7aWcILvrYXN/6QzuXIIQZOPWWxNJDS4Ejk1QQ2N4/+VXOfVP5
QIhKZyt5ShSmGYAA0rfbN0vKWvz50jIP3X9ry6b8qw4r7bItDQBlNGEsPiPBkdHK
DFFbBnW/aFuVZxD+Qlbh8TdIecNJhuR6YeDUgeTq5L06+bhQ7gvRl7o7TX+ylioD
LfMv4cEfNH9LxOmJ34qCYF+Iq4rU1otn0OeNwk3VEy7GG+Y63pXQbrAxjkjjhI5y
3SLENfDqc0F0XomRIP7XUhbzAOMf7+QuBArSuFqhj0L820mq/WUk+o+3uyLXiYQg
WbkR8dhhYrczj4w90LChenwMVNtf2+fR4Nqz+huusM9IJsnmr3Bsbs1iKSmEkBNn
SsMIplk2S9ahwVjM5E3Fp0ikZo9wlDC0yjmNAymlRo3ccWahULlhSPHuYzkqYesW
1WNHDIqYnNWkUld0mrh52tdD0d2MSTQz5j5cAm49/+MAr3beAH+kZUDEMBru4IHo
sSLgSKr95432F70PT6+v/QS83PXhJvwM/XfhQYEjfqPsrKH502PnuQxMLR+82JOl
WNKhukgaJ8HOlSJApijZAVbJbEisp7xUC4GxfF2o6XPSFl21wi5Il01baqQs0Xf4
LKJwrwBPVwrF6era5W5xe7Tbv1xkSFoqgE4HyDERxGILMVG6A35VWEPtzMHI34ta
2zbXF1p/qLrunrbKtdPCcIc5tLD99qBX4gxQfINQnvaanm180nFr1msZUMhqg8De
0zPFdQx35/MyRQvOr8NMuVxhVAaB7dPhJnWN1C9FA4/Mn9gq9OxcibOMKk1jqdtU
ODptU8YSc1UG3p4B36AjTl9C0w7ml7T71gG1ctYOcQxEiw0C6nATWkrmKxaC6S0c
6x7Up8xoVJ2Xc81scxBnOFiJuIhBmAzPCYDzw/A/EgKHdKLhqtluJWic3ZYjogY8
6uMXS8pS8JGEIqL7rWWCCHb93nAsdsSQSYYilRInb5/CyKNTrP3rnLEek0OHmhlf
cd2oVkRgo+eber2S9O6MytM3us/KQfI415W+CHfy28H6ZXPXHQdB58NmO4gGObhW
AoqEi1leTJeAJcQU6h91fCvTYWxM59vjCPct3X0VinwfMUAWHs3lk4/P6ZQ8TPry
D4MbYcBoXdnu9pZOeFwvR9sOC0P/l57ZosY6pq6bAA1weL2W/7jQL9M4XhdghE1z
RrF4h4Bj0L1r2pKUFHb4yv5F3LPrfjKBCm3IfbNnUI/M+BOWy3cq8Pr4qLLFlj/b
+HD/w/o1spWMnpOoIPHTSPkMQs5j7WAbfMJTD2dDFgEbBpUn/uMQIq+NnzhWmzgl
CYPUxE0kpzZUt3WT4LTAApo4VQlXJ/eUnvqRuVnBCya+2K8qQU/CiqpdnIJ2wdC9
aFX0g6qSl/aBOcq6DkQ/CIvYg56i2u/MQPuNGpVnRzB/IXjGMiWCeuE418nafsKZ
Q515jlFKFRpnzA9poeMtMxe1HJYDFaMCYkjh+IKntoNY5X1V9Ebcirk2hn/em29a
ccuuYcxHE2sfoV5OODH0SGNJ+fZLY5nxQBdNNOGJfo2fdp3UoiNr44gqocdpquOr
G4gQvFvQngNNhoAfZ82u1e4ZGQnco00hXPXcYm4CgwEknkqAy2NzCqxX3T8uk7lN
p8akZ03UMkLUYPzmdVkUIl83BmoR2PKLL9HVCZUKsOdJbvUNA7kyO64x4DWdob0i
NFIun0h9oDiSTvKlW8/3ol940U8qKeV/jaz5xD1ePBLR68OX2rN1j+bpHTSVv06u
+5xyLzsZV2r+8HdIVPkOc83K0HHS6S2D9/vIekEFBh8pAfGTBMLqhdzbnqkuXFy4
17UiU5SOZ1t8ZVWMEwsuX8QQzIgoziS0n3dsTd/tUYDQCearUtrrzqucmuQarV7l
+rRBl0Rqt+H9HTkwvdcLCe/NkhoJcCVD7qLJvmYYhYWQ9YkCN7lrQ/hLCUfDFB/5
Acu0MIaVmcFSXW9dU9y1mngkTUX6/77gtaABeyk6fKeTLd+By0Meg6rJA2l9BSf2
3KAvTvTNML1QMpYOopWpsJwqem6Lp0mDfRE9DeAcSQJJy6goohAsBiLTUHi7NuAv
zYb2FiLDwXreQEtAdICNBRy59bpDJq842Tt9s/5OFGgUMIfkIjueimkOXKNi8VTB
nsoJ4dlWH1zn50Y4gQLlbN8ohB/FVGsSkKcVFkyOq8cPR79s76thQDtXBv28bzYk
i1xHJhNZznCxct+6P2+uHd5sed21nLDgVs3YJXvD/SJcIBa4BIHaViqzjFxoEo8M
3a8DXyEljN/uqpsjAFx5hs5qI+IU7m3DZJ3+091rq9s/7616MTFXp/g/e3FBMtAh
8EhrDMFCYzNtajINO2Cc3Rji/BM5zAyVqNV2oxgQFNACO1Jyd0KTbaun6dMNTrHK
IfrUTduyJL6b0ciQi4MZFFGKSmZYPpRv/NP1cSSA6R8O68a3h9M3cags3IZxX36N
qIgRxxklDjU13WoWCSBtv610UETRmO3ed1hcvUuE5hhjx5y76ASDTB4zgQ/sleE1
xqOCFXExBvIjRH1DyMmJGSlUSUE3rt2H8ilp1+Gx6aFxoODfuIb/4O3Ws8IXNHi/
CiBfRdgby20zcObxksxQse5kd8lxqsGAyJy2Zmcg+DS5WQu8QXCxBWXmqKoOw1H/
PC8tN+jaz+8Wygsm+bbomkvTGxG4hEryalATkoZOaTlze3nfpEqUqePgCKB9I0k5
jqPP7wosdxTQ+81gJ/FaDDi7cQllXOiQ6TiCw5GR+KixDWhNjsZ0p99Bb0eYLoPg
yXILHvUWLVNaOnTdPc8DjttAV8cEXh8UrbusYJbu0G/a3cqJrYbYoq7uHnmF4zAt
+PFo0+BwldcyODSCfsYtgGyBPlU7lmN21U5QlVuFg4q5uc5Ul9j6FiZv35PPN7Vt
/HX1fS5gYj6Prw1uQ0OHNxNt14Rs2+UiCI8k7trGejOoUqsGnqvFDSZOAaqPFfFj
zidvwrCGIwNLIiPZXjnrnnVN+bVkEmzMwpCJZxNMu3LYr8X0HNMGymm0gbWSiSau
DHfxN5geFgIh8FRxoh63h5zU7hDZ8CRC7DYDylMhJB5f96zSf2oLgNSH+9WT1ji2
CVViV+Ok35FrxEwa8FVYg0TQGGgNZ1AV4gMfuLxQ491rZfX6jOtpE9u9JfDMk/gR
2jyk4ciY2sX4bDttrYTlEIl5jeZjb4VHpGuGYNwWTZXujY68mb+1J2kfr0OrYlYE
oMHsKoKcXpTNpsiszHe8+jAKTq7mXVw7BiRoImzkzPlXLTt4mZhJV45o5fZ2QK+J
RozzHmQDFtDQpM7hl4UvpFLxHo3nrRNHxwkSgtAvJzAAcnK8WNU0Ulsck4Wm4uFH
fjJ9XnzqlN5A02K5vwwFbuvzMJ/Tx/jgx77w7zTXNlyqSqSNPxzvzx7zWmuUXGnF
kH6lOjk2pjBmyVNx3oMqKqgzTnyZD5KEFc5K1FVzyDGjdfdX9zog6Tlf3ni1Xbmz
JCXCAfa1gS9QSVXubXojvLyxl7lCCWuwftuFOTICb1Ke7EQySvYSIYcR2NJ327df
iDj+fBtGcuIXrlSeBsTMmUADN3aG9Z1AqmiRW8lSw947xtFFyyOYuQwXNIWtSA/4
MO2w+Q+wMzXg3LAUcdDsxd+9/T2LjTHRWAOxhAuCiSNReh+edsP9YovCouNG4QY4
EtavVaYcwKDo/ZDakUsdBu2Rxj8NCJBJeAHOpm5d93HY0wro3MlepUTdqgJiGva7
mY54KL7kh0myHybWFu93Ek8S14Ga9LR5zLE8s9hvnfvp4lXV0vZVUkMVEVicstig
DdFOTjkw5zJGFupZlKeyfkD+cwVRo9eA1zwyEoljtR22oHkqvPQ/XuVVPws9gTV5
154kvcIIQjlSjmuediDiOQ==
`pragma protect end_protected
