// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:51 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qc7uh9B1JgebVeGIseu41aMKGJ7e7La7gF16EiwhyGt3wj6DHmjK9v/tEBhuHgsW
ULf66N8lZtfVWU9tfxOcy4AkGJM3aMAI3onktBF/ENa/O8zCHT15FlmXGcDTURz/
kvXD9k8QLj7GqKLrktjIwWSB6Ais62xZ88/SbvIwz98=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 47808)
DQHnPrWZTCqnbf6opKeu4X3lWfZON3msVjJnUEMaeHXNl/DbFmo9nzQ11U8faPrR
9ggFgQQJXO7qrO3k2zo7k13lwJ+yPEPnI+WoFSbByqIE+r9gTwcx9mZrhAWE8V2W
JJoNl2gKilgjpIkIfuul/actQtAqgUwHpRyOhOvJYqnwcnU558Ss/lqc+kCiNg4Q
nyi/fjEBR9r8Gqq/LZ0X+D7y3iKFVAWKPqFGtpOObwY3xdh3xzV/6KwuvdfG318N
E/SQ5xZOqEKqYq5o+wxbD9hqeMzbNthu6+Wuw7HBtLmFQZ/HusNCYCF8hNc2Sc+X
e+vjR7RQKs4k92J3JkhaAcPGq2XHR1lcHj8pMq77n/0htvIxpn6XkIR956kg0SmV
eAfuh7wjW3ACMIWxvt1S3sdS+mubTI3EmsgYyBlQaYEucD53z8pm9ArBpQTou3by
gGsVJNkQ6QEJDr5XOOo6B8J+X9rMFoZhwXBEbUuCJdc1Rr8OGyTRLMSsBnLZMwUK
gh+zq8ZLSqVtKT+eaLsPclvrYUJR8uNTDIuuoptlxSihZqkj7JZGMyfsuQNvv1z5
JCKzYxxoeDqdpCfKniwUskNrm1QhTdXJbD9LNgHpHp0HRl9iOL19gFELqLHfULWt
vqaaYCMlHs2BmdTp4SUFbIOsUM8n778uel4QsFST6AC+fcVbbGQboawzrf0Y71mq
3RG8qqrhZos/mUYX2q2tKDMeSR3yw0JWggG14q8lSghD7M6UQJyuvgX8/iYftsMZ
fz3AtmpgYCV6fc56e1XkWb88E+sbC3cjegscY/7s5sIW1KL9ualwTGGnhQc/8XS/
6R52bQa0EQj+Px2fu3q/64eiOFUNsHBPhtYhGfIECc0LsOF2v1U9hZWnqEB+AT/h
0JVzPvv4C2M1YiL+GAYpF2qt5TUb1X/nG0JqiEa1IULyXT2/xheJt/+v9/rHtcHj
EZZmrnVIwCgbmdmtHlnB5K07Z4I+ObeTpGvn854I2V0icgZ3b+UsitzBF/DSGSEf
S7r2SaU14dL5k57H5+Ei/EaJ+/8dxwDYb1VG9u7Io471U3VWhQ+ABr1LPCmNv+wM
ljZrrKSK1XTrTyDE49NaARLI/ZVznkCR21mzHTBF/jJ9mREBM89h4qanaj6V5MsS
pwmZjhwxx4nCWtGW7Mtz15fv7T3A9QSwfeAgB7m3qRwNzN3xi/7b+wnX/MGe8zvk
HBvw8HwWNfSSinojOrqzG9gtwc92QxZY8uY2jcBl7d6xEqrfGqnYHo7zuKNSmYgp
iBxx2TUYf+eGOce6ZNY8kW3WJwiTv5vW1wl2E6cLICH2fem7X0i6WTIUC1uyJWKd
6HaWVX3QgEpSoCFPDSpSF3fopTix2MPWOt5wuzclligiuRuGrjKuoh6V6JG+d7UK
NsL6zKb0OyI7oyuqLcWG5VUx3I+X5fiOwRGGfVK2UcHlmX+9XWXgJHbzEEEMblFb
71UcCa4pJ47gTYZInc7+yzKIsQlQwLBhV5o4KQNbFe1GZtABD1Fgg6DxPfddNj+G
HH6mjqdOyVPXDRx5f/q1aKHdAjJ46nSXYVQHyH5Xs/B+YrdpKWiX77czcifjyTZA
a5deBn6RArocKkwSKTZq0S2bXXjlulKCREUtHHuhCDPJu6FOZ32eoPjkLzZ0tkYF
wxUduvA6EiWxnWMKOGS9aNihO7lNjtSNjJlh0m/g1kKpqWPGJhTWQQdGYi8sf9aB
yfyUChSjnQKXjb1KZITpMLVCao7nbCOvokUjaiAbqS41dCuV4ohfZ/k/nOrA3pmv
1jFcT/OQrm5ilMvpT2keCyo2Co6E1O0NeJ2m3b+KSUEcd5+umTz+ZoyUe9Crk5E0
zuROXY/R9aRD74G3yDnNS6lD/e2s9X0PUB/ROTMUiDzkirGa0HOBg0sa0mCBiXrX
gZqUi2NcGWwC+BDktN18IN8J4pBuWovq1dwUMCNVPYjFmIJJxdpWuz/ST6WC6zoY
/RuihwZlrWBVj7Asx1qGC5dLO2JZeTi9EHFenRvWFOebzq98OIrCnoQC5BEzKVOV
HMw9A1qpDdUgmfp309/iy/Sx0VuMHu+7Sg055liawTM++fwqXO2Kiq0oHrr/VwAu
u/7k0UhblqsKrAKc4o4kBhtp4wROyu64EtvQlipRjMStUhsOLUBVkqmQgR1AOuaV
H8qRZ20ucjdgS0wFXOwx3kgM2sY2gqOnfW8B5CBVRM+mSfY+1OLCl0B0kA6iZYYD
RgaZb1fSofGRaXLbVRRrWcewis3cs6ycL+5JQ+m7JtEmCvD7Slaj8ArbvwL02yb6
3+8CN2q42yXHj9w2tTukP3PQxeI1cgP0X19mQvYJJMHkuNpVXfbhgxCftt+H1dQl
NSYi0YvQx9qaUoE40sIxNmoa3UzmeAmK8QHuRcQuMEB806ZSEt8YWMxG322i18Zs
6S5WligdgNjWdVQ/gtuedYbaDo2PVpuWW00G5V0LYS3oE1Idf5KR0xImPcXsgzat
xlOL1+QeG14Ns4ZJ5bhvCo58333QPD9KAzC6V3EDCtraqiphrl6wrp8Yko/qfQQK
YzEz0nFsQdYAc2RnvQ0RRbWgz2sziv59b1JFNlY5Yn0hGa33KzrbA9VfY1HxQIxE
I2Luygc+ltw+vV696ocdPiWu0IwlVcEaSxlHHSTVTyBdqQWuV6F3eZH6sjaGFY9a
paU8a81InfnWoSuP20zaDwUHiwUEHga63qDBfAWr6X+BC+nq2Q2TU+uLcOYpy/QK
Xd/1qG2dwRf7tJWWPYS2HLyJcOuTXd1BUbMU1G1V22TI9yINny/7g0JTMe81XjoX
puDXPokvRQ57rnQRjKRE2cO2v/BTIGx8ulVedndIy9pEPvkUJPJREkTJQt5vxIbA
BMWhXSZ70m9ZwmOLWD5ojTyO/NwQhutvryQZ0G7WCC8UDWjJwVSQIGBaiL/ttSTH
68KRuEuBO6TPzET1dNVBOjEH7NX7ctTfdDmwZf/lAI2+GLOnSp053Z7bwS+sA6z9
HyXIWVQjwj2MHjWDG3wh0wiPepSefmv39Nrs+YGklVB8a36r1HHqwKeiQFkAK2C6
sCiDXhHi4XevZ6O2Sj8bhc81TQ+Y+Lp52PmIb6UAJAZsRbx51hthdO7e/yVRSlCl
TfOdWuFZysgbeN/mFUD6fvQhbUWDsR0+5XmuHTp3JCRbALvhmmjltD9vZevnhvCD
ehnT8YZQRF9BH2xJIuo8eAT1Xv6h5fOsmjNaQqyDRiQcMZhg7JigT8CBp7QDbhP+
d0pV9J0SUkIbDlQsoMNNJONsK6QFA9n5Vin3yvS2g36NC2vciQuLO3B+XA2omwni
2jxN9GEb4s+2cJvWFcUCXmJQPx4HozZrKHudQOoK39IDGjuiZPFgsSfB9N3qhF86
k8qSHV2gUYiwMVqGpxcUaX9TkmU/hJvg6e5EOOOvOzNsxSiIvQNxXsPlNJcn8Hfu
48Df5vgdGHRaRY1DiM8/jSbeVuY6LHH+z0SQsXIbiP/izE5rZ9Qxpz9iOm+ZVIKk
84oUUOnf6UUYYa7eQsdMaKFbqmTRQPXcd0I78UArKA/fHBBcnxjriYG5EjBqx2F8
CcNtlsOqjJPLnHUe3IylDfhNNpHjCc9yy2K8Ij7jXUHTEOVUeRajrEjbS0T/uU6A
557sYs2hOVF3GwC2R1PYKXF2M70w2VzunzqM+Quz3PnPyMLl/UTce97wbMg0Q0OM
5VQODwS4WXIWpYXV+REqid8GTSDlvDrUPAuMpA9ruidnsOc0noFgk5/s1mPy3lWT
LYM9Y/OmFzTkwsH3+k6BllcCUzy+du35qJalzGDAUACuCJkAxG4HFuMOqSpmSTvR
3IfzE6r5Q2zDWbhm0hG0qZRhMc4FswibM9uIEHi3kLS0dFsjja5JFVCQgBkmAOfL
yS6l1pigZRfVOzYS/2ewQLQXEF3IqgUhj3f55m7cKER/KjE7HN1Uu9oA6iIZb2rs
jKQ6FENMLz3SiYV4Xg53BiEqJoyXj5JU5gKNGBKUfzRRWUC5IR7huKsv3DArWaew
FArunwSV7zT7SNhRT7P0HD0HNvPTv/ykrefuFDMrdPTm7eo36Gr6firk4XHXv3lT
uNp79arDYtv/F3xmnpgmnrz7uZwkZKEDtOkETsmo7HJ3JyY42WZGu74rHLamjY/j
jwtF7cdP+5kg47HVk+0IMNj0aQev5qQWetxqLUqa3zkMr6b9bdmWrqxfT6dU4nPM
D2DCCjGuxBp0yrsuIAbMNK3gG8ykIbV6j+15z7JmEQWS9ROOh01QS39+LZaf4yuX
dajU9ilzsDxE/yu5nFwgB8CdHXeDxGtJzMl3NKmWHmPQ9Dl9LoB0lg+JbqVk0Emw
5cPC+SHq4p+Beu+W2zkpVmYE7B0+GTgOi0rt0Nv6OF546ZsaLjvc3FdLKLkQVhln
0VwnYCL56NnuCzldyF9/eQQs57yxNJbkvgObTUqDZpt5TMJvX9sdU3tdM+tq+sNm
JJJ/MF3GHsQeOWDesFUX7SSnVu2dU86B/Hcz9/skdC7n8IIrJgrj6+/eID6uzntG
F2N6JxAdtbh2PGMZZ5VSp1plkIodg7wsBDw9Q32QzsPEJzOY1WK1K/53+yDQielV
8P0jIGxCmnJ3NoW42Fh2JKsrtdBI0fQH8jAxWPP6YtLGorMOUTvt9MoK3oSGqks/
n8Pnn6wT2/9ED92ifSkULvi+cAK+1/N6tb7SOtgUt/ZcTI1Azk6qh54SbY1c/Mqb
gLreJ3TU+ayKKd1Pq3Q5jklrcBPkHiWErl0E9w+a8WGIEyp1QG0vabXPnxB96BHN
1pmf/Q0WUtVodxWqVhws8Z0kn3fMZNaU7CHRTutuQZYWg2lGwr5haW2y6Z74Mho3
UZkXrhbAgahp4UOP5OpOInFh6QDzY98EjwJvlBoL5NGYtNSnpT/yxouv8Wgd+wvd
v4dVsqbQDW3JbynYPZVsOBMFvJop7boflWh/3WOeYFFfRErwEEAp8DP173LNC83M
qwbMoRmZUCsubekjHWeh4+zmO8A5pH2kzIDphP3y4R5gODjUePs/pPm+0GmVz8Tu
rrZVeBX8HBwQ5izmZ7nFAcat3nqLoiNBTA0eHoGu+uOUyQUoJhtOhMOkNeIypSOF
ywV8DakXyXxIKlqjzGr6KjiOEbUtrh4H9gsgraRTq5t2wzvLLvwrqpQtCD0FhG8l
+faTnnYQIIcbikA8IphX82B2oyhDW4kD/0hECHgXZ2QfFIBpAybmSaf8EvrDKU8I
59Jy0rbTGZutpevLAKry7UboHnOq3HM3u3vrkYIZ/Lbj06FTjtuG27325nuJO3Dz
7hjYdfT4qbj+DA7J8RLxkHYlZUU7tuHQaEY234tHEoBtPOeaxDqWc+lNAnydxVvF
MT2JrlBbRH7MwNGQfaZWImeRPD7iq33EfrshSXgoXvzERJnukGnxkXdig0mlX7OO
Lkg6gKk35VafKcIObiIqzSeCP9j8/OdiKDyn1peuPg5tmkfrpG4Rz5Q1TfxFf5BA
3A2o+2klu+Ps7BD6uE/H6jSITVnxCzo00Si/8cLXuqkM3nTfceI/wRnQXzH+/2g0
kJYIFqMFCR+wEJN0vKqwTQv8pBdxuJouBMi5+w7hZsLWKKBU3iI7dEwpssrAYF5s
oVqBpZ4/V0lwaUpF5AA/wj4ADeHUAIToG5gaR+agw/eqZ2L2jWbI5vnvg5Wmm61O
h6ReVAx3F2D+1oEc/FQf7RE2Lvxe8b+7Zh1Zeu4u/J094rCWUcii0zZcmDAfiPbu
84GVx4pv3Bn+7Zbqwgt8dQWkfsT6hjg/4fSyNd3dEiwXhF3AHL1+VYp64FhVW1dt
oGDmghhpQQooPXx0qjfXPa+mZ4TYz58yYp8AdmqZtwYwdk7HU2A1pK6q2Zc7UYvP
4/aeWxjU0Obz3BaSlXVVQcJ5NRqB5VfJVOoc406F0JitUmBGxosjCUh/n4GhA7QW
//ACpWVkFXrKrDr06YwNi438uu3P1nQ1jCD8cofLfpGdHmpeSH71SAUXkomy0s4p
Q7V1+SGlQ+LAXQORCEwbDPqnsgMgHTZ49Tno3tNhkDTD0/VAUNGwd8GWlEy/zwm1
E33+niwj390wyw1lz5K4Oqxb8Ai0vohwew11QlvA9VaYVz5hXWokT/Lfay+NrNur
7h0V9uGaiz8b/02UdDCK7U8FtTs08jqpNVu941LAlfqGVZyGnI3S4Zs0wogYagZh
VloeejWaLibYaMe0mJiD+fOwZGnvJFHDtYcKi42S5XBJEZcLNNJ5R4YsuvmJkisY
i6pNoo/Er6B2p4ieSuLp2nmuAaCBmcAwogZO6KOK7sDkSs+rqMOHGvprLhRtmb0r
DiTiYWUIskwpDjqXBeG17BfeaSY/X921+T+pF4UYZr8ToQ3De5dsiBAK+tB9URjO
tj80z1rwXTJO9upL9WhpF3LXmg91HHELY3wj19qKkSBwMC4DWZbVmT4smracf9wz
yh5xzDZ05vgbBh87qwD9L8z50t+mDpSdNhXA3VSG/ancyNBXtV1Uy4K+/+T1hoL4
2m+alRKT1LADzLXnoQRrJWcq6ae6Fjm/Eh0DjEaWXp66VxnjxFSPjPfDTflYU6k6
RKgG9azqY9HgnFjiLhnnmaL3FgkCx5tPNaM2SVZEICdAkh2wA+EnpErtyoO+oD+C
wzZ6hNreTT+OSgs325s9WQ0kmt8KmKCz+xY+0R8hyxZ4BSb6jY+0x7L7UqHQ0+oJ
dRxX2Gqv0Lbc1BqktB1icGnZMIAQUmiV82jpVv3KQi4iK/PXU45OX3syhrxyoYnS
+jWocAgbGV36SQoxhC80IwI9VmalkpjHwP7H2OBTOwH5GhHXweb0YceFYED6hXVa
oqbuG4Jl4fXeyWI1JGnAfshIy0f+8StWKm4HbLbOaUruNLbUjyJtnT7SJjLMahx4
B4KfZHa31MgH5r/PauS7oTEMHT+Nx7lpusohGEjEhEUA4RW9sCeLQ/P6lXuAvMx0
0Yly82gldg8rAqpVZwlO6IihROY2Ij95HIdKwC909RZt+R6MnsVRC56BtskczDNa
UcagshNF5uUOzz49IPhzHPd2vXqODz9H3k0nZZxCB8BlQeAtpLdyLuxpoDeDFMQe
5TXLv5ub7gkBgnAbLDh4QTKRTIaWC7+PKAFV2JVowYSXCakltdHMAkffu09n1xM/
7qdNSN3jKBqbZKUzSOTW0QFVUb54AEZq3ztjtWpPGJuZ0Q/0lSa1YTspYQd6tzYN
0NyP/fmvc64MhzzBgLx5bT4wTEPCRciL2PChsT90OQzblOZrsiZkUNEHLQVLpggj
gBsAvBU8MrXJCzCIg/Qyv1MJOPFjtqV6C8KPSmQe+ThSdQbMXh9ZEAJ+Z8/Z5VF5
BlmBfn8WLdITbX07x8655afV2poO3LDzYTnjnHq163HEWDGXBH4UM2SGsC0kBPjO
j21K/EroBncUhcIECkWtiOp05vLej2FYT6hxwYGj4x3KACSL7qQTshq18uPLlnG5
0gk6Vp1/YBtglup1YDNPkZjMs6qTi3itxfH0F+YxRffFo4/AWUVCC8f5CojBghbn
MHXt3V18L5jroinR2nzCtxUGhJ0jJByK7+70Vk0sLZU7hsxkc83v0hY/hUiMGBDk
VDurFML+t8ftK53hjLUKCtcvTyvPGfzaw/wdkcBA6plUDN82mxTM84ECdz5/KPlT
OrtoGCeWOoEzTuQ3NKo9R7fq7pQK0R3w1K2oVGr5HLqIhZLrQUyfaGtGyxeDvmJv
KTd79ydtwt6YMhFeHgqfon41c7eu0qMDrWtqMBa7elJdpZzFKrD1csOPOsXfTMeE
werSUNoyR3+QtGAOnM5YGGIwE6GKH3oF4/9f7u4BNnoH29vizS92WbojiqDkUSYp
lHJgEZIS2G+eSs0CKI6iNjTZ60qCgTssrQ1qBCnjOK8T5JpufriBzV0f7+rwnEeO
Nx2sHeUw7vHloEF09TqMjGL0S0u8EW0kBEpwWmW8FSzS+6FpKoJ6LMhMHi8C3Lyz
537R6c99H0ystL6X09RG13dEwiHVhAp3idTbTeFvluPcc/pJtqgT+t/vLsrR3xLj
ybV8V2t+1WQWlxZViARIHpjk3W0RcfHXhQe0Q2jMVFTO+Wg/4CHvE3wNvL6su/D1
RXZZbfCb79odRKrAMbt26NoRqT8tdNhLIz+ARiVJZdRoe9pYwoLPTbNQ8PpX9Ufn
KavrSCyISWfu7xe5cPKUZqv1gSnL8VWEzkS3edvTqMCG92GtgQFf1Fs788ezORlf
+/BEt2GoOBToCLBulqoj+cakPuiRUH2phbtFP9GuxOr4PkuovhTBug61q51UuXrX
FAUifsTXwrfKEDDe7XrY2zV8MDVZGh6Q1LXj3BA9Hc3z6uzwc3qwrlTpSPcfZI0E
lv7IasEtxRC5EC2aJZPm5GGqRLlQo/gVJKOq9IwEYMt4FWJykbthxDHww5SBvx4l
Cko7VTb323iwfC3IbLvTq1AuiuRoMreSy7yCvbP8sep1kUIEzOoNMywqzUgKj3yX
rik+B7C23rSTwbkRAU6ggjFkDtWkwCv44rORuF8dkBrec+/vdW5eMXAQk+NHfjjT
dMTDX8ELnlj+MBcwHoiogNDByzlFAIHd4uwPNi0Q7SizjzaLDPWB7EEFf+4WxWHO
WRGzQf9cSZIRmecrOhbWogcBPPZBewsK10sxaM8yw78yg8sltq7hjlizXyooTlKG
IMd7H24E6X5iQADKUBLA0kfGKpSHwqmmVwhjQQCa0p+10M1DbSYVBNtVTrteHoNa
xKY8YqcJaxudl4deviXKneC9+8FRn8lXcLP4EnEmO56qYBE50pNt98t6uiJC3j8z
zJGFg8CESV/zWvARapPM6FA3mnBun4M989+TnsISEm+qNhEIII4HSk30i+y1e8lD
l5lq96jlmVC8OjhIPNnp+8LBLNIgu2B+rpqyfBpXpUjwqjchm262OHKOoCMUoJTq
DT3zx5fzffJ4txwgcGc58QgOxBkd11sRIpUQdYKX7RIAvXhvmL3T+Pkwt0btfOGS
X4r2H0zNgqhJwaqJdfzCfkfnoNxkSh550j6zn3pX4CrQXE1erfDZZjE3JO06RyVQ
J6mCJ3IkPtS89znEX876m+9NzTrUwxPU8whSoKkzX2ulW8e7/JfWGDJ2sj/pj/6e
gnxGWvGa3TcLurgN1LuG7kh+fObOm1I4VhWO/P2+WXOKRVu38QOlW54OkpSnoALX
ZCypHscBSt0omWW0VwTMFJtLfeQidJjF/3UhkLFqFthYb2Q/q1o7wK7k9a+IzPxZ
1jd7VXrwmusvH2q/oZLhHVSwxCT00IEEoxSDy+W5aC6tJpep5x4poSIi5auNRGpu
/idTtp/3g/LZyLiFuTLtn3ewWyhV7nGmt4s8DZSERlsNKgluY5y/86UjVCfEVDAn
59KihgqTKS7Y8gIirDhbMUZHZGD7IDBJbmp1zwbO7FebZ+SV2uQig8K5YaeyVS0I
1jTG6zA6ad7hIxZldZinrc9ZPrlKNirl2w1QNOBo5g08hdCPDLc7fEwlrYK+eMES
qFc//5yWSLjVeeoaXp7YEtPCh4pgZREn6a5N6ZcnSRr++Ojc1dH68JIiAeL85+j8
wuu7RcldorRs0k+ydOAPWAfK+rNDvYsfWo/xzcRYazTsCTccVaLNrwsJ73/KjIjM
mgU+EzKMNLblgKGajJIDW4Ar7iEiGCMU7WU5yTZs0hKrVc85JqVwYQYCsuU1dcB0
lH04Rbs2W7PMS9ASdxYO3l8xI0hfYJl3QkvbMsvVyrTdEXoTScR0XbmJezJTDdqm
nqK95MTmWYaEDbVppecBJuWNNVVLOybb0xBHJeJYH+ZsmOraonG4uzViojmWTbXB
eBB4d9CWmrr1LrUeNi7mg/UUjBNgdhoDjKqWsVIfQXcFAJH2DGQucK3RbEoOo2HK
Yklgsy9pKtCoDY0STmDKfJSrPBmz4O/jRqjwfypyMeTXSeh9FCpGMT4zVGTF/lwU
JkxMjYFsYhkVAxJdGhC3vOH1RmFXUjgZ0U9dKqE6HDN1EI7NWTuF/YxDosI3Hpaf
Aa31dcAFWL2lCwu2Af01lzpYTfFEq0MO25w8vHxLWA7blPsepUvDf2h7ty5rVdhc
MUdJKYKSBaPaz6nNajVete1bEGrqEyTV0kYeqKwc4VNw5NyZkoOApkmh9Pp9Xvo7
c51J4VsGMq2zhr3b6gB6mdKfussKKPDJVONu01EIwlSR8iux8eS2SXB8BUUW1FYg
i7sSYOwkVFj7+C5Pebh/bYRbXDK+//1hLDQCxSHA+iDOprOflZ2pvx/zfpaD4EdW
XxSuKGUj/Mqzh8PR8oOshtWLFdy7lz6e+5n3RWuVY1kboy87Dz1V3ibwT9YT9SDc
NnJTYqUdKY1x0nEEQLbWoC7fVWL6B8oAsCGRn69+KEU4MeGEXfF/RPVKFgPozwik
+D+xA/wfZDmpYkBBPwFZquphWTNSm4K6P97o2yT/rCZWr2SLJ9UOlRThYpkWsZRQ
4CVYJKRp9npQ6QOnr80mLn+t5njdCPTLdgXLDgbXX/tPz4qHJnWRjuM3wewkzS4L
WVJm4v3t4LsEgU3FprQeSgf32VMKcu0DE93o2T+naPmfEgL8Yvl+P44njMfU2Tdb
eB5MvyQcucZebkaqGULfUjbqutVkSk6nMKIj0p/KX+qvM2T7xF2Gb91qstkKO/l9
rCc+mlMYqh+/8AeVpcdjY55x7eePJZiky6+0TI8P8xzjrgKA6gu5D0zIjmwe3HS3
vG5rma+kc7GeDvWmO9FtYtEGoaQcN8GYoJtCqcO+dfcfwbmnS4yUvQOZRLmlZO6A
vlAw++0YkAc5lX373gwIFSbUOV1tzpCCXvxmcoq+jK9fV5fAtc4FQP0Q/5j6Vdjn
dF0iOXl0xZ786tlsWUZP1ZEQMHWvTBC+sTkhEkCX0x+1xzPxzwFVN5OVi5SDzkFw
uLkDsoDlCyE6m5bhBFIROfHktQu/7NsPAQyCdmEdNKoUvgl/NOh0IN7bvKHAWCCl
IF7LD/BuBwcH6aot+e+GVLSrIyHcuXhr0OXqH3LnryrLWICLWHaFg3pL85mPwtpi
OArnY4+tYINQZs4uXWUS/xtBBjwUV2MQO22N1l48o0DqRdNK93rSEGh+VvLDopz7
mBflhelJQzdph/Gcun4UDfXd76iYv02d3hwlSJQydtSQvF+oIOalZEZgxeJ45WXs
TilgC663EX7ueZZAKxb450QDoxwEmwFPAfqbIlCUMso/+uzUHn+meLyL7q6PjGnk
KacnHYD0vfmiJj2TOKvgBynAYaxgwmy1C85HwMlgmxptGt5KUCVZsIBjB5yp5yse
AodT+mQcN95RhG0GVxuIreaT19F7/71RLXLFcuXcck6jW/QFZ3Xw2i/MwboJ1wpw
Do7RFuXzoFnAYDppbdcCKcga6EpRl8KYpxysgrwb4KfgKYKbddwS0jt0m4IE+XaO
NpBSMl0slr2DQN4X2PIyYBrQJjc0ieHm4oECz0ByPhQ2fl9QYZNEAnERxjsYz42L
hQRyJ7rHI5pLDVOx0y2IaEOQdXDg5f639EuPl5monu/wpYqmHfNT9UuHfluCTtKU
5dwgTdoASYMQrLWN9vM3qzPfjv1tWOpa3fx78odacUuB+gutSZKnNyOk3Pj2/NQQ
Y83Y5ZQV6yNI8e98yEhLTUbLJO/0K8WDVXoo77+egNoezh2sHDUX823arBrnFspl
lRPEFYRYNbARCNKu7W9RT44VJbs52OPsgivhXOgByDj/wGEYd75LoBTr0NLDpV+U
9Xac8yBQe4M9h/LvM5H5Q3wcPWeIOaDMdxDRqD3zD5pVXmO9ZBPbL+dnUqa3lMCU
nWDuPeQeVa4/N5XS+4xzbr7o3pVYRYMHhFSjkWKb9/exK2GUVFCHxniX63/h+jiT
DyujNjgiJ+MKK5Qx7+Q/e8i7zxuQkk4Wd4lWj2+jXNjY7Gz3jvqZoqPC9/62YXXP
/bd+hT89MEY03SrRQMF79S0PMuxS3xYjeeC4VbDXP7P0+Xx/0NZmaICcGH8GmcHR
H0Oz1xOLY+sEZ8cadxOfUVIqVGAXXsm7T7oNwRDz4GdpfYdoHgwV8XCNwvGLe7Ry
4/uC3/x85sHF0DxajX3QwS/0YbRXiBHiexaPLsOgSC0EI4B186W1nzTrCGnwhbPB
6aiwZpv6VOUAHsoIqKFt2Qd/GUsCWOX2wzqBkilZzI0oMMyWGIFJ6xmjySQrXa7K
Gf2Bn3bV1qnoiaG/xcE7dtq0M3SFAggQzT2fzhRpduLtetv0PiVCHKNd36BSQy1/
U+KVZu8okIUnAbXXUMOiJRPYQiXPkjp4pwQt86waD9XAOHxsdRlQ/urcFTUHxiH9
XX86p/7vcn65jE0WCpRtNqWYnulxeDhF4RTTVcQ76DbIWz3GRynF6Jhum8KOv05Y
Wlqr0tXpOWCvwO7IjNMci0Ye1V5BricJnf2fKdxQBsl37dcHG+sKuhwksGpe58+S
rOxLSG636VJGTxxGIPBbmRL/cBINn01GuaDMbpXxO/rAP6D9CP/iFdF+/hpTzn6R
daoK3a83kTRWvM9wdJ+DF+DCf7EsuXhZlypwlXO1KxhD4tO/pxS37g1+wszLcMd/
fSWCxF1w4Bcocs4OHOnu/UObq52ajgEz5d18Syvbq4LEsRcsxR006O9YGtCNh8AX
NGTpRLzQer2w+UGGuF8ANpOVcYAEdRTW6kkUQFtnXWVI0mmrG6hR6QT8bd5GQXee
R931C0d7WHFwCg7Ht1+33oA8wlzS2kh6b6sUd/2lEVojANfV/x69kIqfLe/x6S2Z
VDTs4hk+MOrDGMs+bA8RaCCU+X78XDzm3UDdxC+1Luvv6rUnJJuPLM5y5bOvw6QZ
jm/iOYUlRKQv7igqdtMs23LJ5r8DIqMTzuuyr9FXsCM9+KNakRXWt3Etyy2zPLLc
oL6CzEaGdnpV+RcMNtq9Jnz7mBbEpeWJWyCAsUMkgjnmjrhVtIF3uUlVOVa+drkD
kZDAuOpXBWugwMUQRIB9h0bBaHrRn7aJmkN/wJlZ8AhSd8+TE6KWsss+LcrfmbV7
M031yQuVCT+V+/4HtXcVZjvJCqsqwtWbGBA/rnY0yyZNrxUn7MVtrZ6qIy3wV520
dVwZzlzrAGaLPkhcZlBEY+hhJXph4bbCCzUX3LuFJINjaJTPIpv8OVb7nho5xWGY
zf64TZJCT9wz/sq6FjW3tR/JWa0hD8DIRcZHbKvfhExzaCRvCaNgeW0HXZuJaPnX
6uD5HNVMjULOFAQV+9MXhLHNM55k1C3Pd1Akv8SFbPgsipxYDmFDAFw2dKd3HrLU
tVxaOZpwtE5mnnyinog/pr+BLRvej/GhYBMsdB7gFnADw20fBkK/5/WBP6pLj8rB
qrZZiaoPnp0OtC0JAIpDuhrZ63CczNQGUv2sqj69+8sH+E9ao02PuoBgbcB76dDC
Wc6940HBzzR5uJgNS6XjHkaB8vwOD8UHNk9nncTcDZ7vxHMp8wCTEFpmoLY3/T88
o1fFBADAueaqDJB+jDWoFWZvYr821t1Wr05DxYWKpyTwCIRjZ2CS/HuGJMjRpl8j
zImz2NSvvg2LkPoeWo6mtT0NZ/mW3D6pbMA5w4WETyhKSRsWmIxGBbXVRzMAU3DD
cv0V6Yj/rUonEyOEvUcjPzcqz+X2W/FzLdZqGaqwIF+vSCHzPB+AE7j+VoKBS3zn
I8fU8KVsn8O3t5T9gOMu90T3KOMOLTvfT2KXK1I24PXwMpkes8b7YiAyUsy5eOn6
luBP5e0T0hFYkRNuzsBXEEDLLO6M7n9GRv2K0CcIeHM4IO1dwYGUeAuCkJhzQntt
dHFGeaRuClbuuydCH6eTjcO5TCoDPcvFHFS6CX2ekUiH+DGCi6MU7TNQo1JcTOoL
+Ziet0VXPKeD6KifH5MM1nPyH3hOOQNALiT/AC4C9NndkH+FirwG0uo9Tl6dT8ko
juHMnc0NStz03Sp0QoHrbEtkoNFMGCKhfw/DAGpt0HY2JNCzl2+2Ndgose4vXjEX
3gotnuzeB//hvhNR86kW5xlYXjkVlIaHxo1CnDeFRCP1ocBf0Rp5n5MgwdBOJdRk
iYnRd9mPkRd1AoJCk36oeOxpIxqZWBSjGnEPBXz1KsZSS23DK1vvWmpj83vHDsoa
idbgNl/rDyCUzBw90ZH+TxuOo5EIJS1X1bvawfS8jvrl3QFx33ZQjzEBEzUourIh
/vUm/3HcLBj2UgO5H2kOVdad2Aku1yFTM1rNkbb4cubi5MppywIJ3KCjYTGIyDba
cJYwgfS/zSL/A9FbzBd4dGGsQyFvpMI9y3pr5iqbaijxjC5JdeSFHqzU9tD41lC/
RbTup6lSVsh/3doZWf0nw5/rg6HbnS6T/p3kbSnEWbP+0j3x/5r6Je810CHbB2uy
Gu/LTUw2PCEfYVEnsbm9V03ctPv2i3kcNGFN5TAQ5KmJ6IlzwczWbG6sPdsB9/Xa
1Kn135YDy36+WAeQshogTbVN4xTc7vlm+4O31U0yZlcuoS4ZFMWt84COgc45bWp9
fIa1p63j2qCD8in7cYO0bQ90erSPnVex3t9RaT9yNo7AODQ1sN3iLF4b0AZsb1XX
KXQgtsWDYyROL91K/dFKG8y0xVebgIlT3N8H6uyFDZt8g4YXsD7P6vJgtrIiJs8T
8eqdQOQffn0g0OVE8BgtdOmFL/tg8v/z9gyA6NSvhisyTGVn43hq/6Ix/OWB4+d3
YCqkxidE/PFDPmroiNrh7n3o0yYje9dXJGc9W0BdyeVkju6LmwD31FQp4iOzyDfV
kGV7RIELob7VaA1Ut2NoHLIDL09Ko/KtMoFn93b6gRiasAmqCEVRvDnARjmYSNbJ
mqRnWsDPwr0CPaD7KZdF4JHIqM/rIcr+Nx+uW0XTa/uuOfX2fbLrJ7uQ2+yi1EN9
nkk++WvFkGnWp6N2Fu30+PXnCfnCKs26CbvFOKWD1J6gYPZIztsAsSidgZJZ7/Tf
I/4fowhOCD8PjCCXebXfbFQDG+fW9lBZTLnGn41Nn1IPyNJShRc9rljOSCy16jK3
nA/SwRVOIO+bUZrb7mcu92hk1VHGqrgSLepzE89mQcriOeQq6vhKluAjAR2mFvKq
QqgHR3byGVQxItKziDFExcXSHJJvome/AgHohi/lSzYsEL4P3NwwPMs71LMX8KLs
pHs23CL/jREYv6laJPMCvYztLYRblUfEzV+lWiH4U/c0X7vooekajmh6hfC71WtW
nY/rLcORVUEZ94xtU1x0CAfyA6kyfYWMmKrzSLIPwCZoruCxFOOCVqsrWofyO+ul
iKTfH9NWI7zQemLtsqc3pGrV5+LqCMfukjZJap1nYI/HfvrqbYUnSmn5DTJpVLJH
s+aTqxBN2AWp2ZBNvX4QvY9iJfjaYhIwjS31wMiG46APFTVSH3Q5Rg5Cx5937dJx
WYN77W83Y5NAUoLJUiODb/ANt+4AG9gDFbWy6xj3UczG3HzMJCsQLjLizo/2NnI5
ixddAVYTkx5szrIXq45/tWLNO0mAMM2e3wmkc98C5no2fEjhWEhMxEtG9v5Xe74Z
cz8MZ8axbbQD041CEGleV5YEK8oiXTmR3jlS+EIH0qEWrvj+QoP3gvlAFSWBW19d
aOoY0a8fNUvqfwsGbUOGlEr7rZD5DkvQhvVYDSw/obNJJY1bFLIeQHTQZwb6TlMb
SDmkkVAPfeum+EMPvi+JPndfI1frP/21yScwVzzFCiuUscYotTlUCWUEH6XbH8ZS
MUEaVFAsWfSrQRHnSf2BBd/o+kwm4ZHFqZTxHaBlO3EaMceKLYDroCeWJwG01fsG
i6wgS5jMAXCRW4wxxD5YBQkqj0/RdFVDWO+PEcysx+JZ/40c+avL82f7B5b1AD0o
cAIwumzZFc51wtZ1vocOcoXYmowF6btmHQ+lXa4zwLtkQtCAm54zBtBUyBuYnaXD
+N9QU3b3nVgCF30Aytj2B0bn7wEUwMi9Wee0PuO2O0JbvTLko03GGJAmihRzNA1X
VJjX2R0aDDJguPbXbRGMUMejiIZHCfWxafLXjcFsqSq9o4ofduX7vp1ujNvdW1eb
X4Doy4LCfMOrFWz+atad+h5Et9UW4obrgBEnuZ2l7vJ/Wb68g+V360OGpz35rVwv
X2GM3skNaX5YdL+CAkfLD1H6m4Ww6La1cGt6SkMwcfMOabXx1wlsL1rbHiQtohfB
3mlIwqukavEBCugi6z6s2LY0uVfcafiM+tNcTb2q447s6un2RZr8eB6gdzaI0pTO
fGa7tkvWXLdH5VsakCGO8UjgngBPeuD512Sfeub5NabWE3F4OIOL3GbpuXFcnZcK
bPJfvKKsZv+fXW/ZuQhJQujT5s263tkH7SDsHa+rm2VtnEm9cU1m2VSp+wpjuUEu
u1BGsJUySH/YhBeqMYcBs/BIziYVRZgEColnX5PiXrYH5ZJjExKCNaDunJijYaa+
xwMa3Mn8Xz0KLtprUvukZmkSuF4wX3dS66OvA8LHIquRLXBnqo5HzNT1uY0G661f
/hwIi1PKKHhTW9rajahNNhaj/fQeIWHHiggEAFijlxmzj0sJkBg722g+PD1eLBze
AYeNrt/p/kPrAuQmO7VxJXUoVn+PHl5Wat2RNKA5Ve5ellcrh5afr853+wIckJAi
ngDhd3ePuZaHpaASnSpiptOzB7op8XPF8ZHHMGJVSkOmMxqxu+JCLpiGm5QOqfhW
27/JznyPt5nZCJzKhRu9K0iXAoO4Qe2DgCSB/oc7/zewgWUj9XCSGJdxT+Zr83DY
35fl6CgkwNuyFHUv7rVLKzB3HOihhbcX9KBm6Iixd/yl1h/OT8/ot0QOJAw5wzyH
ET8di7mxC3bhACaZgIr+ypkFJuxi/vYIw0WAxZQiIDKWdG5qYS0of3C9FAg63oWp
aF1t9mGP5iYIbLgwXtXXO5RulW6AAI2Dda7qfTwXxB9oVW83QtCRy0WmwOCamiTm
vrfAzDKgEGQt3sgJVSXPchRrWTZHpa9VH9jVEwAoIdpeWLAn6JYhjG4pfS/LFM6j
pjkLW3sIXdcblnnZBKV/MCA1G1aVaRYz8jU7ETABeTDvrEOdUMZNPI+ITXTBw3qm
jTSM3Qb/TEcRohpeeYIdowwPj8Idage97UPvFCOw2z4/nfk5fPxjLOA9VtUZU8QB
K9vGDa12C4e49AJA4JMFaPYNGdHpXhkMmcgNdniemqgd0E5PicpW8ZmjytMwuTzX
MrsGr7wdc16nZHlb32Kccx26Nwih9ED0omyLoP2ottOGo0RZajQM9rYH+K/ATyzf
XgSTfxffLQxAROFisAYUUXRS6qPIHXTMkzN7J9EppFC6mq4YU4zQX7EyJHOppEhB
4i5Fp2EiQVilqRX0FTk/nLOp6kdlpge80XXsWxqiQC1H551FkMrR/ZNdQEOaRg+s
sStLY72LqdWdbrejvzVNEox93jIDGEYkSc6FPSk9GzObjD3oRB/TFzuEjfs/b81Z
+DQZ39Vc4zaPxiSd7J21H1A2EVemUKTTw4dncGQ7kSAC+cMkMpDn4bQJAr0+7TEE
+GDYGve7vqr2Tl43HWVd1cCvFA1Pn3v7bLI5BonDK7GBrK5zeKdcACK7yBfqk95v
5An+CqFpLTJCSt8UAqAE5KxKu5AU/oiaakFDN77HEMX5Wjn7zekBS1sGWcPKuddA
7bkX1edu4CyWUytmPEKG2OaFX6Ujnca2Ae/2Dpeh6kRSBWKMELXbx4muvyie/oO4
fJUGNHEez1hzNn74BHEs32Ka5bZiS0Q/sOX++osevUI5f5OOPrNnL0jP7h1suuy3
6h1vNFSKjXUPkr2Ho05sbSA/HdelS027lAdplxVp/8t3dWK/4j22kDnDzgQnqYU8
phBEqqbKe6hbYd7uoYQGEFy4xDg5DD0ASv4CPhyYiOQkcy0YKew1FhGIQvrnflEI
RlbTh0qq//IBSFbZhPRSBmDMbUXGn3dGJHqhuyWjx9xuhbqjomAG/EPcGMk/I3r8
whXUHeQZti9YnF4cVQodqu4stKvinDAegjfpZ9dswejYWvYfiTOI8b78knN7ScKX
0TBR2Aj43Fn+xrWybWw5DnlbuAktkimgtez5o8OousKRtVU9rC9gjre5dULzHk05
oDOanpvYNVSJC6ZEWUdHWaQBNZ1Y8JSPmTuIvh8PE9vTZY/7pwyikP64iG4He85U
6MhuZ8ZTZ9TiyAEQGKhaD0Q1+p0dXcKZClvpAjTwKL5B8caTsNb/ox21j/oSBaPA
Ss5smwhMQSZR/Mk0PmvHigvNObGxlqWUmTU0OEMS84MqzsHrtJPQxyeps/iqDsam
zGEUC0Bugt7h40FSsUQqbzkhXBR+LPMnkWnVLOqKx/pSs2kjv0m31kunbAUPqv2F
lT0P3qm0UvLOvv0MlQukKI1eisfbRYpM9ucuzR3yqfd7Hd4Ei9vlYkn0giqGfD6+
uE2XF++4GBchTjUjvcdckcXy5QK9G2xEbEmbBL+QArgcNfrBSd5tMidF4RnX0xys
xQRsdOMy9/EhU6e26oJF+fOMDl4odKMXADM2Gaix+hjpGuxL5Lr1uGOmsd1pAGFW
K0jhnFwphmSxqF96lSx9WIwgq2+jzzr6qp5n1JD1YnKhdRahsZnwHk0sP4kcN+K9
VlptKc9+XNtXu/E5mMk5+V6xNLJ4JpYVngizJXUY0eNe9c5RBoXl8BrBnwzQWHCm
5liZk1LfMPWf+fyT4RVrZLBL4ovEVVp16mUtkmxbHVJSW/aWWMjus2UAToKRWe7h
fqWn7WEuWXt0/3NE57N3NaD+bzhiP7lAChErUhPzHmCuwkq4ISZyGMugtTy/6VkK
u0NZJNIfbw5Hfb/ktc/KgLrms+uGVZRTN5+HXKF5v3HeZoyWsznv7+V9gFyoxYDU
hgto7Yqa6OxVhxD0obKqvwESPK1mrD7aaLf6+oPtmZpVJNDMFbRsU9jFT82gxnew
o76FsgpjSBlMZGKVDEdDOfeg61UWo3rIRBqba0P6WiBlCrUr9nLvbF8gS9yiIeAy
QqDDvJM4Ue7vN4bUZYBcWR0cTmAby7nRc1BTjTG+CJSlt3Jzn3x9wjMX9L/dfSDJ
KFtXVSahaqJ/v7/8uluhzFl1OREKxlGFvdwqsyvTQ+ei84evEA6ky+0gIepoaugI
kFZKDQ/1T6jsriZjdML/GoWW2s6YeJjfHRFu44ecYkgJZ90pPNPM7UXwxAf342bH
kZBy8Z33e0S4I5BREPd1pHVbjXPw6W/cXn8GNCubiVQExEl7PSNlVLhHK29aVQWJ
dmIWYSPppIgEm2T8xK0NgJ2cGq6pUs0vumGnaDAZQbyJdxzq8Bks7sTjSplUBX9U
CRbYNxcx2BBTmBNL8mskjgFpEc3n9ZYgVuOtM0ptUUB3Y1opziE6VVwx9E8/ofUd
PnLB1TmCfA3CQdIbvn3LRb5+f9xrIQ644N2Vl7cJPiWmQgXiDIcj4COoZKzqPrrQ
gUYS5ZoTlg36i+IE7+tFnqRz5SylsDaFyvI1FULMWOBOAqjSd8lqHuffVw7g206i
UDp5aaj1hpw+XgIhtaGRMJzq6ioy6pm2V7NBAI81+oewOCwcpaExUbWuQML9XrGh
RhlUuZpKuiZlFU1be9YaDcoIEWAsF+J78sT60Ohx2erIc45jqtyKiS2Ui/bJpWhe
9F9S38bBU3obzwjrsF16iZZJh6j8wHwuDvkqCUl5GxBU28CrHy+Y2A3C85nSkua9
Y72VjBdwPDkjdw6OHIZKA2cOMICVWCSOppxVHOkwAbY9+pgrAfwbX/2a+9rOCcvh
MinhLgBS3M6q+E6TNWyWJIX+lnUht8y1II0rnvDAkwadQIlWvDt+qKDC9IJSblOh
ebmK8JInXuUlcQefSBVHmO3VnMhNUiHtDGXARm+RAqV44QS7ENExI026VvCExDO0
nGFTQzL3bHirnEhCXlbV5pz0i388+/CSTf9nDbMkP5duLTV8q2AJCTqWygKNsa4W
tIly37g5vKu/iKYTg8kwCqe5xHrsueX+svGkCSoktrJ8mg0hUV6WYmii5Xk/N6yr
NREaWMhBp31XkmJ1dY7zuZluW8uKLdSmV47iMX7LiGOOslQlsxserolSRbsjHJmf
JL9ITVXWiWsd3j44ZIC3mAQiJleoCdS2f/gfpc7IDHSBrDQbHlNwn+I4uIN5huih
SyzgtYPcV3m7KZgW/dw0m4Oo977Ub7I2BbpEvR2NcZrG2ad05OShhbC9MIL0kncE
JlXjySWREOSOkDSZzFOw/83W9IVZqqpj4wgqczwcpGnArGOrdEa7Z0KiL1HN2vA0
ZJFVdB903WDWRPgDVAYx3cPsn6yjt0DY1DTA5tS8gP2TmwvFaIACSSLeSF9hAYBP
4EwbFFiOq2EHuUyRoiKLzo4v8PQJAIxbf7uZnGtx/sySeWmaCaKOtu2QOmCs3MIs
FxBEvYYYkbEB6irRTShOh7SO8/0nBO5wheMl9dFumumBdRewwg1DlhLhtHo5z37B
yxEaT5D9OxPfd6Dhbvgi8eSR3XlkTSzEBsgSuk+WiKpSadR3B5cx+EhcIfZAaWWS
ghSKxndc1B6jcU8qNFFF8taCEh7H2O7c49tURkfwZ8mss11kndhygYgzMKs0QihP
t/WXIQrZZeIV2egS55tbnhcfrCQjHrDbdP266v58pFXVSVsjt52DXzHhA7uvBiu2
29+87QZodnG0n72WGf4XBMpj/YW3yNCyiyoUQveFVILqh+a35Wv6j+jdLdYAGF2l
Moz7GU0ELxjwZZYveyqtiRvJLHKtJTYHdqdtvniafRDatwjFrRW8YYIPtruYxH/n
N2/ddgWfLmlxPBlQLlvWeDveyALnnrB9JzBL+AUpTh8weZGV7cBcZu+cVvM85F8w
CJoZI9Y1s7qDj5MnnkiuVo9vH60b2zZ/t31ZoJwWJMQqpptiNYcXSXBJOUuA4ciy
TQKmTe/0tQpHu6hJvZ/LgAqARgFaPIZXM3UwAobYc3Ch25spPnyHEvW9Z9dWG3Cj
S7tUZw4cJNndu5jppD4f3S26kmVxt3y2Y56SFa4IhbvpJgXa6LL+2Mb9LKMVD7UM
g/2I9k4SzPpWgFJ2vHr5av6fyJvO+SI0zRm64VPQq3pOQVmPlc46ki7oe9DKjX3T
5v6poJxJuGGqMrUExMm3gLf01I9tXSDQk6HptHzaRrRhZOfWMLOarQCs5lZpDrMS
R3yfFA1mACfqUtcgK1rSS6VNjp0DsefdnxSx3LYlp/0OWehg+j6iXnCRdI0uQ8Jr
+TUwhVZwz9KtEIQrTG7M3SCB40WV8jCZw7wDq83hNeALzNhgkjVC7PxPPJqPBVf/
E9AwzybRHK9KO3SOqjSUlVjHbUJgfPhPRj9/d8gONmFlcYSQMikD7iLjXMI2EgZH
kklDeNpgN3FIqIJRNMCOT2h15NE9pH2CkJ7Po8PkRySL4rG41KZVoEy3ARNHgfFl
1hY1Lqdktbc7m7exjBLjA020TbLEiIGYX2a23An5+3napM664BbAmVH7C74k1rSy
fjNFKG143vY4euZLu2EC0OTbW570JBpjT+4SGJ33+lTxB2AA/Apeh94ajyzgJIzQ
YWD4ofkc9e9DOV3RNsYsVameFEqh+EV3NhOBwxnRKDpjXaYuIS3xQHrtRzdtie3G
8MHdDUHb/hxseCtb+/lYFjQTjrbc23tzdmQ/Dt8nRt1hwYQXcXzekX1rQzZsYz5R
hfSveNeONQ0eaNweuRzegVQRYcthruusI2PaVOcBs3BdewGgJU+WVl6XHE1s/RIW
4Rk2ag7gjdsGvxUcDn4WluOh+D/VfhUSFx8BzJQ8jVJRhxK88iwEkarYBt1zlJjs
a5sfhy+77q5p9o6oPhL40nBgjQSF3J6ahd9Jhv4FIiBD1IKxvxlP2RPcZa/4F5O7
qcvsdoV377UswM6Oagn4js1Kd0RuogtVFFOkvqibypNmo3DjgrMNbINeuRbTeFLE
YcbJ5trJdQHqboEkKA950Q2X3VcbB1md040XtayapK+F05HslhK9kB1SMc0OsZlq
KtF+l1A6igqp/+f6EQrQWyqfGebsEoRN4DwCX5pCJWS0I2Zbl2Q9JpJQ+FwzqPmc
be9WPQExUpF72BFigbRVtNABYNziA99f7MYbO215embyp1CGjPBrGogqCojEhYHZ
AJoAa02AYFo9pyK3hi9YpWV85xdbfQVg5y6XoP7cPA0P7Rq4RtQ3ELIwqpjjuMDa
6srM0sN5mpUx0hc4COrvkq75erRMQK9othhlmz5opqlPuNrN2EG3RQjTIxbV+832
ovraIHF7L9XG0AdJldJ8jvXDB/0MuVUqh98WhaQku1Cw4nj5WIc19D+O9W39LJ9q
24n8QWJYAwykE6Fwmg4oMQfcMbWsAjPwfRzqmPZk0BJC4eut7zFzfwtDXu9do/ut
ARo6h7MyrLk3GVlytZlv8QGPDwHuHmQ5hqtfDSSX0YJlqr8wn9gdsB8Nf17Ao2WA
KwON8etTFxYwfGvTRHCRKth1F5JsGnItH4UpALVYomigLGWeNxMcrUkXYqhHXKtV
NoSYEKZswZcsP1101qlECkONDbsagGlquNpwdQ1cu6UO+mDyKzE9Y61E9Aee1OBY
wV+eo+W4ahg4OIfKafmTyxmcu23oWLMxccdmSp0jxJic0atJ4BoWATjPNokkW3m0
YS1ErCoGwn8XRRRMGKqCS6buji5PZ/uTcbH8NHyRCD3s59SCK0uQdguCGJ7dRUoI
Mv6XKhVDhRHMgMbNoOgn3Mu6IdOe2q1ypE/D8RtKbY/gwJjhwQuh4BXHt9EIbBVT
T8N1zyuYXWoEFPAW3gDCYnXwk/JspGkowIRr3RMuYrbNjDK7+JnZViwqyCq3Msfd
946ooKfTBaWGZ7Bto+1NIDU98LAA1ss71BpjBY202UEeRzq3UqYa6WqDwbd5cw8T
6VOofvy0sS4Dqi7nxutyScLEzh9VNaMv31Xge60vDOwqP767EXqCYPNbTGBbxs4V
BNtfrKlQfWq9HpwZ59rjaVJyyJqAJsLcbd2/W3ASAAxj4wGb1lyQ3YrE7QdHR215
lBIZoYX5NF4R1C8HqEOqatmqAooNn26OMV2c5W43/ggO/wnL02NfTelQThkpx5a1
6Klz5PXwX9e9ZJ7/sfP9x+awMvM3nYzIdYVyVCklPWrsPFdKaVOqjHeX/NFa0tVE
9X76STQmitEsQerFHram4ogdD8nI66oO7CB33Diw06YOI4P9uOWiZ0R6b6T7zcwj
JsGXzlbGmxW1DNc4tFAzPdseJ5zpakchU1pncv8JcevQWrp1ta/QsxcxfcEPVqUs
YhuotOESZvRvst+aaUXD+twV3GWTUnKa+CArUWtJErN7SN6xkWhtcoVQc+t/h1m1
j0cp57/WpIuE/H32y5lEL4V972WIZ7phvhGOZVP4sB75LeLPeLb5Ql3DQn64sYMr
W2Bre4FZRrCflc7K+KMn1hn5GwGnbYfJsnKZmCXNrA1Ea12Q3qY54/G2zLYSTYio
vsm89wje/ep9H4IM1GAqbHsMI9gxaQyXH+71JN8LTDc91wisae4rwTdMQqk6ZFoQ
aR4J/T3zOnquL/1EORy9+m6I+lgoLWUKxVdG6w5TgVldRWIsztzurZrwPCkg0aJZ
7mbsNAvR9HTPcuTL4sd9SLFt8eb0z+1miTQp6Bh3gtaLNBkyTlgQhIRjz8I+vArA
0fUUDpgk/5+ojgzgBovknFbsUeyitor+WX9x+/0qBFiwikeO2Ii8mpT+QegdPQcI
hz/vag6LK0AEZLedNi6thCR2EJtoUSuT+IHtHcNOdZyBTKAmkVk7Scd61IewlJpE
TULaYrABx5DPc58myd9RJl8QIzp3XfzCwsPrpe06mfmKVdkKRZyU3KRxHsds2aRo
nbeMp/IBM9wV1SPHkTbUIDjEa6bIUK2wzLwBc1Ek17gxjI/SaMh4WQpxHh1DqIlb
8bHl5u4DrAyPFciAJwKvvafwC8GTtAwZmURRcE/KLpLT1E8B1qxgy5+SCx5Vmiv+
wK3Yd3PnvcXO1Uz0DilBWKejnY2g15UBCT/ZIrCJDawCoEYGAPzSOP3dRJ5Ukutr
8EeS6xODH9XBMI700rHveda/a+ZZG40t+UVMMZBAiYRJAduGDu/Ld3jBtFeETcT7
lNCXbpGeCSPmbYbydwwPEzpwmEjEUF3kaitYnKq8YUW/brOzJsCqR0FtFAHXF15W
Jh1FkIfvs26ahzJFF7kfcaYbk9d1pXuX//Qzu33xPetinwZutgg0QqF1qlxHZKN3
6vMdCyoRj4mxZ3wuwdY8BIeDHH4e0uqAfmCL4mL4GcyFYf7uttYANw2iySIGNXd4
FcSVwjlJstSA8g9Z+y/zzbyuqPFIyJ9JwqdDW3FmD4iZhkGCFcXPmzOuCAjvLv8F
rlZBiocr4eLA3Wof/lW6p9/0YobokOneU1sTH7C22KHG7HzmcP3mq2lFuEk6ghvv
hYaQZa25L4vS2Ef5axQjLHbKq8nqYIr8xNagDpd+LfhklLAkA+ev1j5ZuqScgCxz
apL9XGtd0KRNQkd7l7ow6ovv98tGRxWOLrJ6T3oqHHiua0c+JrqDNBAJF48ZT7d9
Pb7B+DXCI3fMIB6PBjojVVi7cbl+3tKcYUAJVW7vvbQGvPgqkDbD+81VD3+0DOYi
9V+CTvbx+SI8jGJW4octgNNiMGyp3G4x3h/OESED8QxMRpuYxVkVzXZUFQV+RqyE
E3ET4ERTRZenhdFgYYi06/nHbqyVTWYxv0cqly/xZym/1113iPzNzC0XoeMXVCnH
AVlTW39eFWpm9SpJY/P4BvsZFz+fKBn5t/6M3lVqB9J85kJxiMK63gg2Rx+ESu+l
WPpA+sSSZ0hpMgGHGEu+JbmjAxNtzQjJya25c6Htsy0v6V36SWSXuItLBSrBa+fr
P+ecQ/yIJMnYlNTVn13S7dG7nNuvldDEvkRDECxvMYzmiT75TSnGtfTPI8vQLXzk
kau8P7z+X9woWX9FlxvUJRZk87+NaFIzGC/TXIeBbrrBZ2k0GLPfHRX7oWEGtvsJ
wOdStRjziKzxaF1i4dhzTaHj11sBeIxxO1Ac9MN6NxA2pmOdxQEI5et9Wd7AKjY0
m/b6Q7v2KLHGbE7eQ9IwlRQBrSGs1JGyHaaexAb/gHousSnYu5n3kpcs5yUUehoR
9//TcrGWTa6DYFYWLEIoEXQh4A1g0VB2VYVg4ZnvwrW9pxCG86yTiBFUFwZZfp5A
7vrAJ2XcOBOQ0NSekLtyYSUT24xEJ707K/IzOoVi01FCrH0qVMUUMxdU+1kRlPOR
+8zGDr+x7HXWYc2AcYTaCYJcZC3ktVKUGr536X91RgItPaHWdjDEk4Lr7fYrLkaB
sMqaBwJ3EO+e3C/+DPFTWT+ok4myD30bB33ArCRo9FaMTKQcWGh21kR1c9NBsStJ
Pte4XlR1wuZ7a+yNxcrzit7ut9bNxqSUN7yIlPL5ueYHoysMtu5gy0/x3fFHOoeM
bp6vhpeGWIRF2WDIbP5eGXBhdKknQ35Q8iBjwV9i0awCnUXdxy8y0bPbapr53bOH
thpMvxizCs2fIS74Ck4CdNz8n/2jMRXfuAQxYLAHYEecAIdSInKyugPhA+Nj36wx
1Mq2F8+884EJT4djrOeisP6TDUvS+PurcZT2njEHxUuLaCripd7etcB69CoJi043
hsVDxSlRrWeRp2NYWjCE524ni3n5UjbPTf9Y9O0limBeo1F0bt3K47/QBrtgi34U
gW5EiQjApXjSfWf2cPrp85gmuoCY40f3Y7VMNRH7Wzt79ecXas2wwyFul6eCIHM0
7f1IyCMLE4ka1EodAAXmI1DtUv9Nx5KkyFbZnSonouP/Z7Y8WtxqG/3lIMfsd1py
iRiW1+88LKqjw+sr0OXxyDMnpNhMRmiQ8GGc9jjC03HjhFe/62pIVKNZ8Qu7c0TB
4D03W6XgEtfBcuaHAIbkeKzUoAT5Gn7JH0YtJ47FmClf8EggNkZYK+AY3dPxzSuD
jhEdO8Sf0EpGQb0gx5C/a+iMcLyCrmfIL7oWOUZa6SwanhkLxn3Ry30bba714hGd
X+v9fSkr60aJyDq4ZzgWIt42mS06qxOMdHXuQoZl3pnfLBY3GCQcmEPRBTQM1FWc
Lgrs6nLVmpX7Cgx2+WSBRo90fZoWxoACEg1n8VX83hKyXFWStramSkz5Fs6K/NtU
Cpv1I1PEr4lb2tsxMmXuT4h6+3QIwhWc/Ya92JnSRors+T+ZqS5AP1jT/7WiYy0w
IdfxtKvKt2iIt0VnxC0P58TsVnXKPsak9hTJvCi3Q72sdVfUTs5F6YdffTP5GDo/
lprU0FxaO6bYmibi0YN/uumcu7TXwjkAJQCtW2sHaC5LJpEg7+kh564JMpoynNbI
OdjOP2wXgxL/FPWlATLyNduFDXhTAkEd/ObT/0kKwN2wNMvVAuZZiqaEcCRWOol4
Y4n6n5Ey3GtQRkzqSwg5hin4i89FoFlgw7wfS++ucxKgzRp5Zo/p9ttvUpjbAtd6
vnCuzhZWYXktPe6tnk9Y36M2smIwWvCyVJNGnXdwIB0zzgBQfElw3omRXdY1B8lW
hX/oWwAMXkWpD7/2N65+bpIppn93uldXwZbKmEIzBI/NCCWzChLO8g3qi0bOK/Os
2b8j4tLioqUCFkCkjNFnS9TJPOg8esjCROkUO7dbnf/c05TvpgABJyHSakNW78Dp
uFs32VhQSEfRjTBrMhVkHv8kA6JXojMgxitAxdXvef96/bsJXAvTvbmsJcUTtu7b
GB3d+/0m4UIA5o+aYCzeK7jgAg2bvPTXlLTHyGvGjSsXFPVzWK4ELcpnQ0vo03Cu
BRHO18bndrww4AHV8MFBvdMeGgPNh07YTJiEPk0rKJPTwVAsBqmSgIHebLCffYw5
gbwG/4TGepixwtY3RAH3d4G1ORwPAUmUKp31IvS5+0QdLtxJ6S7Jw9i2xwk46KOh
gxoD+Fcz8LRylTLlu3IguWiiQ0sQ7BvbQGQbI6jFFrCOyn/iv55JNNVguk7AQsNa
SrujWmloxpBzK03vmuT3Iylwx/v0Umf6hFQz0TALUyRp0aLIeaCt+L1sMHA+L+Gx
bqjzB5sPzO4OhwbAkx60ERNMMHqaLNCgfwPV67DckZzb/jeuUHJFqMjHPo8toK0G
n0wieRfv19XSMYePhGez1A/HB7bGxci1LJNKC8HYJ+7kkN99bDKsL1wNKYYHqy/f
iKHWNtIaaEf5g5NDox/vdBt29moR7e2ok/eEOsclOLG2IlZel60419OKQY/RCrRT
CUfMTCgbpSWh+IRdsGmEJNPYuC34DB7Ca/Qy74OwaCz+kSxBFk0U2UTPG6Z3jByP
Y1VUXvg6cx2h679cANc5GLlaxZY7HNWSh0xRyvc3Y4Ve0CZLVZ+6KIskmtyrgzz9
7Hew9RZh1sA51eeS2/snHVqMgJq/BJV+fjl1NvbTJePsIl3pYKXXTF0II8r+bu93
qxTT4hHNrIGskEW77+M4Pqvj9me4iF6KuvCkFBj6EnfxSCyh2T3NuMrjBIrrd515
i1TPW3AWhgLpgpz3IPVNaKhgu5+l7W49BmVY370x+jQEhZVSwxYlWHK+7na5Yi6q
Jj7qIUZxqul1j5QoxI7kTq++U3RZ1nycavahg2TClofxO/kAIm+fkqei5aq6SpYL
unViQ8uYpc9PHiFE6AKDXJtWrtU+BerH4CtTBcJOSNX8iskGsmIB4vOC48nV8hJR
v058AFI5u+68upuuvSZD/msbpecw6dgHENl4TaYnxrokVn/mQ1vKjkw/2BoV6hjM
qduBNiujSidnDNj05SkiIjJ6jc/vspIELvkz1QLG9PSGyM7XnGJ7WxCOIqQiA5Vd
8fvoDRQIriWeSMiUloOoghnmspcv4QkepYjPf0fGWB+d/w38NAakxpCCQ6TCs5GA
8tbZiLnVs+g3SMNVSmMv3dTjlEnMeQGD3gMQDsq7Zo+pVV0y3bdATVIjoWvKey14
5oa/fUVs/B735kiIY8UUpENUA2q5F8+JGzLAF+hbHSygV+nhhy6MsM48r6j5s6w8
JkKBbV3JMDnENUB6+q4MdIUiOb073DrLlAkhEIaO4LPhdv/PHBxzWtARNuLkmzWR
ssEPzPezaSxBQ1F7pln7i9eAJAODMUReAy+lSs5MYOmbJ0LQuaGuPOhEDGJXxAUI
3JSPkl/V8netU9owOH315BrERVlH1ZepJNv4r9k+u8wVdijqbKicKcN7H6EAeli2
Ec7aDOiBae8T67ySw0+KwW8Kt88/dWkQgmNOsnOSPo9CayPusEDZ4Ze/1pAhLuN7
3XZlhAbslolTBY+if/ADJ5jEM7wQryrurLsULdg1LyQfgYxOThBjnx38qVms+VMP
f4eHXmhmdjG6eO+TZz3lJjr61Rauwq4QlRCFD0Xfs8McXkTm731k+guPfbizsakM
8OZaPeJYlHa2p5uFL2JzLSFjtxFooKIoSqjENUCkcq0LB4lXbBmK02WRfk8cO6Hc
HsO5EbhMgqLeSOlmEt8RWTJtAhiS62PHnB3Uwn92HFDPMJWzYWp65p/dc6ROBFQW
UcsRSXvwnFpmVz/fCG4LYt/LvKVhOs67r50gScj8QJ/+KG8Ha3kmGgCUT2a8ZLmY
00xIV4/S7kNBpcfWoOLq0M94Jn72eKXcM/eavBSXJTftcFMf01iSLI6TJuYzjF9l
gVnBrV/6XYxk5OFe53jvXGxv8yMSOpdFCJNwHuWt96ccLV1kzZrmTEpBqOoisQJ6
r+9XupmNUuBiZ3JCrZ/Y/+pAWZO1F6xOUBHErPrmf3ei4pwZIZzk218ICHqYE3/V
Z3SbYkjhKpUF60CXC7MeFDkGRxwtWbUOl9wUvWgt0u6tr0P+SWR/AAYcWzJBaf3q
bEuWb0hAlsaSDhcZUjT/F32SduicJxnuKjvCuZBBX5QUwsL0y9YjVCRPAOJ94/FC
eOjpWeQmXRrolagcxXngqs+CwkSNbiUHzXdTv10AAE9PdqoSRWf6vZbPGsQeHpUY
qsh+PR+r6oZO/YphZowDaAINJS2DpM96iLEvy9qYB0a6q2LEpMSHPXcJV3uD0ERo
JacEcDg10NDgydy0LjAURwUNFV5NN4L0Pb1db4SyHFr7iW2yshBPaGBiUSZkfva3
1wZyVOCXGcF2tOcb4kO6xteNnLZnDRFFetR/Z/4CpCTwl26Ibzlgz2uJ7iUsJsES
vBravioo/+NKUHVTbPPZyhTzMpC80TOuFXbfBVmyWZ9yMz8UwcKUuLrPmwK/Vl03
nNqn2LbJ07Va+heQXfXKv2f60aYD4jC2x7M5BTOekDY/AcsInLMEefbachFJYyLq
vIi7Tw//bClWj7uhgvO6eNTOCJNvRLR3Ol9tmjC45rB0Wxro2YVsa8BMR7K3gWvy
eCvuSIxqBW18RPH2cD4HDK7eb1fc6pObtzMXWZJVCVvK1hyQdtHg6lRXJCrRIfSw
TM85VusDj1Cf5bxbYwsSR9njLpFKYHbbrrQ9JEwgf2tfQRVYl2/idr/LGw3UhTUS
DnLxlVfEuSqeOs44QFRynokpSLxoPUMU6leT4C0whjBvoIJZfLid7ZnvfZecPGwz
d8RQ8nNO0LX+W4d6csCFcbIuD83y0ArO3J/iou2H3pTtLYtYPbFON9x3UQEmzpPD
4fkZX2G/PvXcjocOB1TJC5EvaDA1FJgvSs1iLssds/2H2rtp7ZKkV9bw9jKMDnfI
93uDt5Nn1wNs31tC4C2pI40K5O83WwQZBSVU2BQnKNKkf6HhJj718UxstO9ej4IW
4ezQ7QKzzlb1V57uD4ur8+rFgvxpU3FyP+2qYZVPcTvOKDhqJ8rxkrQFGOO6G2uA
AkxP9RhRpQ5K4gf8/R9P54c0xGQm6BJmog1Qn2ryAPkHlC8p5PB6yMeVGnwjsz4D
7zo7+KuHLNOt92sXFIQyK+QLnbi3GnMsQhwKBWhGqKNJ6eVgWPVb7b8Em8Cbc3wd
bKhfiKL6jmyMz0mtNTun0FzcBLvQVWhhBRT78rnKAa5q2pviBwOPkct+hcB3MQsR
qtzrCFIw27HSL6J+QrjARRTgpR0aunmL8cMXWmiK/8RivrPf4WOpK9SnummPh8B7
V5CF+HR/ZNF8VVKnIkdG8wmr9gxUzCAF30uDjs16GvkWlF1/PAa+n3jBBHOif+AA
k47rFBqKYewrZ0Hiby8FgaVZ5MpPT7g184dvZNl5Nw6bgXKKhJ+8jsUcDhv+WODL
FBrqCIvJD6e5CwtoK3Afeu7atBcE37U5RWj5gUxKe2IVcxFRiVJd15hzSabciJj1
g9SqaqJE7kuSG2ktl8h2d0Rr1NxPueoSngFB1utKIfGU8GQp/2g639inRfEjTY/7
cJvhNBbmIrWRKq9NiPXHGT0EB1X+R7DTfkubhAPdU3RPxms8ViMnJyxOhJcccVhW
tkDi0MRRW/t5OoDrnqMkDZ0l601azDvMb1V7ZVg7dRI0dW+xQ/gnkqiAQpq149IZ
pXniAbbvU6YmlAHje/BVtD7WkJ2cDp3Pq7SRCUSX7CH1bX3JZYGWiAbQilQwOini
ARXK6E0o+IWpXnbo4WktUDGWogsUgzKVOHFdHQRZhZQfXekyH0s+xnZI03jrvaqc
POULbkCZ1x/LQGWpXpYEzOh0gHw4N1ws4YmweLmaV9WigsV3dbT9znpdqwOROYIC
r+q3AQERTUkVcEi03/iXxhvgSj+Z6ArLPllzBxmQD2hXIp1nYMi1z0pbMHgSxTEV
qUBexekikwdGqSRak4Pc5BLseNyqIOXIg8CjLWCJoPaisKTShaTrtbt+jvrsY20B
TxHvGqUHXDG+zF7r5DvEJKvY1Vrg3OQ9S531mwpwkBn7afxJ3sbD/BjAHXPux2wp
CpOadMxrx15QA8ReZavX8eo6S3s1B+9h7e0YzsN5IyaS5cftToOHPyr1R7AJzf3/
TSwFJzSRsLCT3oke1Wqa/E+Kw0v+MX1RyYr8A6xb9LsDJkpW3wXKFUcqLNi/Bv/B
vRvD2zs7y/T7//94B76OH5bWgl0s4SjbFNQ0eYsDpJc8lHx5GcjSDEC5IXIL2K8v
GaJWeVFBJi1wTKuftjX9hGL0JiUWdbjSj/P3IXtVzEEExQ71eRyw0PMREHFUy8iu
1ICycZ/Gq1nU9A7cyYEGo1ioMT6O08X67pn1qLHEXXc0FttSVhXJjCW077CatZMo
7G8z1sNIP1NL8znRR2jixzXz9I6cHCETGj6r173H2X35/XsD/m/tUIZW3aQA1O1N
9fzKDP9pxGT99xBkjideK0lBNLWJl94m5tDNwN5oNvPFKiI3tjx8AKClYRR+wMES
wVEP1BDmaKAM8p29CjiQCBYCfAuwyeJIZXV+uMK/6+6B0THbD9Z9OzZBQcTYYfjH
kDlin/QvOEKP9WBJqpK6e0t6g+sfmUYp5X7uXpKA63VMWHDTsXebYSeBkcJPh8VN
Ol8mQ5Bby3mePUOwv6ONnQBVoRzABsztOVcKYqoawTo9Qkwryhoderc2YhoenW8/
KUjCwMOWIEBOChenZ9vQS3JgvVlxS5jWNCPGKpC1rZce/8LM5WW9dBManqSwM0q0
h+Mrii4EATLpT6W842auN3ZrCzxWj0aYw8sYGD3o8FBjvFaOgeDzqCAtnv9f5T5M
WHuRPWUQIiXj2QleRtzA1x+w7T5j3wHMJJKZjW7TsHi3gWIAU0DkCrevQJguQVY1
E8FKRNSGGbbIiAGJeuPHojSGgeyR5nSHO5fmi9NuQnObbzsUOkaJFhVDDPIqUk68
mHcx4iDUiXxIPtgmxThX18kvtGDSvq6G0+l9OL3aQMAYPSEdffkekAiJiDkhYI1K
YbkA8KkeuRtcUO5zh8UhFEnHlaHW9PVtlJbdakmHJtdH56iZmn+4mE5kbGU+YKYN
s71oFff5KI6e+PQSo/riFcp1dY40qIMZtQukgK3UM/eq7ntKY/3LlMBIMqh8N8zB
0dUpiBnndFwuw7M+gPjNASM1HfpybJpTxARcwI7wMMmQFCDs2ILk30RJVOkg2bvW
RISwxbgOo3VE9aZTijG/MgNRrB9ohOWNpraHruO9QBDcPIxpW6QQBarZulRHylpC
rbY3AarQaTfzg9NUm2bb8OkZyuIevIOOdt9zXN7PhtMppLRMkgtd+Mf72vSxKxOA
G83bDd1YcvlfzvFsf4F5ZzZ7KbQCsCNBarX2YCA2T+XBSi/SNizcHpnf3EeWMBa0
P3iCvkRMlPkM7JYzSOzzezq9V5RGsZEpSGmF9c9pkxgDCmhm+xGbtZvJL++7AkaF
9QqHTgPHbiGb4w/rLvjKPfsOzdHVxa0rMn+4TomcDLjERP1UBvYa2Bbs6ihcr0aP
akBj4HP4twUgY2OaT5dfrusiXSeRx5kr0vcgxCWS1RHUEzSbHr2acOkGLtSdfriF
+1y65RYf2kaFzqkwOC+gH7ra0Dd9uEpZI6FyAamQp2t1o2DgI0YG6RUeOCBb50KO
ESW2ylLP+i08s4fTPPey9T8/mKPE4KuJovP+94ExiGP0Bdncv69G7XALDBAQbfQJ
Gz2GYu83wRamM3A7k2hBPgWRGcaVhWjqMJtkMpnL+1+bYgvVu5yDOVHPxljFQVZt
QlHxL3Hx4zj65S3tolUS1Uf45HbEM9kMvMu/Q7Iq4p/pBBly24cnc7Zj88YQDlT1
jdWqOzc3tqy8ykKPefggGGyuSTaw/8yMk5C3ACnG9E556Ja2BSrF2fl1WVQMiFFJ
WP9UkaESws/A4q2rPSyMHH/xwyvD2kDXe1HgBcI9/2dIJQZjF73q1utTQfeHS9SY
AnslUeS7gAZqgUlWW4/s9Fb6p6zWs0q3jKTLKZ0lhCwrmH7gQeFTyhEkCNqOjrpD
KIWGkZcLQ4jV+zI4H25Hgh48LnRDHNJ+4XZhKBKfcuyX9qoODs1QXvVRGNmfQ82Q
qaHIU2PjIybv6WJoIjSaZ420P32fd3ZN8iKDMCFJkE2nhfWYqjSTOJyMTySDS9Up
7cT5FentALDOyNRGNJb0Y0/cmA+lJSuueu4htKWg4ZmTt/7zLwhNDgP8WOtjyDj8
mLdbZ4QtENO3DeA7Jo03PTEeYG4dkvc/TDbNwL+b9omeghy/Gm7scjKjeKbMUhTE
txFuoku/f/MBI3ExK455bO1d6BysAsb5wkjXm/eW7Q0JIcRt+OWiiWWi8x0lFLFa
rmwo+In7igXJ2KgfZZIKZl62x/rt4HG8O7ifunDF2C4iLTyE+f0v9+cWLbzTVlUK
yJVi16+vTAis4+KDXZs52RV7Jogzb28RXuchAO6i80jp2LKZb58qWeGc4Qk8rYFP
ZZubYZfE9HGWROkI2VWilCeB+yFRa3YPzs76E67gpgd4IIV70ei5guwq/vrGaWKs
2qcIxbz3c68/ToaEmclxL/2mSjxrRPEfosApKWnQAUtXefFF6xL2ZE4xt6Y85HjS
GV3HDcanBi73/eaqKRQ/iyQuOd0BW6KK12A1CpaFbv8Eauy0k490PXEaCx+8gk2x
obbmeRCJKCJXMFLYEEY1KMYDncXZ3u7Nkq5boF9zrEvGHmfOYy6q7zKDpbPloKvT
lGbl0a3RsiNZVQaeq4wQytGQlNgQOAgImIdyrdGKxAi9eEXD6pXqB2a2J2uQY1Az
5YKS+vTn6LjQiPWfhSbWIOTM0Iw0ppWtVQcgfnbQYxXyBgo1pqDLtK3Jfj6ASz4p
C21sORXKFVgkBw2PumPx3WUEJ8UvPxJJz/fVQjPua+0jlszgEEAjNt0zA/3rGRCq
aqq28qWgqNR+UHQeDP+eTx8yOA3Ou/eKUgtPzj/nb29GnDPE5W4GluNVRY+ud8Tr
oLHiYXDXHkZEnYkI60G7YdnMk4G8/TeFCDR9M7SGva27V3vykaMXnARp7NOlLQl3
WuZOl0SzeG3E1uFF+VYjMwMKK3MRXfTt8RSyTRLs95F6dav8uCylUoKhEKxEcBOQ
h6OxvCjXq38ZJ4u28XYSydulhIKxhK12W+yl04NxxDHYMAINsFTGhfdPYNuETpo9
b+9/PANge7/HHU/9+hHyozHERZM7miMtr1JB1/akDg248epw+KzsHbAvMLpJ21lr
84QVoCC0s7tHsQmHlZIBjFqcGJsiPxQwoo2aTVzfPwQ6Q3kWJduUtXC/e2EKbYZV
tOAjZ4Hfy9+E3VoJPYqgJqlstmX2v/3hshhxG0r+MWC8NJx0OkcqSeOAK/X76wan
SpNXhCzS6J+kqsbZuHIBuF5nh/QoMPT5PC+ZFqPW6JmhHzveUTf9FnrfpgSMX/Cp
OX62p9wt1hKgtB9IEqSu/dS5ibjl4MCcQKeaj7qgh+ivgfEelzdglARkR1YfEXqm
AISMPJ4qOQs7RCfs6KfihEE/7ncRk0tT7TcxuAFH3WYnQ7D488MopiE9fYC/Es15
YlQNMdX1iH99KdRGwpHi2qTb3Sg2hkqK38Hwg6hRAivNFf0L0QOqLcs3bNiy9UC4
wbWlIzOLYiqY5ooPx6OObd4CUbe6Sg41QUOTgdi5xD19EYWQM8Ky6LMuqwRC5TFP
ojcn7uOsqV8ieiqOcbx2S9j6gCGxS0hmw1HbGPR+7C8wMSom5+abczCKCD4tfL3Y
abm7c78VCwepbSeWrftCk+dE5aFw4JyPiCmCqiiI2sQLWlpdlSOTIXKPZWVaaJYM
KNbMCqOclZd3BsFcvVzHIcFSQLgWWn/vtRYAo9CiBfPI7U2FDikl3MmdbC9NbbtL
jCm+yhsSZvNf8CjQBqT738r4tO3qWFN5+SU2M8K3/GF2quHCD4xVK9Ia47KJUKtm
IYCuOZN2jQsP53KBAdUdNwVoNOlT4yLza4lAepwI2TKXbrEpkFQwsRvTDjgFCIaz
2AYp8E8vIEFha/ULpfj7utEC4LNjqvqiyZWjEFWwMZ9kplnGqETVg8s6X5GILfp3
dWGDL/jnQWF45X101gqX/I73eEwSXpq3T9yQHGDGYscrhJFM10/iV6ITmdkq5DEy
1+ar0Y5oFM+h2BWlt1cg6RSAPw+/8jpV2tiRmCi873y/H3YoIE9vip9ydOhAnYtV
V0TFrow3D68RxB8qGV76Rfe2dn7tRr0y26JAKG4nNIALjZhW8fJG0wPHqJywp20d
sYvYmFYd/5fCZ2iXPnYeYItd8lOw8AIYUgWLUo68HfiNx+4D5DRMOUy7O1xJp787
fc9cT8Sfv2gfGKJVe5NFs6FO0g7pg+8O4oQSpVksR9Paz50i8HlPHt3kpqTlqui1
f/bc+mo4NrSrvh/6fz1taZxMd5dWwc46Tgsb4zBvUQDY1BYqUsrHqjsGxhFP3BK7
OOltOmE8/lxrlA2uNhqvuGpsZhpFMhHghTFnyfBoh1/TTHB2GjmxuRUZj7O5xqgh
NCRnHYrEhJW6MuQKX/VID/6yJhA5EReWYWSwha9LLrDOo7scHGLYQB5UKREtAGtf
08srI9OhJPv2BbEr2JHDCVpSXP3JbVeSwQq91jz+vImyHAeHyU0tMxylp3a/GLnm
/D9GQSgXA6gIdhx5s4sgZsXoaozNlOzssxM9hMHo8EzGXs6bA6TuHqBElPX0xIaG
J6pQXDAvfkcpmPXTDCO2NgYdC32WQQEK4RVRniiM+QTroBuZfg+21TmJYCO24ROg
gQG/r+QBfHVUMya1XPGJDQn9BD7aJzm7iPIF+3W8/i72NRkj3rDkbMCX8Hb+ogGJ
8gacVGXAQgc4iLAAzWcyAn4gsptFztV2RnvHooI3WKV3E2MUf73Q3cj6+gQ36nbZ
nBUj7K7Ry2A/rNo+LKpC9AxhtIRkYOcwVlDBB6Nd9I+bHhFgna1SfIiC0VBFK5kX
PQUsUGc+WxOUYjlj0FskyhfhIgPubMnGWhpRkP/1oLTurZVVVhzLDSIEHCYi1x5Q
q6MMTU0o4HeBga+5MyKImZX1anLLK0nmi9pwxaT+H16kpuS0Aya/mBxT2O8xzKO4
p/ZK+FCwCOngmaGunKIQYi7Kd2bNSgK1XRsALjyuKLpXF9X+3fdxZf9m8+P7l+NQ
T6ybYbciqAUHjQZ/auneEHengaXeTZJ4a3DMRCTnsKg8SWSXm3fqnxJX5VCaq5sJ
KXw2g0wDOCTO7mwpyoFX3tCk9s/BbT3+Xht9xusJXgbLEslTEfMQw0pyJiV8VnvQ
U0WB5HGmuuiRwOl4KGvzsjOcaMIlr3QD4Q5uSPq3JNInac/QHcxey+EteKG+SUWy
GtqaHJs8q9xJwVfqn4v428KgYTh4Y9uR2yxlXxkb5LspZ9VJ4JsLxqDXA3rR3AoM
FqAP388k0yJHJ1Llx7lhWfNiLwVdtZOMhJtjeBaBIM1uEk/gBRMFfo0XzVLMuzZs
dQZcWoyWev8cKrqLQNyPEyAkuLSesIbnVIqrvsLII0MxLzvvaNerVy1BYXWo68aG
MPhwRzb6Djt/QTH2Jx04ipT3AKjD9PNZ5hAiX9isFigH22rgcbs0clPQacV1CtU1
r8keG+RAffLnCrxk5sJ5YzoF0UZTQ0PP4My23WbAKKJlUjXa1O04t/Ege9qTFp5v
X6iNdPTlpngnkNLzgXKX4eurmVMW1pnVuPi8ZF/G5yc4QOST8sO1vRPaDwaMrzyh
ove2/qWxolwQVVP62/LOIutDAi5khpUNoEHdX6//E6aWAS5ab7Yod6vrtzE3pvYb
LKgo2nc+dgW7C5w6TMh1IwvdU+SYBXN1AmFQwblqGPnLtsJL+kaw9w322i6dDwcu
/j+FLhgWy+1D6hWhDDtoSSujW1QqHkYrdU2xIb1hjA/6lr0iHeEhOLAF1ZSmkoxc
FtfF1jnVwxPIWDnE7RLSoNab65ZuywkleTSSNrl3gPkqs2p83CccdYU/Wfkk8wHY
90B+zN0cO+pmnROMQ1GZUNR+j3+OPH9sJT3n6ZqCTaHMMjcteSXDxqtxhf7mYyj+
5NDxIt4ftFOHTztfexS+VXL+MVbOxrQ2kStMjth5VtpUZsGk+xgsi57TxD2B+mpV
7Tp8Lk91ECpH7yDp6bIN+qtFcJq2eDPSLRZyNRrZy5xsdSWoWpi1ZfPGStN20dc9
63xvjB5snj64W37g7VT6xcN3gQ7rcbzC3tLDXKXIfhnDtbAD8zqNYFwPZb/IpA4T
g7V/H1luI6ZemzRfg9pdU9UfBRk4qqQruU8DhYcvHXuUlDmJ47+zwRNQlUMwEqKl
XO1c9YMWf1s/VJVoABPHaRMG+Va0/c/icFpPn/bIn/MsBobth4e0NVH5h811uXLc
inpc+DUj0fuhMiXSb5etlWTc0OrlysY/TJttZEzE6a80mak0JKIAUkSB658E0crq
6jZ+RSh11YGvw1Zz/MND4x0OOIqbb2a+Tss0xn4dZao/OsFALXD/VE04VrLEBBto
a5/pTj58h7O8xiQtQ7xvOsjsK1H4RO6PdTi4GTL+y/gbixbquV+XCchBhvK1ZHLI
B51+9kJUCcHXUiaqIjEjvgmCQGHCgID4QM59/64jecgWLcn9hQMXiqsAAkhHWP5Z
esDRMuhxtQJAft2Ho1hDnSjYk77u03UI52MrxYAaXmd/YHdJQdNBGZVTT0nSUG2K
gfg2FzeyQcZStVxNlcfZh0P2vIG/5vfBYuydUrU6gmaPcvYIK59BJpDv/6IsV3TC
gmZwnY0f3fOFp8eofTn/1n4NHY3Ws9ppq1FrdLNungfyBlJpVo7a8bT1wSJE2vZx
aZU4VzTZtTyYiTkxu6YzyknPNai3rZQ9xjjzIREVwHYEqK0OP4VRR3meNpYZ91IE
kX26v5Ibdfrl61dQv2y2RttxW4HCUpFSaIFYkZzuYXxj1Ylv9X8mDQ1lRGf/+w/2
3LmqjwiM49oQQZPYsH7S92BjplA9JYmAx07+FHpWSxv8yGDYf7TOt8jHnTK+E9ow
3OPg++kkudBGpzT+Qvd/krZNZpzpSUPkO08hpTaRrtpIqiI/NXEokv8i0IMGqaSc
HBvGG9Yf0Za0Vymhz5sOR8mVDT+ElUaasC8lgMBlcEe1qHcZ2r5GIFzZf0FZ2wdx
B5c2DDf8eHFx3+o23hzQFzP9snp1bHHSFDvTGNhDxib34lQKI23GklGsGa+pq7to
NwdaGeEOSv+4JszQHbpkCY9J55cWin78CIIWhgTOEoNYgQH2WwHnCJ1SAzdky/h9
h/sFakS7aQ2MDSoQWbUs23TRwzhqoQXdv7QF+i+KzSZQ+lfOMrf38AA9ThaNcZ5I
sCPllic0WYK8ATAtOxGLAEMHJZGeba93O229QPmI1EoE4HhS24OMmpb6h71ndB6i
oew0VFXfEhEDGFqzCjvjq6QZlvSlrVBuBlBq6G8b0CBbum5KVH4EouvD1ldiTZeV
hw31jSd8ZK671P/Xwm5INOgYhVz+3qkAZQfFBrffOqxoiK6zXFcnis/1TSoT5+Mf
3ENnQxDVespDHZjuYCpEDMxUcRXraHHGdkrUeQ4lpfST/NCMmKX2cHZbz5GRCFPQ
tRP+yM/o666Wf7PrWLBHnx1ojbqK126IiB+1Vhop0LKgI1qwn+/6+s4gVGGj7MgQ
oBCIr6Dgy0tDI+KZTl3w9gESSuK0jc52PlBSzYgen5GTA8V6qivuzeZHFJsJZ0+l
B0Pm+7N50wvhPiSc7jZF98O/7xK5SX+nMpyXaOH4ZXRtZtq8XVMWy5c8JbNOVF5J
gjIHhuRI1P6X0IQMuLbzRq/7WM0fZMuDatimZvGiQanYc2otbxCMs4i8tC+3FzmN
52VVGFEaDoFXbylNS2UXP98BpkDEeQy9SYGDc5jlbXRGrKCWDsElywlsm0HlT+hf
EwEfOiHqT8kDvS6nydmF7LL/fDcdtOohJjs+hx26upuWqaUvrE4hRAE3WYa61fsv
V2FrSFjupsbS9oytDVt0PvwIdZKgQ9knK6yWQRy9hDJW6AMrIWOXLHlYbHgd5lGT
1SphtkuMPvv06FDsP67TlZ0L/KzvW5w8GTVD4q8wp5LMZNxh3vhEM4IfAaIlNCyF
2N9OJFj0SIS+h4u4pQdvnIaGKDXZkGp2iplK4fbtTq+Cv+6A80z6jC5pCkVORUNh
I5RyVLJtE7Gu4zANBAHHcA7ifE8AoO4CUHSGN9g/mX5XbdqDoXExkWrIMqbm4KDx
YDfyrdaZivfRMvJKvRa/LjzmvRGVjmV54DsxA0um0i9ZroazZ/x5bQY0JzT8DROG
q0KfD7wCZT4RyObtAYW/aTNqp6CoeyURLlbfXoQks0AoLXe4nifUKUh2vjVNISkg
JwvpLOD6gMtrM+atgwt0MOhmb1SIAzNK92T03MNbeDrgtq1j/tKJ5wziB2Hk77DC
PydWiQFtoKMyHxSQrll9dmjp34naWXJ4pvJQq1cOcHBa1t9tJOdkuOsXrUm7ud95
W9YY2ifWGhIBd1FBQ9PmCOm0wCDyJ839zErH0Mq7bA1pEDyAoMbI8yVvT/b975+s
YY6K+dDcs5Wd4xnI8iVsZrLszuXgWI+Yl1L4Cvv2rYJvMikjroCJxS27kit/N6SO
7cjq3VdoHD1VST0fNXhwy8SIlwsW4PuWMOt8POet7cGbPZRRHe/W3bKTyxrvEKkf
iRIluaQmpaFGRP0+dVsPLEVlfRu9zAZyhnoofy5cCCUx/q6pXAlGgs933J7chm1f
x57aPhPjknNxvfcYGuScIZ1LGo+ZLOwYwxgQv5TTmxjKK0S4l9gxO/x3pv74yYi2
dPuVLkVpdvxqEMAIXhKM6q6uMMwGUJSUagqQiDKqGCRgPmI6rMyyq8z7mOPsptXx
Nn51GGaXn4kz9HeBQD7fuFfEjuQ+We1184y28eaTUo/9JJ57M/CP9Q7jbb/FSl0i
urWqmTp+HYDizQaipPmF+gxJrJ+ZnNXWwLYumaJPj+OOomgTLQ+Dy1BDMKr3qDB9
pL2RkHAiInETJPI0SKnAYCWpKMUGsZh2n977cIBwEb51zeD/m3AJJh7dtWH9mKVX
yqyi8j4lFaMBVzgFSfFF7wi+xwePMEWyxABaDdtxevXyoLSDPIH4bwhir+msD7VE
3FYEJOJcS0WZxPh46478PZvd/j3E5KEO0Ioqcq8MpIH8Hy10bN8PFDBJMx4skg2X
OZUBjiBYpy6VKBzNExSp049caCUnNG6sMpAxQwDDgqa4WOwk4UcjH+kduQBAyeza
G0RxB5RTbEpWLmjrpSC2nAUciwYLbVHkXCiAggC0kDIDimnxoOXdFc1FxrLhcY2B
dJB7jHafkUhW962ddmyjE5Mon0Q91ISvz5xL4NAg32+OKGdRSZt8zyfzgug9XLUD
9nv9u0Wdk/G49TfEzYe3ya2loWcChjb9ekbZ1tDs9cGXGBJAobHLsx/Y2iaoJRkN
JE50sjcG+jmbnsWIEE+eD48fulUP5XPP3wLXPM2rGTWqyakyvNUuKBYLFKwegabB
jaXK362/uTy+MgdC7yR1jiaFn87d0pqC8h6/PAMTXws3cRnNU8zkLz/Bp7P9GlM3
dudlk3c20ir4mAjhJKdoKa0EJpD6C7o7NPvDZf0KvSMChQ9KUj12/i1N4RTVieWk
FW/ByFLyZWqEb/7n482WukgvJ79JEuwJTPEQIZ3db74OSG9w/HDOBaTmMz+DSE7b
q6TqI/5dP/DRi94qdFL+uLO7HkdRxmR+u0QTAncm2AK6FTLJqo/rDf0vuNVdudwV
EDYVXOqNi7T4edYBpNtxQqUCxBCm0tp515+05xHXnpbXtgqslGkO90loazWyi49K
PvrYsSeJKVBY7cC6TJeZ92l80BUCUQLmbcQsTzVSl9jPMX48CZImqiFVfA6lCG/c
0tcRdxyR13OK+6FiYnb1eSrVXKTVMcWEiQ1k6sQ/oa9XkI5byTdJLfQi26XKFFQm
VvI+OCYpld+LxWH+JUqKc1zhrr/GA440JOOsWbe7a9kVs7muld2Bc2gOjjA4YKZa
8TDDSxxAqCG44XTV4i6m2/jN3vhjTcDS1/RjzBQLX6zTOVc8wjg5GFY9IQ1zjIBe
SnjYYBecIm89h7drhvnffMVrpdeWkbionl8o3XYUfZtFulobgpAan+zB4CT54IHE
iSD3MrccLbygFGVAb3rVh0dXERdqYvcWMMtj+YjqlipT/gl1DQgybjKNm2O5gdXb
lVP7+ao4d45b7NceXby4aIQZkUC6xX/bzpZwCoV0W1xwj8QlyQ0w+Wah8i/e4af3
YcjxxgluVrWa4iMQr4UT/Iyozgo3HZyzlM/gPN7/fzv8wXRXDmCw1CUtzlU0UcCf
l7jJoiYWSBrmMi2PH2tqzgOPu5yrZKSDdVONT+rghWdRDOs2ct+rFZwqsMMyP70/
LdnNrj7sdDt9DokP2M+uvHsIl5rfADZQf7Rilnrms6MoihjjmRfbpQvDHF8CDV8E
+bZ4S9IL2OHcKsHG66zghMU7PLmnzCsJqLniUqsZctKaVNS5O6GJ8vEYXE11Gna7
z5u+RW4/3/0AA3BVke7Nt9Qfw+P+T1XaCBko+eVhIgRJvd+6wCVxE3f2WZwcv08E
6LsZvhXOUYrrO2M3Mw3sNYygKJA1iOPCHa/DH/rX9J34wuZNSg4uT/vYaKFGj1cw
ps1jfzd/fxp3ARvvecwkZ80JaZfQItar2ZJoMmu/SconUQiukO7+tsK10Jq/sH/k
jpAC0V9czaMvrcDPP4TpRBMXu55FROWfLjeE6mMsyaABw10N1z/pAViM4rzhS5Zm
BHpc1HglriOqXl4LmS8CsOoMojxXO8b06OaoqC1OumOXf0xM8defw+ps3RYq+1Y/
gGQPC+WiVCFfZfn+gm+7vjDiNrSwr1JJq4fRlq2RlF/IwMLhiLBiKXC7TsWKzURL
Ci+I2YhIMDRCmEVNLFaDgsZFSRnLxTkCblDJGTBer2qiL7CNZ2vmvKxEsAA6ilIB
n9zeIQI+g4kLnP1oStYLGTDeFwH72gcLdP/KAUwTvMfjlvLqSdV0cgBv1VWjLt4o
7hn95DqRd1YFAsgx7Fep1TphXFKiCEXn2lmq61rrwBIpkKvQMNv62pIC10U9TN5/
fk5wQU+mhW5P58Hzg5zdrEzMufumpNc+0h3Qr1TjLDOyaavE0uICYaVD5uHhE98l
7O4bw7x3FaePJlBqaCg/3uD1MuEeiqWlfiv9hV58MKBLpXhvejk/myVMCcYj4Mdv
hoiT+BEjQu3h2DfsEl50mEQg2Dzv+EOcSJg3TFwNnMm3o+8cIzMpLOzbx7jXuzI+
XP/JTvFLBe1Qmsfoyjhzu55j9NstE9u///CAXpmhpIO/g+esLG24E/SIQ5O26tcf
XtVQX2mrGyglBgIGk/FTZTIWsWCQAV17J0VLBcE/dwkQ6709tTcPr82RfDG6GWE5
zFyQ+NukwTRs7blsQ4+uZF2hH+RZ/cGgEVopepHdqU3N7WGK0a0LNfLBofVnE+CM
d66qjrtbHcetKXRUAqtdZCT8p0LHu5lATPx6WHyHbCR6jdyXUj595Vt8Rdq5D+i8
PTNm0c899QnVihFvGptKftn8Ej2EjwcHAOEjqqe6mQV2fI+uJh95lyycNxvxauLi
3EDkg+egML5lKlJ5MHiM6wyWWUBsTovKZyx5pTq+zwL7inIlgGcAcJ4WBsz+xfBe
QBYoPYl/ijMH4UbIgVLLDam25RXuNxo9PEjlgSUV4Lp1/AxmPsW8ARfX9mjXfWiC
f7ju+zJtDUQtLXeUhcae3zJEb/s/rdDhI8u4cK8oqZs1ZLXPp/7SRDXGYYY9HCii
iyO8kOWSUGivnf5wsrxG2EAlMYDYW3W8c4MQUa4bSLS6c3nu7pUM8omBuDU6AC6M
Yk39E7NoPzUhEbsNNOH8cBGfdcFYchj3qz52f4TI3flGDMvEqYVs+M9gMSkEdiVb
mC177dl9/t/nT3JU2rBmWMnqIIR8xaawKxgwGiiFRMtuEaKE/moyFoB6YpfmTdZB
BXSRkNG9nHHllvQzhBYXaaQUL7vARLopTPpI5AJriDi24bU7SUzVzNWvGmItDNwg
hPx2wQ+/EWOpgvcl1PWt9C82DO/IyyiQ1jcJxioqAoCqp4nBolewjVaE71cwFMbh
L2UCxn8nfwvSKUYtob79fLlgU22s84y43kezOdRxguI0uRDbO/dJzA2GcXCokNPO
pZJw0g+olVozV92u/z6l22GC2IrukhHKF04IJMBTJSMyo8r736lMZvx1WhGBsQMo
es7i/X7BqNkIt0ba6h9QE9nbp/1YPdhf2XbBmRtaVAJnOg+yoN4N5e+q8nOMQhdy
CJJT1Km80lf7RsuVQbmcP7HXrYjlGHndayQQhNfuyj3u5D7V4uxINPgwh1MDpPyy
lC16ETjwJIHJi9dAWibbSA1HanoxcnZBPGZzS6JVNrr/u/zh676mPwAoZT5pYbBQ
4bxRvRuCrZEzcTUIVqIT9FKiCmMpfHU2iEHXGOxxCijtF5JR5uY7kAoXqEj+Infl
BENl4gwqb2t7Ox2coqoNSqGsQYtPkqujD48KoU9g+OdLSODnhUvYWvh9deDUfp6O
s/eCv7454KETjW3MXDhVrv1ROJkTGbhmtUrtjf7gl6hbHl/6ev8bCNQey2u/rLwM
CBAOTgBrIP477NZY15d5V38YDkCLlByazDh63qXZGb6eYaBZUjXox43UP06rKup/
urjxdEsW8fAeZbXhpRtI8hzoxHi5UApQowNZb4JIovGvWIdk8p6YomRuWDYsGJrS
IbieeUaHwzSINKivqUdcoVDUrlmTUdEAQI+zsOpV2VqrtjqPlvDjxwDDkRm6hetE
RLIoHUgdVCso4vWKFu7lWgw23RHVU36/U1vfSywIxFBn6KNneau/RPXO5DiRsilw
s6RkvPBKT3WXPTASW6z7m/mNQSiphsqlVxl+MGz5Lh64p2cK3LVceZFklcHxbbZF
cFEBGZjXQqzlBxdwwlTa+lSEnRxYy1yjUrxplL92u7DY9lzOGoDIr3auIaqPnY31
O22vxOYXF8IXtQ3kKTca/bJmcIdYLxM/vilV8WmVzT/IAKJ3u4svk/N5cccUgezR
VJ4Z4PvWNJnzEsVuVIefoiN76a/FfS0vG28wIpGkZ8ExMdO+NlyUT10rjHB2WmFe
AitJwB0CGIfU6VS8pfevz4tRMfVNgkYNSbp1IgHE/qk/w/jZ6oRJF0uj+COY3bp/
lCyzphNhmBMFPXGBA6YN8OPMHs5gbdOQl5b+esO9iDWk+4wL0ec7VbJ+MP23nE4u
cEn26Jsp5mos4P0et/lHLSnvtiX/Ldn7GfI/Es0CVz04cik4UgxP4ITu27qEAhv8
DwwZrqCjfGU7aibn6n8RZarmSUTQscH25uLWsejecz7vd3kWT+OswZdtkIzUgiXE
9aI4PMibngMxewNeXNW1ZhUXQSy/kooT47cX2ilk30obOPB79yV5cnuF1Y6RsjDP
ap8tN+8R9GkzOIkHJ8ZfoW2ixSFRH3DSNWAIuNWH+gIXg26r2mLu9y9hsX8mcuck
Uz+aFdk3mRBFZVFROCu0wWe0x+Ct1S//XI+C9WBAMZVc6UTcGmF8EO0cHA6bNZYf
JItxL0u/yzBkXDYolrZHKLWf638e/d0UyqqtfYhtdWX8S1gHsaNXjMpKh4z3YbPK
BnCtDSMN7cscfyv7INomH+u6E4pnSitOjAtwTTPQDer0TrdgZxJo+eLlY3j7DASd
HTTj+CHiKhQf9KiOIMlmZGwlDG8iRCXhelP7cqrFasg2b/Veb8jDe9YlLGbuhEVQ
Bh9bHOQAe1QpuhNQeVjuM8nWHvvrjm78+AD+Lfv7WQffS0LqvTlZa4IZhD+I+87G
LB29eo8M2suvm26iPIyOTg6ZNOmu5OfsloF+J2pQjXiiinpYiZFl9xObvsepzQpD
M7HvVmedzWImNmAX/mcjgpmBSDaqut4BNOZOntP+RywJl78IgexHwe2hgQq0Gb/v
wUjg8KAzXrCdWgmrLyEpRaD5EEbkS26JUQ5BqrRTMeElEvefsS4D2L4MLVK1bq1E
+Iae3aZBpyHn5hLAmBHj4ULP8A2+c5TOhfsN2FE9ZMKokhcq7Mr3g+H8TEtDV0DN
TGo9wxgZdfCu6gCuxaMrG+Q7gP5NZVAjkRB3cazHTzoyuqgncb1TJ2M4mo1HU0AS
rfT8lBrjkJDDYY7KDbmHmEYdCBMq3l/qt/MZJngoN/6l2tNaTnl97JoA3bxhMNyb
hC/7tpFza+FSaq3UUjSfE2z2v/2taq6V6mB8ew6luwn3vkiYqUVRtOd+C/EP05TK
JB/PUxWtDUO6rKqW1ooqPe1XTQ3PEjPTUvQpRbhYjR6z9mX96sGFHAt3h1azf85n
1erMZK5A3vp8VVD7Bsb0O97pA5JcsHXvS11rCsYXWU3Qk3Hs1/KfAtjGgAkalL7v
fINEuMgyFp6WSuaAktAhQNha7IA4yE/kmtMRqY6KF8sBscAClZtxF4WZ38sBlrjl
2Uq6o1S5eeOMYWYsrLgMqWgaSqFJ7jeEPwquzs+VKvgvQ4pRl9dQsYihxZJnICwx
Csale2nIP1LCAraZDVkmZGtXJynqTuewGPiDDmY02Hwt+wwjnyXJyWw5f0DZR1yb
2aBboyfILWN2SxC2iT8thQKsvEPOMr72JqyI+UD5n6EvVhIKXb8W+8PaVw/Pr0og
0SOU+xPtFvxuIDqho+BvR0/kanK+/7wLIwRq4uVXFA6B1QRzrQoRMMkclWv7BQ+Q
MZCw04dpFbn7RkvIWfME42DRKqyrvmasT2c+JdJKriEuOczZhyP2gbsMQ1xcOn+t
naNp/T20KNrrNQyuAC8vyl9VA0F/tr9LuKHk1eyRsrkW6lxkz3ZJHVWsQ0yMbjkc
tJBw675j67eI6aZCq4u60XgHK+cdlGkOlfsPDfujb59D+Azq4nQScxczBbCbLQN+
v4d2xeSIISClEhmT2DG3G4YOizBUzJmdCKPLGgSo9Q/oL0DmhH+nR9H2F1Y0C9Y+
EXK09j6USeKKZiY0BJmUCUeLOGq+IL7jINOqr1UbW5+ye7gchWFjIDCjeAgUlPJA
av5hnfTojI+Q4FCDLcz6Wvbdqt+M0D7EBQI7xgph/dMrHp+ZoJTXcspKBSm0qrGP
6kIQzgW8PgtGFjjOkcXUbHiLPvOo8ALbMXlcTPR3iVUyh3aNTv8j1czJyJcBmRY/
sooXTmeHUdUEudBTkLoFXFXGLmVxfI076e5qMAfCVbVn2h/NXmn121u5QdWm5mUu
eJoYdr0vSVuIJhnZlH2sldln/nsw8fF5SRTQ/V7hMq5qonaSlgn0D+fcuSBB1iIC
ZzcHi+T6aDmCFo7w7PxBrCiTzWu0hpG1YWCyYPAQkqkD/cVMYBGtQ2HfGbNmyrY8
dF2mMihGGJvaKOmpUU9v/napMghcuGqaFnNORcaz4AHHohc/RMKFJDfaki8q8uZf
JXZku/9rxHhdBbAN/qzDwYxwNLhWtH1TzaxcaaK+TrEn+cd8xl7sDG7b3xdjS873
D8ZGGkVWUfwKGvitVtDPYBpjh8o5JsSVH0MB26Y0BZPw6iDQZHEtZuAs5TA+EeMi
zNd15tqXoF5FOccK9W4UQIILMQDqEteHEMK19KP2Q5jWfRYDFYZTh/jt8sT6pzJp
h0FhIV0kzQP3u4cIdlJYZJYvxU3pOzwAm0Lpr9BFRi2qX5S2pIJCyCNPn7677a6N
xtfbged7VnXigzl6P3Bkf8NTi1A4S9OAaE2DA5F82w4A0RLwq4PLxbM9aiPBrgpf
a87AkHTaOWc98D+ZRR0/OaRoaTqNVczIAZkhPguT6UbxKGpWsLsKrAGyP09zUcax
+4BOzJsjwXaLOZ//So5dWSpz/yTQiNtcE4F4F3su4oczYmpJr2yTIddDdB5FOVcP
ih1VWOWmf5FHdWt8B/gGnO6Ci7McUBBFSRyY6dOcJji56KLBDn0/f9eVIYkxxio2
VaHXx21K0fpoRkmaDlEjXdICluvmWks0tUwNZr1A3z3zIsW9DGKZMNj1pcmR5aK0
aKvDujio6h3H8i5M4ts7/gwb7HGvJLWwlvuFl6z1LOOInVvW1213taiqtwexuG5v
1BtYr2J3PuX4KgTRjarQZqeiVWbHhjGoJ0m7CqGjB6w1Yk089Rzsa7PgV/zvP6+S
tpup4J9IhyqfCBdLyk9T4o1N8aL8Rh0Dh3kJHT8PsAs+/+qi1jWjf8zmqoeu59rj
blSiXqQmggePWZdqw3Mk1f2NjNGRiGNP8bIoRtoEslmdH+ae65VzsRg36Ud6JwZz
/ORquNPH2VFMIGgKMBbSwcMj3fdt69db1xDz+SLEUAu/j8KK/5gRdjXn5v0lh3Vg
PFfjnu/3wEgHZzLoTgLF1TON+HmrFMYq9wjVRTUK4yMarmvBM3THIQLNyAbf6TeI
z5Sd4r0O21gf+R9xyJoMhgrmZ0kQIbf011h/E3zwsNOyI5n2jAhlrHYf1Dq7pO+Y
DCCZbFSISKY6JBwgZFubCOC17mOMioVL4dDVOCDd3oIesQNfqpirlTOUVVpx2go8
EIwmopbBXd/SNvtnjQKu+RWY1nCE3ltc18zOqOWBQZsMSfkAAvFZ2lXcrmkhm4Mh
akp/4TmZlGfYrMDEJ6Kf1ITHP5ccZljQVWERtueQYdn40QtLw+Ap45vdpUXxFPwo
pV124LYAnxaRDLSv4lcISZis7DYYD3H3ZZxkMHxDWbYaxG8Xma51caNTerVtqtFp
PbV+wFt4EGHSuHuh9GwD8Y2ud1X9P98Ro0aBWmsI1wKFfrc27y5xSmYGokBpDEwB
XdJNJR/6e7nUhCD3udFy9XyVTcF7xhVmfBkZrMNwiA/Ve4Re2FDk+LkBx87+jLxM
edoUKM7HwxGnHkmYa4jMeMzwnnPGLSjmyCEc77zKspPnUNteB/RhrrFyYyD8dh7J
hRzwvNdg3a0bI7MuQabDvEH66JTSeWw518tds1T1mJAGMB+mh5U/zU+1WrNSTF6I
0TuR2FWTj8Rxe5seYVbWYbGYh503UStBBnHwQZdWTB8Ln5wIPYI5rfy848qHElcm
CAptNrJcKAQ2nh8sYNmD2I4ro/WV6awul/yy2lNdWllLeUjfU3n1CckQs9vYLygE
jHa54SYGjF3GFj5trQQ7SwQGdcs47H55wQWzJ0EthCq8Ctf0tm2fgATpgb8scW9p
5Ycjc5UiCfZxv4pOWYfepb517yl0n2z5+NW8E/Nxl2ZXAJjN/SLtvl+R5JwFJeF1
7ZeEKLyh+e2pXmJtvep+v2y5IRLO3iIrj3HTvbIXajLs2X3d3s+puKBUTmaLwVc3
W2g7mzM9eV4rPlq8wD4VquR2banFkg/cEq8ymaVvsqJ242IaBiEMwHR/C5xNUfgD
VMMr4PsOVrE2S0RuL0sUFKn4VyZ+9cPUUQyAo0As9GeLtXhoW/2KFoeFPji1Zqj0
ynYPPCFW+3AuJY3RBoiAJpxPgCwzKteIdZ/mTxkT3Ecs4D/XHa2qYMaaq0pQV0H9
rlOAcYN4PGvnsGmKWOwem1HYDboHegWMtLSYP57o29YMQnerM/tt6mCcZTzAGll5
4rRvFJzjWg8ytSVxl549HWhr2dCGlLufdPGLx0/Hhr00qsYEnCTltWRXplEL1gdr
9n4un817U5SC9l0tEH5PgO6/OSz/amp+PKKoIFMFQrNGz1jwP5v4AJs0CID5C0WL
9dU2M9XBcHfLDdkrRa7ttcvef1G21teWlW+IaQj6sSMB1kflndJ62ML6BK7dZ63Z
Py0n6vKEGk3Fkwb/7ZsbCSEbDgwoVzCkwbt7cPOxWcr/84r7nlNEP2nsnW6D9pev
ZJNlWjIvKcLz7hSHYnbYr8oc9uB3IETzgiHGAtX4GoxF53Xr2rV2MZIADR7uKikv
D3xRbylRYOarUof68S007fikOpQ/JyXpw38v7kAhO0l8OHolfHzGpJdKxVCntjsZ
hM59mXNqVT+PNySs3TgJWwaEuSlf5Q5tE2TaFZwGfPdEjDW0zyz8xYmJAe9d9RKa
mVdNQeem2Nsoa2vdC+vVZmI1aB9Xp+c2nmETMYJ/tkBtw/AjQqU5BqgPwgHehB2L
RgfEv35BGA7E7aLnbTwHThqTlbRTRuTFE+pKocQDG9T0cv3ydLTti1K4sy+goM2c
Uqy6tR/kiDJl9qXzPrPF9lwL7I8Gd0RQlG3c9PteELaYaGQmRVW+0v6phowgjEW2
u7T1rUeI+APWvU/SyCFCWJqm34teXvwWlqejY6q2RLuA2lkjJuTTQrSJycEu6aLo
EdpSNE0x1igbF3EcHfxiiqu+NFM15AUGDnYG9C4WhNlcVeAbRuCHnozvdrP3ldLJ
uWc949WZOzy9ut+NdH2ZQ8krnzpDxe1XhQXajwsWr1+PTbXWUKOttT2IVwcz1GGH
l13Z3XvKczURPVjSQJQZCbCf/UZ7mEjScholwNtKbAPC0ydyGqB/mNQ6PySzClIq
B0/NctHpVqqJPBXTIXQHrcWocgnIIEdSo8FA8v/oHC2JdY3ba25gUt1Z8PDVsOXT
uaxipWK5q6F3T35OdBYBT5Fls45loefnaXQXDhrH7VygIexqWNONJosduFM9JcRv
pI92mBk9Q1K8wNr7/cjnJ8P4cswgBFE1zBagARVxpvUq/UGfdW8VDnz5pmrg3IZ2
+fh98i6zR8XG4/xHjF2tLUuXue6Wp8TG7oMk+jkUTT6dEw+6U1d9R/U284lR8EQd
kgACPU02N3obb/e8OZezKfYKO04D3h/2VcNdIv1UWmHSlGKUpbw5KIWBZrQTnhha
+TwNlyLl90MGGL8JBzyzkEdShZHuFFfGORw6cCQ674DIA5+4x0xVcc6DIVr4j2iN
LJbULQd6wVCThdoIZ74mCiTtu4GHwA+3rahdMUaD1zfw1Ox9lUWdCESK8DyNo9jl
R+HyzaMaaFH9I8D6IOlPGlA5g38ifN3L642ctsb0HsxhcMeCJ7Lsre4Dd+sCmfpk
6kd5Mq3izZb0HwmdsktgDSplnFTvqYXl47xLaHwVYk544El8um9NywMrgXqr0Rv5
TRljhxbo2nCK8+irKy4O4sFSfh6Pkb7arrHZf3cN1o5wllHnbpPTM+UqHzNCA8Iy
7YJ6Bzh9TnLzg7vBHk7nA0Ro5JvXfGaB7Vgg6v00HubpyN5XotvHjpMx0jN8hd/4
UfTJaj/s3ElyWryxmMBcERNtozRKFz90RfHZK9jLL+EUIXbOtJq0j8UK4N3q3ixA
xWLMcMChDZjRxUOKV1dO0rVjJpPJpMTAhkox7jyw9YS1/HAxyBYGWd+Zh2Y300rr
aT+f2kfWlRCavEW++sUjmZj8IYNB/xAcBrhZ6sgjjGqOqa5xWh2GAfu8TkLuHbY6
e6hXBWTurJdO8YxheC3l/9k4SQsNBJl1i57+bJYgsh5vL789ujVOpSgSHItn3cdI
G3BDEdvACdEu5yh0N0g4zBZWnrbIRKHBtvLuZjG4nJHRCXX9rFiC+dKfmnf2yBHh
wktOmT0WWVReyvrdTnAgGqtqYqS403waCas2X0VS3FWtowp0zRTFcIaWe5F7UIT0
l4NhaDLoGZQhMVu7LuQ7yWH+9StVbJNBRxHXsZrKXlJ+JQ/uql4UQb/clt2UPeoX
87ea380v8TE3Y+psDo394LSS7mP/VnUWN4h9cIlmffxMggARc875UQYdRFZGEioQ
gY11FusA5pemLNqj4uD5Z7Nim/2+iCMwi12NRdNe9BHUQPsLYPDay1APTZhZ7c3D
z+niZrQdmicsS/UKPSjHf+FVb7zCOYIOp/Qho8hzc4+r4NX3tCPn/whdRfhM/s5v
pXXjoEbsw8fwHfrVDinSGqwXQggPuDQKpVH0DIs59Cc1vr0+Wzz88yS4CItANt8j
oEsD5tb+BdYLADpMpo9l9p8J0GwRH9Hhh3Ay/GkPoSjdGYSRRaGlTt5wj5v3kh+v
npIXbdiD6M2Sd5AUt6yoNK05XXYPWOMlr6851I+9lP2o82RJluLILGXYgpnkFaga
ZHxydg3B8N6S1pwmEP5rYn7Olh9+RRjhj1KcN6dxWhObeEj4iPrWSah3F4YZz1ah
tcvBnRK+cxtd19atVbO427lOYXPa7f60M9CEVeqNyzF8dKtW7NrSnGG/8MxPS1km
jHpL1SizdWpglqxpX8NukfqhVheoWrQCu6isLBq917JMApMZb60ZXsW81xuLo0Rh
DWxLl8GrGyqOQWOdgnNlmX9U9Gro48nq9geSv1cf6jGyiTdpA2hQFbbU5b8lQdYY
P5J0EoX/ovb+OLWgkXeypNvp88PIJxUiutGoOjWOv8SGg3YIEe6/ZDBMfiOHVF3r
aqwhDyAJPOon/7XVZoedD0jN4pInpTu203HXxQlA8ej67RDaytZfc2LpkmJkkXnv
vbycuHyoth2/lQHeUh8ZeYH0K11hEVyvWSJU4atAi7nO2+hDObxXNOKkM+2pm+Br
qUsaWQzAe0YxlfZPZyJ9jRUyTYd496cFWCZqvdw2mSDYp1Pqnc0367Tw+9+Qlnrb
7yHC58jj+ItyWi4koGF0RpGAnfHyUaS8WhGzBtq3ESWnNqpNv4ioLzusKUqkQQap
dINuqN0I7gNy4ZCCcyUyrZJPkg0bkoFn+rZm7A8otcyvbjGmAB+/86rmG8t7yXRh
RIzm0zKkCKVXSSB7nvxaXqsokdOugGMAJsuv9oynIjJA3pjZ+2QcwLCxAqH/XLQx
Z1y963jwM/Vg4yJPqBkEFNoBR6GIGXJ4yi57DnwoyjXEwm1b40ZKIxUQ3Ru24ulW
7Wa753tku89j72gllNwxkgJJNj/0xO86Zndko+y3cCbnpeNakAj/HWp+WuvDTfqo
sTdud4aczTPZheBHdOfcW8he5zjFqzjZZqk69gctK/33npx9TAlETzt65k/Soipb
W0A06XgZJjBwDkxQSMC0nSDDtphFDlKwybgmV66F3XM+Azz5Kq3xM4pg+YPblXdS
nF+cjBj4Sswt/1Ocsk0rzhrkaCOuS7kGnPL6zCfzvMSdvMkHIpGX8UDVx4CgCS2W
mabBgLTFuoCfaM/ilC0A8EfgZ8kxE/px49h+5N0mDOMvt21EcenbPeXMA820AZHi
v2yQbSXid1DU3/SqCG6OhKeu0wq6t2hF8ff/YHkipvaZBErlTPgy23H5rwv7GJut
O4/eKdQoJTiAiiGv7um03Be/LW0oZD3VoJqM8VlRo0xoZmFC0rODjQxAqNl0I/dO
I9IVKR3p6BfqeQ4tNdxDsf8hhbkNHXZPylhkauq0dPr8HeBJ+HN82a4SS7RJkmzA
79lhqgRbuTw75uL/y36Tv/E6duI/MDAP877vgbxCIC0yfCqlsBfCjuJJxFe/LYFS
fS20xfaBf6io0XaAzgBzVqIHgX2pY90JS1cBBN6dJ+bqF+Y2vl3jh8m+WhgWr+6L
luaecEqiIpOAxxmBR+Vewp7c5Km32/IPKHFsZEkKGNuEHSkWwGdZSAzKX/ZMMos3
kcj8DfCNZW0f1k18hwjKtk3Pg2UvBOV+F4DjN9EYNni7lJnXL6dzpm4mT+LRC9Lb
c9U5oZGgAGYtE2IYutMMWTYth9G/L99mFMO47BkM71zkmUb8fnjKgsECgCW0R4Jv
k9n/yJY2zbY3udPhP4/3EVs9GYo9RNbo6rd+sW/nKLZaqIQH0giGD14esIX6/MCL
oPicPxe0I7AQpvsWQNAHowp456u3xAWkOskYRLUzniQqlVH7e9PzvZenVGb2f0Eg
ULnGOkWLpBqUJnUir24q0gLKl38rN7GAj4Ng0f9BcNbcxStzSZKTYmlqP9g9jUNc
7aTFUNDBuVSCialJpSjLHH47mKx2dx5WSOWmLWvinrObu6oyFvbI0n6+YuAf86dy
uUE8D9nO4wKIpfzwNolsHSFJI4N9JUJmMwqnKyz34O9y8ezJihtkPc2Kp1GTuP3Q
KxwHIvqQgwzKDoQ1/AAyfxpzgdw3g2SouFZd3nJE7AuT/rWJmBmmL7chWl8ybnMq
rNDPSyJ/Q+aO7rs0yY8FWNZUklK8w5rFtAAaMVYCc5BJekCU5U2S+v4O6Q/2oPGp
Kg1pfhgkyfhgy3UdVP+oBhzdhy3SglRkcATfp02QyfBXSuXq7/fy0d0GBZJVPuCo
DtAHdwKsv2tNOmD03XXuxzRrOIl4E481YjKNYbv077DWlkoZYNmRS6ZvBqyHkQTA
dMftrvFk3BJWrJVKLmOEG9OZ2LajO0VKrWy1GGWVxg/g98soWH/u1HnEXh/GAGe6
E73vh0wKEFK446OlcYPXYxOAa8wB5HKU0W2OobLf5hdTf977eiFjuu6dAPmQVj8j
NFay3DLg8u4Oy8vBy/SZ8mhbufzRTce1s+dJwFZkWCwOhK0lcHT6bUSuoB5BLa7T
tyRVA8XqXIxRhJcPwE5i6qWgX8xjx+7w+wY3CZx6Y4HTnBnlZU2RVGJkttGpEl2E
0qhy1CEBTg920BbpwTdefQXBjyFNeY99k8XAIZByM41X4qR9zmthlWMr3salCWOv
VyHzYwLpZqxXgVZifGxKSRLKyahLxIAjGsEVYM5DdNsswG+kkhYv1DIzAP/+WoAM
z1oO3Kf6DtPUnWUyAEQmm1UYxk19gtGPB+Haaf/zHWrBxDJwbJImjpwbtDj6CAsv
fazU198u4fx1Qq3Xb+MZCP1q0mkzGSgjOqU+OOjGaj2ugSldm2QLKHQdZkQUmNlQ
9U0NiMApmziNz8GeS+rwBksnIRf6ds5WrCJFZUMbG4050Zz+U5kQF1j5AzXIwTec
6O9/edEAf7DzlRWRC7VXCI0/jZusAMu2VP5Pqtrrl9Il7QJqvMKn+GQP2RCnCaxU
f6bougR4jiGdz1bt1rWty2dR87Yi9nL50FmsgzasWlpY9VLW4PrEuXWG9qxV4w0H
McZmTPY8N/kw2yq5urfi91r9mdLsn7ucmJU1z563K1kWQnyn1RD40FrZFqOHbobD
Kqu1rMnNjZ1X/Dyum6+haVSKyYNH9hgXNSVEE0g6gqJMLcyWFGsdyx/S+gn6E8f8
D2UnJU9lzsCkMCj70GethHhERE8pJmHOre/wmGixaeLaqCNVbTz+HFyhqRRk3FsF
6w/CgMB9k6Zrg5+pKZ7Q1+ijFhALo9xg7gh60uDr4qU9/m236O2G9G0qFDCFymGi
xNt10Bxe77yiZm14ko/8ZllUKl4cbzs/74G0IzZ2kd5BfMUJvj0+o4FrKkXTj6KS
4bZ7T8yu0bFB2iI7pkgNeFYrcXAIhEtS5BjBS27rBHiMPmDdXzFhH7rdjtDmehfo
aQG39Wujj0CsbtlL7NQi72Zyp5Oz77z/yzJU3dBdElc8tRjK7AOP6F4cN/FKjezk
BRwt35J/y6plfQENWWvgBA7JJAf8jr86jiZmcmv2GzjaJ8wpU/iVtH4I+qGfYvMt
tsof6f6MN12MyYWZxD2JDM1bXSLXkQAaSdqzgC5p0jYLGe03CMAsp24qxz6r2nCT
YVKd1Inqa2C7pgR3Vyo/lRwP7A5VESBajU5Dwg6poOLonbsgFFMGDQjQyfipia6V
jYprHyUs8yqfc0IMn0R2nZc/LjBQ/4TOXfhOK8x8cUM70KRVw+iB7gsN/h2fYAYt
FmFFe2/+B0sepX0pg4gPOh0n7rdw4hPzQrC6wqJxY2QmFKriNrujhiOf8ZQyjKjR
W8iDVS9n2dD0NH8YJGerSAU41IvCr9GZMzBOlg+S/ndfuhOp8epnA2i8MA8hBGT2
Tl6nvNabNH6y06GU0SoagM44sJe2X5FgkWVC3od3wmKjAYand5maGqayB75W2bl6
AqPxYuG56CmPxat5X9YtCpL5WwO4Otb0tq7m+Mn9ksq0l7rf5llkirFaToH6/N+s
IbB02f+qf4QCjyHhDb8PD+UXBacIuIk4fdY9y3F/92W/fz45am4xTrwyCrV6IJU5
RpXL/uN7xDcLTwdxioHZae0AraeR4LxlJ7YDtAoh7+GCtWQzLE9admRnkhnzkBHf
fH4wEIUkTmbA0a6b6Jc9tqi2N0dzTR8+nduto/BQdCSvvBVawAAu+R4LbfEHPIH9
XyMdg/gEX5AcDRPJkyySdbhsVEbOfFGJanmHDbsN76IBRFz78hhgZmv2jLOrmnb2
vY0Tgez1D/36hSNiXMUwJFg+V5lRA0nY1WhZLsjuZ4eOoAPqZF8be8mfC4jmvf8L
Utwet+1qPLXh3v4iajiRGOowi1wKFGogrIZsglDnAHZLPlpufRYo+JCa0zzOL46m
uG+xaAcrAjE8lRvEz0JPPcrZ7W/fyjHUyFim+w3nF+KvPl0TEy4YnjkhN4vUC2vo
gke+Z4EhnGUm/abmH7aoufFqqXCg7mYZDWrgePYuSm2jBN8yCFTCBZcb9hvZ6qbl
UpaLwAoHPaRgTvIKjyLi8wZQXO/H7HYQbfheqJ+Hw7xzQFkXPmFErGWMl++4+HC8
r4QR0mcJ4tjdBJ9I0SDvLnYSHQYmPMssGBcviY1yPO/4nuYzDJeZ+WWXeBdBez3f
dMm02p0/+vhELx6rDezYnyb/J38kFCPfqg1MqSPM7UxlYnETP4dqerg1voC22AtB
3C8o2cVDFqCl0TxGFRJeVluknvSfoIuZkLj0e4Pm9fM4OyQyFFSlkYv1AmtYlnwq
/JYGKEWgstPXR0pbQq6NnMc++RckkKeAEJ8JU+Xe6WYJH1+r2Mcd+HDbN9CWoh2n
CHwpJT971Gm0xjjgG6UPx+NFpGGbu6yleAtCdhJKStdceJb+gvHKtwoBPTfGPEaJ
ITF05mc9wkBX60AfwFN+8dEDcv0z8uuMcC6BLyUloMsAP8gTHSqMJPLxP7nNquQD
0BRAQhsCYYzGr3ltBKOalRzcvpWVMQ19kbqLUuI9QsBHUWeVgeA1EikSHiuNkiQZ
wcCw3njCcVCV9gcM+PF7nCCFUQwVQ/ErOFqJMAze4+5WGPmfg+Ch1QmcS/HzY7wb
iWm+/iV75PamFBSwLyDJ7tS43u5xbIAk9B0QituoJJbHeXoRm9snCcxZ6ZqJmcR0
iQAGzBLVtZJyKSl1igQCnpbXDHqBy/MvNSbH/qQbALYKeSRKJs/BHRxppdKtYceY
M1mOKu2ipGG3xxjb0iOYuVf0QeV4m8CXnMD39bC6NHBZRw0NY+FypZcDRA+TLVb5
xfK0c/Py1q0lSi83dj7C0PTsRRvwSBY4tq1xmPE81L2tJA3cjehn0A+l9xRxsGmk
hIZIvrkyM7eUE1bWqf7sn8RT2Hlhha/lbKNFV6j8gJMBDZXi1Mgi6zP33Evwbhc3
RZWATwOTI1VVxVSvQ7e8mm9hC/2MDENO66i6lXwgdNJdKzkDUrqFV93kdn8OG+lA
mKcpH+WZGl8pGZtS8ae4wxiObSLDIH5TYuTAFdncgViAG0rdQYSQgTP1Ehonc87w
oIN8p3+QDjA0nWjOyACQySozgxZ36LiL2JYFkKWYw4mO5nJyJ3EWWMm+0+yuolyh
SNz7Lkuz3aw0UTwQ7IHMHPtbYaPk40+rldGnsgtthKlWeyJCF9eHSnyuiCReOk0D
wQIjp04meXeeIjwdonJaHzV5QovVnkDOAVKN4G7e6zn/ZIW9fYM8yZxr6GnacjZc
uoZE7KHYK4uhtNQB25zmgEGhddvOnuk1Ra7mvNO7cEiiqQgLJKcPUzeQx0FhBETV
C6hsrPlNFE/fh3uYMXKv3zWfaM60cfn6LNGkix3Rp78ct7vQoELanoPu1uVxkcGD
s9vuv6eQUNP7RWV+aUMAapZ54sgy7D/SFWpZAmlj2Kk2Lc0nuHd/mxq8Uh9IIoH5
XuF7HIR0MFUPtH/YhJOHLeTDDrpAXoHv3Ecfo40kbMoWvKAGfaydcHpm+psJxqeH
B3c4IPdPjFE7HON4X69HVxEcE1q4NEjtNvvJnMDdpu/EnCOvVWXSquIcrW1SSzgQ
orH7+FQlrxcLhffoQfcACliwk6+Zp7uB/J9wxO6aadEW0sNW3o0Ac4jAblqDzNv+
k8F4N/OUWLYmItjpK7cYwuky1d4HTUHSDnpgQNTElQALRkeFuJTj1hIZK7a+1ql+
McbfkxO3GdTIvBSSKNBs+9DLgo93hnSJe3RPMJ0U1WtaEp48+WM2p8zUV2PU+a8A
hOW52n8pNXUoF+T+UG5g+KtRIO+WTPm/9H1Uc88CEFdeL+x9CFlOjLYwED2ITy7E
apmQBliSpZ2lpaOklo2693ePqSMh+B5ERepyq33y9uV9+rT24e0sIcySt+aBbL/i
zPj6r+Qi4skUJ9A8JsMp4YIqMXSaLYcsgocIpzAA9QqYdwJ4zcDkfmWs0SUd5yJP
CtuqAW657E33kRpKHSJj0tBDcF1bPDqE4k7xCj64PeXt1uHg2AvkF/nTPbXX0v87
j2xAjUJJfBfIA1soQzadrVOk6Kinuj0KrIwfXMSnkW7CFQf0QY8Gaa5HZEi6ddlW
UjdiyMYp2ZPfl63R+ChVpAMbksBmvhByj5caWsJi/cien/LhwdpMErUnJb5frMVI
tcnUXee4OZNIxLHpQ0/tSWAQuRJqbNiPRT15zTaJw7oQiI7CcckDTZ941Qv/8CfP
P687rTzMI1NPXlK9G+i0OnCKqXsgX6bRfMbgqnrkYQMPDXelwoiMzfjNZmzNGk32
oQhIgxHpQU7CAPeMZaSj/LrzNtT1RRjHQCj9+ULz2KzUVzotgAqEYHz3HlSJyj2M
2avCHVCmUXY4DvcqJ5b+mDTvdUNfEeoSLUMbM/q33yNm4VI29oi4JE/qI/APlhD+
ANzR0yNyko4osAd+eoKYBrQ+YMnVNcG4OVUeTVZYU1K4UXrlWSXHNfXtDgumir/3
HREHBB6oo5EaGMUZRyzzIBXQvPUmpLZRWmbGQ2JwCCIx2RU1tMp8jK7gfTJizquV
ROMKCB+g7G/+TMuBn52GNhnJPnZDC1NVGwkNm2VyUtif1QfMv70rh3KTCSV3drDV
udv2bZLOXwl7xQvkZdW1hMlU623RHOWMn1+xmX3pk0w2PuIIdc9hOu5OHIeZpVay
wNNgXl9nHgRYjsGWB2y0wCQgzntdGUSKTa9QxxvUXrNgh9FtmFdOc7IbpzqnDhME
FUx3VvNrQIbGIsSy8acrHh9ELj4iMULEvC/jv9W8upl6+OVKySoXvoai53HHK3p9
szqo9A+EOaZPB50uAKdNFsO+BzsJ6fB6stn7/zzYUYFk18hzahcuzI8X2voQglIV
LEQvzHvUhR9YvP/cq6A9gwlZLvWIMez6RxYNw4iEC4Hh3LskjecZ5Z/4HHpg5oqv
uClp9b28nVLbCavccmRSxEA4SQ5gId/txQHxOQFybJOA2aIAJLoDlJG/BgMHJKWT
451osoOKS/bYLpwqFGZRgjk3FQkO7X2gM/fYpxLZXenSpeaOjrS9IWKdOLgVYDyK
JzQhpZi/kFj2Dhb3G+c1qRjKkuW2ez5mhqSrUYzYzcizPledqJVU6TYry2vnROYq
oJMRinNsvUv63jX4QMrgAqkf0fGwi18rEXVgsGUxVcyznacCMVYjdLqy71v/bflG
wMny/KNa5xcJxIFLvBEmiU4Q6aKgVrcFK+cC9LwQTnNKrfB0IO8pzJ4cKOtFOpRb
mktKZgb68w1ktdX7oeVom/LKE47f9UEwX0caBM8k6dCsEmCTOuKEXLcja3wROWdN
ifu2p1W86CR7gUwofwWnElggbQZ+SoEcJWqfQ/3LgRXejAxT8do43EZPZd2yTNDA
FgigzigUEaMgbm46uHqc/kfx+mDbvDWJbAwD5BOFFhXbZjKVwRSnZTBN/087PB5M
FbW/Jwhb5tm8jgAFXUnAwR6Lpv+85+AYikSeFjPn4nDNkAWO7L0tMvkQl3AXtC4X
FQeYHTnKJlJStp1Zj4ZY3bVp8y3dzRVqXd17lzjC+yD5mKNwT+FEQ+hhXiCafCuI
9mRXkJim63ksKH7/1o0x8cGyL5sfY0nEz7B6g4k5YgRG/IKOhnAwamb8pU5k8e3N
TsGdq8uyKHNmWTeR1JeTpu07YCfh55TyRod1RbkNRY7fRo14C4Fn6KN/8KE6xmgF
XAQmDiruL4vuz4xBZ0DT8qxuTxzG0jjY7Tj1ZD3igKz/a1oL+oZs8mv/izRKanY7
NuVimxxqqXUngb9N72TGAeei6vRlchWFp+Bw+h4m3vRdTGTylKzjrTPPI3Tfkj1/
LLuHFkO+SufNf5eX82DMmTjFI5CnVe/Yip/k20/2jfcZcPUb+/T+36ROIMN+kSj6
K+ODFyzq8vtPQSRgpXZS/4K1dgafIx9ca8YYIlySSGeSypu4Bvb6L1cfCgf5rwG9
KP2y2amHijOE3nUBAgBtpTU/Q0s8ZsXrRwnPgpOScw6vMWHBEsBOgJgx+jdlF07I
JkZ0Yyx3v3GT7qOLKeci2oVHTluqiv6T1k8vjponz5ks05oWYUQxsatmsfJIBuTU
S79OvGubrnR3XYRYiCK36nGOn18FiF6Jgq8JEkSRP6DWJ2fjkKvQM5y0wl9+8TLz
+t6wmT+aSvh0g5r8eNPqbkI8j0ZcG/tu2AnCCQomb5sAJ3CXYDoSMYX7V/e0DxBW
lU+AxtnZvi7xLYdf/JyQImY3jA6KjsV2668UZKDEI2DgiI2PBAqfaB36+61bmWsi
FH2MalGlGmB3s4f48lPFklaeyjd4tRrfqhzNriRpscCfUr0rGM+MnvjhSXI2Crtx
s0Yz2job1rUqeV9fbKoHIdZnyryQYvCYFykJAMR5FkGU50VYN+KkJY+xl6LXwa35
D6rZfZ1Cs9CsrpORtF/6Mi/xU+qDCkF132j5z+aJt0/gU9HMhWX+C3C5Z+2G6Mqj
aF/t4x1d0TBbGnJJLB34mlnF1yOkD/GZmaaPU28IXUWjwv4zn9hsW8888YUnXY4I
oxePvTgh28+YWbeY8eXyoaSzofv09DRNcjiWtIwMEta0Z3hAO9AtLkZYl1OANLat
V0r9VzD/dYdgEg0i05mhRRNOJvtr0b31U0DvYMw+yQApVdTRJ2dPBUp4zg41wgiE
7J3cVSt56GDgbswM0Rt7WbUb6u+v2su8lS7Bd+efBDXFf+/XeZByb0txXu3iv1L7
N8WxZh8wbvpTGV5lpkqDfsRTbWmwAdD7vHFK/op1HFtrqZZr0CaY+gWiCbYAuR2d
0PqjnktFkX4f3sz8NaM26MJ+lYKsOwI0f/d2l0Vc1QhHsaLrSjipbZHO89kckDf0
RY6mIDrYgdRd+qQwGmIbVt8lrwHHv/UAZAiCtdw9DwfwNAYaZG9fU8/U6r5Tinqq
ZR+kglgsm5J1ObC658vweEsZws/d9Xnc3/4De1xcd+Uir+JO6WjXiMRWpirt7uhB
88xy8TvC8uRyyH/v4OPYPsblNOgKUvMuOYpY/f8NynmZKEnnN5bScRS7fgxKM5el
i3RZU66pYjcKs9eyeIcQugVIgEHLdZpfqQJ+W7H+/VJDss4J5lNsbR2IbkEOD1Qt
en+qOm5lUC995Aqp84mW20SOcA4CR8eXVkrM9Dwg6xSaTdonniIiTkAPvva4ec15
GVAX3vX5M7rNmK8DanG+1Q028Lo8uQ5TxWufSxUf8hJPMGu/rSB64Iq54K4cJyLm
tsXB17KL2kgRjhmUb0vi+ahO57rZG/UoBiV2hUy4KfezjSw7E6TtTVl4dN9R1dtL
fp5uyFGFoPya4MKAKGbb6WE+RY5vLzmKot8C09dqwC5XU9pl0yTAEuytt8oECIBf
DMH8gE3xgW5ThdF9pJQboahJrpbECHNTXkvLjfA9DViT8zcHwFvcUbU0O9sdzBFT
EOMG9KawF5Rzq98l4Ld50+V8OUhFAKIngPV9Iur86qbA4heeEJLDPstZ/k8aHhU0
KYsvV0I53leHypm8eT0U+cEn6s1zVTCqZyToQoRD2+5GRa42+E7Z8Xc9oDuaJnRh
4lfB9FXnYdJPSlDtugj7yiQNo3E1+X6mwr+pJFofyl7PZx01nXhfbIuggjePMWdr
jt4wFAwafaI+jr9EurXen7I+9PTDDbyMoCX0K+5GDSNTYJb7BstZGnQ6vGbHysmu
HmW25O74l52NWf/rRTgvLz5ZXbuGjpT/OFc+WzkzExRr/qbZw/NjXkzJU07HPnU3
I1jod4SKXTjH0YIGm9nffj8OyqCW71p20s2asXRLDLaIcq7BGZhKRXmnDo7xxLIJ
sC3h8+vEqUSZJPxdHnQ61fieX71Nvk7cuhnNxITdhyg9aNd9d+jKWLxkSY8WkNmK
i4IYmE7sKE9J6QtH1TNnc1GNpi7iH8FK8gEhPyC7uFmldcfZHcxM/V1wYN4hPxmB
uCg2E1APZx2UqUZASzy+jXMPwdNX3zYEwjRbRb0yg2MAyIQhjQzVGCO0RGNWg4O/
WqzfYlJu1dS/TvawSV/x+HK84KwkZPxTEQe5giKjT2gAg86gwSaSvo/98Kq5061s
Z7cZ6usfb6iUQFxR0WWyMoONGLX3ebo4D9/RiCqNrQRG8D1yKdIGBnwe8LV7NW9s
/qR6H+FOn7wYigygPCWTmrVZr403pfuyUZ6Gb2TlK1d/uAGqRShe++ogTCynvsQg
jlTRgCefr5QO0HxLCK2sG+7WKs2Lc8UPjlJRayp/s9snz3pboPl8l+nuoD+97V+V
zXFQ4T5Cncn+wfx0U3TKvJR200C0ZuTAK1ouDHyL7sI+exUIevOQExHWQaXvJbt5
nJq5k5vov1uxtQVBzt4Jm2JAWttEzrrTx8AiSdoowb0J/X7G2RsV01Isf+quNgX1
8v990nqM8YJKYptWGgCfhky5unSqcW7kef8Ej3ZT62WQmzyQb7BKCFZHZOdh4gB8
C8HVgja0/avU8NCdW/Jq/PQpRIikWyLhD1TD3b63TUsaDpX7NgorW3IKXFdSNSHT
q//J2zeOrfkPwO8kKGlt5sl9SuH2lx6V4msXL9KBP8XUzuPMjNrmjsuSO8GNRFod
dUphWoaIgubRreN+9+zThTei3m4WqzLN+K8gVNh/8GWVWA9oVyIBqfrfwwqPdgYd
tGbBmq35j3ScJDXpsWnuaXA49fSsZAmo15/8j0VfSJfTCLbH1SjSSNRpAM/aRAsS
qfojLA6boKs6FiVIC2ajtlAvioaNAA1yZciEqdAWwzgfl1iB02Rhv7xlyaOIHla9
DH61YkWjE2j2pegmtaMB+H75N+9m/o93aqHapO+vsPw7g98NT6vPbd+877jq0d4t
Rst8zN678DIMCw5Q/YXtfD90N6IJpYLfiiFCLUwkJT8Vw0eZl9x7b2i2GQ5EnSUS
3F9EghWCaTJLWtUL/oPDR2xWtA1mXAzXOyczChZuRCKdcd1k3+6/pOv9MVU8UqCQ
+MlH7WfvwD0D0VImtmxTxl7gl/2VSqwL+KXL4ky8t/g3Kgtg0yjYn3Fq5Hc6/rqo
aEskI4K4mOQ93+rXk61U2usaoFffvd5W/cStCqMtncYLixKkovFZApr2UscLYLAv
tBLk5ijWYKQ3Lv2yvO2o1hBDS6Vq7p0uomv6cn/p1hzDobBDIWH6wVAn9w/A0fgI
3PYzwvqE/mG2fT++jPgUXRGfbOGr2guNPlb4BRqFx1RoyqWPzBkDlOCuJMdx+LtQ
OXBkaPLlgZRmSGlQTFrNDgi7pVOB3scOtB1L1BlMzVrtsGDZPAsdOPHaZsXRnC16
qj5ymU0oWEoPqPT5I6J6Xj5fP3pTiuXAgQBvA8MLLRCM+fr2m88BRhgACx5sIL81
ZsrIgH7I/eUdGgk6AzaoWxWHBvxXlmXvRbCnNXgOGRg45nMIsYZ9SgbI6xAHoJS1
J/pXtwxq0QZspEAIGsSkmvHPK7AmQLwuXQ/qH/rgmcJ6ryGfs1UwZZ9OHTwQSmT/
7ciR7SYTL/rTQ6lZsvhln7UdDoaaNzqKk2BxKp9MiAW5Xuy1oL6V0642Vu3vcBhW
Ku6l2IPx8RD23fGzcptamA+CnPHQsQxlMuHt7P6YSD8cP4Tj3cmHqhx8k4dteLTQ
adXX0EDpvJ+fYLf4KqAbc1Pj4c7Y2BJdPl29AU11LaXvTnprvpdcutxtuioKKl7g
ZE4N7YESEZT1nm23WuqYbvtVN3MA9C+2/GEF/hlD/Srhmq21PINlGKK01hrykSz6
FbF+4/nHyeDmz1zjeXU6QEXf7EPjB0W0aH8aHpxXuoxaViTKFfLTcADhU9MuKcPN
R7c2YtoMUCNB6t8t/Q0H9+jc5q059LM1UAi7H34sfLg6aPpU6kGt4joBlKNgtOnt
yF1hzyOEkUvmwSMzrJ06gRVPbue4K6vfYvCFA4HO6btGZOzGH/SpPQZ+PPKX8qzr
TjOSd4YfQBiY6H3o6MzD11yJwFivvhLRasN9L7RE1d6m84j9vL8dQ5qtud1rML53
XQIBfBoKm6s6N85mYWwwktThsY0pSoollnk7+A7v8TkIObgjJ6upLppvEAmNSBJv
daMl+uCwrWhJ5AB6W0M/lh3HVk7bJyPbGmsKYDrMl/Pd7ZFCtr2m1vCYMcPZN6O7
jkNZ40fL59V0kxJNEuVJt5luDc2Jw0rlKRT8wMAUTJheaE+c2H1XmTPwUL/tcxto
K4T7lT1ZiBqpkhNaWPgRSAK54XnmVT4biz6boCiBm5fHOR560Z4qopOgGsbIeLFy
SXYCq/4tluNreaDB6MgyOh5H8963VB3qGNwKX5wyefxHu7FH+dHQRvbWrR5UsLGi
UGzC+y8bLVrlqpdQR8Z+duLWiuB7/eYp18VVMvB9EJj+mJ6kGlhc0CR0Qrem78Va
jZNlauKzvH7eGsvJjE8XfEib0JKYwsDHtOA8/l4RNgxnohmNyM981xeirSmA6qBG
KBNQVOnGA8SEEj8/nVPXsK+oOOWAqSCR9rH4EhUkOHMmaBQ130Cy0TUC/uNIdGVl
J+IXEOqdw13GxWNBmmS2DIveyKXk19slzOpwDL+a3ZN/dZeppIT1Far11wci1A2q
Qax+AZwP+7HYPslmyeyXVsMRjr7+zgnPcuG26DW3wflcw/uP9fN3qCvuM4rlMLkr
`pragma protect end_protected
