// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hm3S3ZbPgX6+dHH5fJnmWKv4jVw3LDI8l24fny5EIo3r7x3NzZ+eM61Yw7xGCPVY
t1kc3RwvsnhpGG+Y139Ktzk/WhVGSCwC24hy9F2L3pFlWLCXhfI7ODso5tduWZB7
Zp+N6BQEKu3lO5KrwRe+z7JenHOuWIZNKu6+svfbj8A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3712)
ZfvBOUbt9SbPRK2OAdckr0QJnYqx+XRIpQ01qkald6qijNauT+kBT5cuOfHkjumZ
+sRvp03I4htdkzHweL4rMtxjqL3wr07UWpg2hvOa5puk6HJjB4zguW2eDZljrQuX
5FjTp3sV5Z70rLnHnI+FYXVXHvbJVsuU+AATYlc0W/2MKGodYMI8IwClRDEZ7yL9
1TG2xMcciQij2nxR8xCjH8nmgUkpQgxxfWXWoqHn2czaoFNqA+qCFi9ryAlJK4w8
2+BkWKxR26ihvEvpZf+BQnv9tmRfpvCah8lqljv4igspZfWCrQw54UxflXKNcRmi
iO9MCkjfrd/U14EFsT5m8sM39680wyMAQVZvzu4M0B6iB1MTQPtADvqG5UxQ+aRm
wy/f0F8/ne8dljfTDg8NVEs40XF1uYWAJ8pHqsYAjMwPmSrL5zwa6FdfaZy4SFsR
sXQn3klS3sir+lpBh0noVK/3HHwxVodVosOoxc8cCU2HVTbmcSuN9oVZDuUdQgr0
M/TXgMKbjf90FHH7RkvbIkXUCK17D2/bmjs1D7mK7mDF/mP8FZF5bDMtLpn9HQVW
wKEB0OZV0zqhgOEOcabAXpgANXqpM7Lw/xt3QDQFhNTWrQQPipA9kdKboGsaBdtk
86IO50cvn8gB4EO0fuRS3sJJy/VaMcA0YkzqZq0UGqIi7kIokWmzEUvdl7fWlTeR
GtOrJx9XfNVUxv7YZbmnDzucoUiDT2n+m8LMCzB5ONHPFgaFuZU4hqv4dYmELhfA
LY6qJpkqmYSrVmk5wkDvccE1SGLV28f7CTgJmhvtlQ8K1iBBaPW9gkTrLCsGiG0X
sGQUnyvaWcCkcxq7iD1OuPDUImERTXR6b3Ujjdbj3h031/40g03kjL+0YVFDR9cJ
aptv5AkxZCDrw/fnsuBvIdRk9vphh2N57Mi0qyLCQseKAReFGHPT+wdzMct82WTj
EOK7dLrfb/kIWvKBEAAYUCgAdpdHaUmx2m+4lKKkSa2VOk4b8veMvj+hWJBmZu45
XwPeT6zIAAiCbk+arwlldhdu5IMjOexvjPt3cU8OP8KiDAt/NPg8S7/eoyGwrmUi
ywN6kJbl6cElBAB4apkvRY1DpOiYBtSQYzPbq4oH9+sW0dk0NQAE4PjvQxd3z7lK
EGqGkUfXihjPBxEmib0whR89wIkM5XTXoBlgQXhekBLcoYvC9+3I82bfyUZ9mzq1
EvADUtEh0jJzG9QfybUQpH1McLNxWodXdU05QcdeEyEk61MEWYIT9HkRh5Otey+t
On8XkNYChosJEaMTY0F5Hcb0SdAu3TD8EVIUCr/soLU8KBVXjyDR+fP5VGLxBgAS
Ji+0NvXoh6VITUi1hS0YA7Hg3GQtlPuzfkIkWLhJpHMb9gzDgF20/yK+YgEmT6PO
Gr9PvgkHgW/bOAeaeJY00pXl3l03h/elkn2o/33T4a+Uhch9KURaFaNWRbjtw76t
YnOg1FMArVorpS/wfyCOnqTK7DB3fOqR86FjQ4GYWU+Y52z/NQTb/z+lYc0N8sZk
flD+BRIOCl1Qb5NPYqPMPITyT5UXqc44s90NpNk1JoK9vfFqT9YIwWpq0QPMARgk
BdDHmMxAT4Zo5bSsPeOln8dVkMzHyoHcTLgUDyVyfUX8rFsYDo/UdBfu0BR6hNWC
jA0dcFI4Vqrl9fBaW8696Rj3lIeq2nNUE/J00bgjBc8vKd42jLrNdxQORJF+XqBU
mR3Z9YR9j8D+dzoElxgeG+7b66rowyK/PIwnGP0YOnHpGZLgGvSpA95Wkq1g4qyR
FgdF3tfgNHd6p5y2579R3FQ2tXXlHTNWSao3DKOqBvFX/AhxddDSsHfbweSfmQZZ
WrbTHcl6+37Pv07Acxlj63txSr+Wg0GEDQ1ZvPFF07WlcFt6KVbEWWWxNb8eex8p
PXwRzKHVaLSkUO8QCXIYsx8ubXGBzRGG8sxgAZDsLjDm7RM9uRxf9G0+aUEKNi8a
82QJw8gUQ1+DOe+4/9gDHga+NNTVoRsVDC+HcNLJNCnbxzHpvU+GRKHdMgnTrFDW
1orvLcg8JsTD3it2jqDtIxIK3joZOvGnIFaMsKf7YRfLOFZQ2bkNtG3XMT9c6ZFx
kCrUD7r6bvWW3c7gdgi+A201iTAganVoAU2ScZL9g/SrLN8VdoN1OA6iHVcpOkkj
4924vdXLbfEZlWqBqcQ0J9m4bcGqaQRI9GyMuGVaXWW7F/76sP9yLROAgshUpTL+
8QDMRnLIcJEAN/yYt6aj8IrUyfcgn550ZvnfKHiKbu3L+8nPTapOQkLJbCe0kzXp
Awl3EjVFkUz7WDB4oovV2n5EHQi+WdnfDpPQyLdZlsSSnKb/wC9S05pk+e2ixgSx
SOdantkvg+tbtVHdz+eedRWDgUxbTbMWaOcsA+HImyNFhg0E+jl3crcoKffjmdq6
I3ArXB8XOLwb2JoL0vcypQVEN7WRpR/tuOwLPJMhdnoQ6X30xTzZ06ABGJ5talpa
q5CO2fUvyu4ZS5MumnXpHDn1LGNS890Pk2QJdVTLOZdH54UoIyObe6h6YOx6w2ZR
mLjjV/RkJcnLKtdZxOj4Yt1zCDLrIcziIeRBTVcp/UxU+Tws/rtF2d1F6GobgdIn
Nrcnmxo/8rweQeCEVnBgoJi4/LsQKqxEdt8nDRnAM2Z4we9Zkq9tae9vufIcrxCi
7vVXDZFJSjbQvA2WHabes6Urwj+LbPK9IpG3VekNxQYD2ruoo4YNuKXV6Xg9pw0O
HQQ1K/NP83eI4zN+8U/aEZJOhcIULC87H0DbF0cupTlJ0DAHjpNRUtx2UL+CssJc
ibOoSerrT4sk1H2C++933gROPgiwi7ky3J1qg6dQvS+OM2YmjV/pBiY6cZvC2lTN
AWWXLCVjwaEw+SfZ/xIl6/brWwZZHmrkt3GBxH9dp3NhKM9Ltc51Riie3oZbhApt
nVLDJm92tnn4HaVOoYjeSp3Lwj7GhB3ylC1Xso/9mDAh7QTsKN/TYrcmGKCb2ip6
tDv29qbhcj8c8U0Z+9cAWpXBHRLJ7QxXyDPkpbQRNr7NTyOdfxHn7CyRa564/lTU
A7m6+UO2NyRyr2Xq0UfJteMP7FrNzhU9Oczcm7Qjgxqn53nN/fgXfKXRzw2fa1qV
bn8IIOXDPjzpGGi2K4hLglmMfCeXJHvKpaC9OU9Yi52XuNa1Xhq4MoRfH4h4IOSO
OkuIBmZZ6E6Wx7YkgGioNYdf+HiMaD3sCQVWQSmUb5a9xqUjzUyV761vditCAzJ2
UzU1SH5B2cOeHNX4rb0tkB6uoehhwUZqNqEpl7wbQ0CeZKPobxh+pqO7ovEYsdD4
Rg8iiuyLm0cgefWDQo4bnUCFqYa3j3S4E+6+3W0NV6VhW3lumjW8b40DlYtl1S/+
//6etWp9laxhdVOTr9rovPdkuqUnwDgxCAUHf3BpvsU7bYvM2+UW1ZqUEo1n5sAr
5HA9pN5lFw/pzjk7u25c7ix8TOHeHUMpEnyo9oNuy2P2YQtbbERmL85oPLroXFSo
iKgqkx6a30y30ODdAaJ+5UFs5MloJSUP5e1tNgWh0FBX+BG2i3w68S8dYNyl9O1D
2VNvgM6adSwUrS/fwiSlfx6yLgF3FKYXsP2PimkK0lCD/TtLrGr9Md1q74Xbs3gC
l0Bd82Y2wFDd95035G1vgjnfT+dQ4ZLlEq+0Eo0D4Iecq7FXzpt+RGJXiM63I6aA
lxihSBaENdqhw1JKRIEMpQb3s61XDGCTSsex8rQEENGHYVSgnuMZmuacWYZiSncL
U3bNEJN8eWCuT12s+0MQIggyHVEHnJU34rs1FYPZ26ZlCNK9+9zB7JTNthSIJMA6
sdFFBZL6G1UlDUjBHIPIVdRNIS0EL7DCrnxjDqMCJ80m60ZUnFyXqDDZi02g0/zx
3hQYok7ucjdO/9edh32ungfzoUU8MZSczH/qMNrlgWmtPEjhZJsZQXU55cXEIU0I
ApvtHJNclWIPeZzLZ5qtRSvVG4r+0H54PDCb7M0UQJcFLOWWR6g0QBynViil/wNI
8SbTOEtxZnwOq9i+yt4c45oKXnEOnp3XTGzhkc2dV9UuqiJ7gNvpC6f00HTIzq1y
PLOEu5bN6p/UChJE7pCRn5hpK9ld6aUh6H00JjIt+F95wLoN9dKaNAVMey74yQFI
GfExLRnpwNXEvdmRM5SQC34EYOI0f79UfYFwaH4a7C0fRMJ//DUxwMkoe7LrLrGA
soB0dzY3VjU4QBZa7K0oGLV1OGWyLGC70V/XM1V2KdK1FSnN23TyTZw0Kk8gh5L8
s5UwP2Pg9H7Lb+unFZgM1DhHCRguBuBpCzWpd+cLepshe+0JzjmbeXZNenzDuGrS
Pb1dydX1pLM4i8reaer77h0BiEHShRGk5sZViLaVMe5XQfn3kDDADIJYCcQz86cq
FuINkESHVUm8VSfYDkLqiMn/U6wfoVog13conm947JdSxsRZPYwI9jGQeU1+Tzh0
9FNmT6gmqRG81pZYIuah5siKke0rhcFHSxpcUdq1qfiYCJHmG5uoEpN2GNOL4BXp
tB3eeqaaBl6AE413gp37v2O4nyeSi4H1zeaZLdbM8Gh78QcxXjfGPmb2YxOXunJP
O6tCxT2K+2TPfvP0T8x8cLcJh0To5Z+eHuFVyvHmbTKoZDHdval8/JlKFq9vymxF
366dvPLSQmEvRR9zSagftf30Q7ktaaJwGuQlittg4IVyKKhoZUPc6Tc/4o17ISfr
mbumdg+RdTneqTOMHsj/CONeH3jTp+LHBn3xu+Q4ogsJuf74FK4ct3G+YzfbeJse
sVWrRq8GrWzGovy/gwM/jwkVluE+2S+OwUfktNBJBYpMcmFWUZcux1f0xbZboS7b
n1axV2TlVEt2DXuquxKTdhY4R9/TZM4ZPmhYygSdMCI4g9Updqu272/kkCj8MzMS
PKw0378JpIMwHSJZZMWUCA==
`pragma protect end_protected
