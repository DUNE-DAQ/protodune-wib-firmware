// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
anO5H5F4KUIn3S2MIawHwwuG/gQKoUbcRx1sXrZ0p77ou9tk2SsoDDWEC+c14wLG
aBWww0uJ8Vq2Aa4C+rtgxiNRe/pu7yH/8dhvaQ99Jsu1SEfVOJn8La9okncCf2zg
+FiWhV0D0sjsqElxchQNulcim3iuXWLwUetBeI3NAks=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11376)
VoG+7qPXuvxfmn5x/3E+KHprTM5zZHJ5MYNbDWmDEAuc0yMvZSMytJ7z4xkBq2Dk
oI0+AlR6OGRNVYFwHEjbA5wj7jufpMVOC3Wwijy3N8vyPl4hknt5etWjAKp34VF1
2Ndw6Ai0TUJPXF7pfaEApUCd6aVNrCCHDOJ2Fcz7lvfYzvwmG7gkfylTAjEAl73D
PmFgWrx4mP2ZiDpug3LwRQpkCupBsaOss7r3v9qYegn+uPNYSMFd9CNOD+c0D0gm
Dy0RZAS7c26ZGy10tbJoIT2MkO/mRrhBq433lWfc+we+UJCXE/IhsphWfGkJ3bmI
6Hq8yy/63Q9quDhEavqkvjmWZomtIJkyGs0zZ4ZyLpjhtjuPCnXxhs/K2eracb93
T3z6batlC92PwYgwZg2g6wS6uf0Vy3A38GCpkUBgVLjyHxyJKQE5k+hQgBf2VvNx
WsA7UdHHKfckOq2dbNKEy+4jw7wrxORnmNOXfZVk3CVJvxMBZz89dB39HaKknhIt
oxxvhKZoPFGA9KNLmM30PgVVWtyMTRwlg/uKsjC2Lfjv4plAe0AcGx7EZrQoqXgZ
MjJ8uUoqaDY9yxea78IlASHvzBYAkfzomP4gkG68EevykSUkm0mJyQAoTBjpscG/
2nVmeKyqsbOfbLyBcjP/zTHKHV3K3KMp0oV/yKAgyQr1hsToXpEBzi0NSBHd+atF
Ni9YdIT6o+CG0ghigl8h/HwrZsb+qWJVg9FgDVijOTKX4rL9zP3t8JrjLB0h6/Pr
z1/Pf3Apk69deh9D6CWQ2gg/e/SturjK7Q3taiAm13eZpzAQ2l56xV59sAoM9Cwg
urokwR5bw5SMS9g+YqHqWnFuaMCLuhtQAfynhQuqykdLyE4A04QkKt/YZ3CMCtL7
4gnRl/Q66zwSEB8hdlVOQxZDI3WCepjfLchGR5CF5WkldHllgw5TSyDnkwQQ0Wny
GGslf/hri9kwET9B514M78SaC18Q6ZPkG26HYuxoyp63XeLzZTtg9KBUkUI1qzBD
qTS+sxVWJYJJh6abPLmStAlghO0lATk7hI/0eHwg1eR90pS4ruHySdD1HTljyO1n
xy9xU+Gz6QteBvjMHcR0lqlU2at1z2TARlXRN6pPwM5HBC22hFKaONTfb1K7Iikg
EnFWiHK1LMThmGryVmO2/Abuvkft52L8rAhwN0bwwIXH8SPjsoGvxVaNwwRvg7mj
Cs9hgHuJLFjeFGWLWqLEnOg3whEmqrUUnDJNTCkJ5FiBROT/qWyeqiV9W4AAOnrN
OJGc/8Qb5gBfRlw7JotW3Cay5Ck8pLpPzlug+CHqjyf2i7lL3XvHAK5f4ZV39XbQ
hH0FeTB3FCFksnLmHKDesWFQeFJ8cBLcY/WaQ/NJBJ/02qY8IvX54KvYYLEttmxt
ajWNqGruy8jHKDe71+g7hEcLi2BrWre/0JxSKxxtpCM2AK7Mh+kNEyBJtPI+NEfP
uyMS3YGjKzSF04H3OTFi9sgYgZyKYP2gMa0EVN6rzjO9sZ//0cySKETo2PvbifJA
Iow+m3DpQThDwoC2UiZ7+wsVcH7cPsskQBxF8jm0R1/IfyraKCTla9yejVkYMxD6
JQpyES4d5KGkaYRYxZ3zHKI1H+zjthxjeXjNDN3aj/q9S654a/m3IBwdMsrhsRs3
zpbV6dQB7wm2um6LDygHQ11ptsx1D/cZ5Y084S38VjJHIXj2cbeo73VnrCfk4bOY
nJ+HgBIq++ElbdRfszXXI+HxaeZH2f7ZJT+VbgzzPPI66smVPmDOEM7bVwTJo1qx
V2SJKbLHvYMsi8nYv2XsmPRgc5gaMWijAd0o3c4pNeVB6rH4551w0K0OHLf5oyuC
zg+r8y2VIbfia4cA9PvGgWCkbOBG7xVQTb+zvCdU+qY6DJ7zxHs/HkLlxvrjwYux
kfHu7eeyKZg8vdvs0e2yf3J6AVmPp0k9CpFRX48mCn4ftF8bwDgPwyGNaNLyKYht
ZWSBn/FoduziKJH2BxWyCXtT4jSYPyVgGZ3UA4NbRZK5fmccvx91RcJ24EiUhaXk
hRLZEjqpFSGANY7Iv5jZgUmPp1HVjcxCQDAkqPvT7SO0aub/t0w+KmOeX03c/HOQ
A4/fpEuy0SeavQd6SVEKikCtCgxVxELa2CL729XioYI0viYa3iXkP3Jyqpks0wDr
Os5DMfdIVheonWo4c5FJSm+leBQt+F96qNCPkVhWkTCYfZf43MD7Q2gyyfj5Dn5l
93WNN+8Epfde6XBEcTLUMiVhHJQ2JhumjWU2eIpMM2m9yzSiUz5CRV5WC9xC9ARA
YidihCOUd28/KQCOBGe9Dwap3lzsfDOtQQT5s7/o99oso2duMEauhrzzdevnG1pw
Lmem+mv6JUmrAntXSgiosVGZg9QBSGHCgIg7qt4XAL1HsVD33TJ+LKC0vAdyt1yp
LkiLHwTBB9TuHbiDntVvS2JatSaZ7dzmQNElsTfX+Vet7sEugnq/3ArcQe6EgWvQ
1kIrMXH2QIfpB4WJ9CV68Aug2O7r+wK8vOPaVzC16Lv6xp+UYx3m/usgp25nPUoL
kjdZmCYfxLGig7DjAqmJb1PBODSKTbCg9Yrv9YLZ/ZnBwBRujMVGYMq7J50C1y93
jA3DNy0MGIZyQ8nZCi2/p4w9xaIIWifkyEgql0w1PP2r1eeAzEhl0vpvFVjxLlVF
RNogleAQ2oheiU7hVlGfW+m+fBVdS3aCe5QSOXiGfkHOL5DP7sYNgt1AJn6mxli2
ubhCPZJGTuuQx8Rjr8vNOo2wiMD72INukZ1MVTFkl+WrSZcH6jMlWC1Kl60IDrlx
rkBwVEcwdNzIUNv0CcMkWhdmlt0JFccc7CDJaou2vZUkuNOiSJkj2+OvepTdppQo
4mKRqPjzIQ+zan/xbiBDOEEXkR6h+2aGmmkn8hLy96MqhXxD9lYP0Y+mynqVMXqS
C+0PBRdlZCKQxHLk277rLhEW7STGGAkgBVQJ3ElGh/i9Om1b419h5CP3JgKbKBsC
wfROVPjOEySwLNWQfmNKdtz0T/INNLYilIseAO9A96wbgMgNKvCqzDPnYJyb50df
qCgTzO4vP3lYd4ChWNa7u2K8plFSb7g7Hz1aSNeWEV+mqy6CJEdVM8E6yW8ATaYw
7i3N6lrlSblsP9cAowoLcoAdTkGvD4y6rMk5mtLCDx8LMz1nlDcQxHv+f8Dh/mQX
zuEi/Qi0ZqZjRROH7MMpEBBV3ad+HQNR4/bQjeitAbhbEak+aYGifx/FWhSv8b80
rJ0aQ1XNzESpR0U8azEa58Q+86iUK3MQhqF3kzrNeUkGnb70E1yK+rwpKULOtlJW
NieFom6OYdYyAMX7APB8d1kfWeOR0qDn9Yfvh8/nyAyoLMam2vp1KvpJfaFQlWDE
8n+yiWNTzZ6sDmk5tlxEbdpZ2GDL/e3LrpqVUkSOD37ryRXVHYktS+3oKSDiowBS
bkk8vgo1sO0YgLspbuJypKzxNwcPBJaN780v05caDNDga8zpRGpCQQEau+NSQr2d
tOcpllyl9TxeUBn2qK6IejfHY2gIGggL1s/zjj32sNRF/KCwNoeelaDUxtyRLkgS
YumQLrcFgygg735lxgYr/YJlKX9fu4LpQ2mF8DxwmcpAo1w8U1zbKgvzkqR7e0/2
XHNbkOvJ03tXEu06MVCuMrENYtCiX6OLKXQAfI8lIjpm2AB1fA3oDGmHId3DhP+x
UaAtyAz+tBCCOl33guQBVI7rKoKMvJtrCHsTkB2WsoffN/eDeMNUGE4GXTxfVtaY
kXXYj8et3YYLv7+fGsvV7Wb7OJz58ZtBL8gWtxKrbEKWdGjsAeJh/pczK2jV3cKt
5dcFq9syUJE+f0cV/qx6BbVMa1yFd5F1DELqmixceH8IcK4fH+nO1n8vLmaoGeUV
K/BxL1RJ2B8kou8MIlZ+HWEEBs+44ccs2AQAn1iHXmvXTEVsZJJ3r5U7jroBACFA
2a7otDpN8b8M2Hz6iApL4xqgvzF7drU3fGYOK1Yvu2piND0MqreKwKHEdzWUPOk+
mRHx+EBRkRF/uutdwBYi7+uYuRtdHs5hh1vm54rSinCFSqmdg3iTtPKZzcFfvmtG
6Ra0cF6KDPw20dzK2B6fhS1Ecaq7Vl3YHRkREIop+fbkLCdoGK/Huco6vZRs2TaX
enqriY8xZfzsPZYMZrUBDog6Mi09V/U3uPKMptjnaPIejwnzzPymSJz4RyILRyGv
VKJ3zCXWeOsMY6Wqylo7c/44YlPhTzkwnAuwxLaFj5dky9r5iwq6E5KZc1UNEq8C
IdgZ0GWJ1mKgF+8gqJzMnGBz79ac3VTJc9t8hngXY7QNDzuhqPjG31qb4dIF/Jzh
9+RcpTk7zDp9qPcrrs/rJ7xcbryVJFiQCKTWbTV7wAt72No/fH/MrbXF89OUe4PR
U2rK0KrlAuR7TORdqiB8tExLehQb+ZQbH8dmbYJpQWfN1hjJ7zE7n0qhaJkRwkiu
sWHZST3NSDQM4Hz7ZbyR9JNctjCt+yqNFG7Izo1f4w+ZkKP8XYyJGX0UvVUrqxax
iRD7rDQ3xpBlNpzwsfQeFrZXSyEV6/mk9AOHmfDaTTbbYpTETm8StCUHd3Fwfhty
SHoMYvLTcIgaV08xU9FtnJG/S4CQucMnh6YCViUxvrWHqxz0OYATBDVqh6ZAlHPd
s2p6NIKP2oRcm107r1FJFuoj4CsLcHNCzrq320rWFEzXTNYWOoe3t0H/QQPC7nIr
Z9WpxHhV+GRVSL3Y9RM72SUzC2SkQerNnNNayvhP79YBcFzJaurtrgU7Bjq+xn59
6DvUwvgok5EkBxVc2vA/ZlxDj8npAYeet/I+8VcM/R26zFEaW+DHqK/6Ma57HqVQ
e1cBtCKdESWhXIH7K2ZG1q2Q1yDnSyVAiUdiupWdWg4R8z3MOe7rXcNvGGthpWwt
Vle0RskpzNnXN4ozsaffQGA4Fk8sdaNpIZqiYv2mZ2dij9ZNf8iW7f6Qcn1PBLcG
U3khgFzmJoiDMdPZukv/r0IdQNokEtjhCOSr/uj0Ol61Hop7KLEym4yteJ6Xv8PR
yQp2qUJWphzPJ/nl1N8oQfs1vw9DRdUtL3P5DrDgjpraurVSITBO7yEVO1sA4nUk
7XaWm85wJz3BU8uiGdB9rGe52PjNVX83fN40DHFCRlBtqICnTxfjApxSGZHMovLc
5XK9nOTGnQULWoS2albRtgGkTzPBfxqREIscZMUHWQ9KkvqjZkhOkv2olfX0ztzy
i/r3lCD64v+VZTuiXQUmkkMIsHjFFZtafq6NpMtgwZX67Ue1rIxDwFbE7hkaKx3z
48qaMYcCBbdz/hSL59kpuorg39c3V+0UJmlsPWWgZj7GqkbQyVGnDqRNTOU4O0+t
47UgBfeWxO9z9jmYeQLCO8kLl33wu4mEG8fhmRrzQBgN7e+Ubm2lhIrDFwUOigIx
c422uF9d4GQj5S/sifzq/WhZsi3Qi9DgAWTxh/wm6A0ZhPvS2tuU3Owozct9Faxy
Jt0qJJt0g3CYD+L76W7BfwkwRJnZsB5Wnk4+XcUV7mKC+BQBWYWPznC86GlcnRv2
ZKT3NJpuHEnCRGsI5EeJX13vogCankBodoiHP70CJxGN3QC9ghH8DLaU1tZ5vCSM
pF/rzhgPXbilavvBzdHWAJIIeo4AwUvHCwybFbW1YYLQArwNPF9OkD2F5A55HEam
Bl9KpGhmLCZ4IMwNAghdxpYCcShTdyRLNcrrfV8plEnk+VdUHcazhQVHILZxUuMf
85wYDUWK1B8pAHrYKTEKvMX6PxV+R9W1XZ9TXXxqbHp23yGAdV4l0JgeZZDT4xuf
5HcO3iUKuAq5F7QzyvXi5sLxvMIF/p4F7Ya7mp1lOD11DIYEUIBpV/+jZbZuuFGj
nabmQqPpXd6IrzxdaIGdMfxax/JPa0dkQ94Qhw4AFtpTH5OpMpGSUXdF6i1cLDI9
kJYNciS+gtsQLkdtsYzD+0wi351VC6MPo1AjYyG8g+L1WszEB+LWGtrRvXWce5CM
E8QjItHdR63iXDCPrwfmBlf/6rF17gjc0CgljHu3pP4X1rM9ClFrWSpRdhi9jMG6
jaU9eWSzilRIUZKcUeF0hQIMPMM/jC34iKOhqZV+K/cc0Nflmp5C+g8bJzQceebc
ErallKs6J/4X/5e4UipWNPkqWADmuiU64gyD71WWOlrbSG7/vdRXjzpTC5ycszig
CODTP4c6lByL2L9htK48wTar4k9Vh3s7fAqfKV4OMCN0eS53W4O6jWwqVSC7ENO9
PjOZ5okSrkSwZ1FSjJUIYrkOd6vklaWHSfXPG4YjQPUnD9nXZ7hkAFv6QnH1Vm8o
Mke7RgWYwwuK985gNu21vkPMNSqO8x+ksBi+ZK+VIu12rWa/MIFPTLo+mE12c9TS
WwjyYPAids3gPG4qbL+j7hC3rfROigcybcMKsTZJF/7gyEdewbv7cLWbX8S4tr+U
rUzFFYSD0D/6YrBQQzlqBg9aN+Pbz0cd5UF7pNOrTYEKhmDZMvr2kOTI7CKb4twk
H7viZBtd2F3JlUE7yZ7G0iwjLkbJ9Y/ImSPxFQV8cRhNhcTmG/ylBjVngngv1buc
+hQul2TzpCYEcUNTunT2IdTHDL34fTc43Xaf5H6/+OHaLtZRgXc9cfcefhjhf7wI
iXxHVb896KU9LYRR1JczI1tuI11KC9wvUu/17SU6nkvIxRlWWzvNgM/xg8yCSNYJ
k7MVraBDRdAE1G0RoxOt9Vohq3Ml1uMk4KLrGLiF/NUQaErOqriPCOHN9Wz77eHX
zTz4nYSdCWYZylgMVT2RRMYobnwnWHahtT0cjuYmzB6va7b2kMSX4E0B7QWZDkL2
R9nCXGdOVCh2/wNmR/+sppsennLN6fN/VV6qZK7rwxlIb3FwnAMqmkCfVKzx9MVq
j6uooYnyfExlqm3yo83Sj3a6bGi7HPp0zpH5faExDaqcj1hSBCPZhIlnZHHiEDTa
KhVGAPG1DtaMdChslr4DJjhSWlIUasRbIZ/sIpgVEqf9amBgYN9LCPpx8U2nFSnF
v2At4MoLAS6isp6q5TmI/tn2nD9uNA/I5MxRUpj6e+i1ODS5PKTM+CTkRMZHSeyI
eIqvmya9wRHFYyKMlUcArGJvqVIuJYC7xpJOYOE8Wx8nYviVV9irNACc3UtvHIpF
PkX7ssuqomruZ6XHJLasFLSB++Qg/IHHVfwRSgbmTeAAdYyDmxcyS2qknJmJn73Q
FIP3cZ+C6DCctq4sCfvN669G7BnTyKBuaj45W7R+gF3a01zBaoLLOzBet2lm/FSU
o/cGN7yJ2ZzfmiqnhUwn9zHXfQC46ZlYTd7FIrc5Ed+BRT58Dfcb3THb/jpk7JyN
cifQcX0ame9cFRlafuGFhqA63vyxdJU6QRxPys1Qlnek6MxneBPgs31BJ0JZJZJL
KIiB5SEWBaAniJ52UjCEGWOYU6GkyR2KwXtKkDBsxEb88sf2K96MrLKdOUZnTVuk
zVhrlgdpMKqEoBCqchMGOj05S638lP4n+87vfssGikTH5vUmPFGM6m7wMgggGeDo
mPGH9WCfiHr297qCzL5nVKhUMA5GsMDaBRWg7YCz4uEVPGxXHe4+jH+71WVyhu/x
dl3pVoHe0KiaS6+bFXcwuqzzgx3li0SbYdRzSRG1I97FZM+bY7j+gg9bdj26J2/1
GiLBdLMO8KUwkyR4GJlV93IN0LVAwBGvhoGQWok1izkRpn1cXtHVo8P2CnUk6FcN
XY76MoMGFAlTo78HGnaKU5MGK73LLamoBzPwlFbtZwxzhc7R1WUhwMMwH5b7czRZ
U8iEDcpckisjcu9oHBjihkA9jvKDbLzkWB9lQVzKpN3MjSwjjHxiuDgpOhX5nbkR
0IWHfoiUeNAzUMd6Wn4VG3JpA5uDFnaf2068oRTc3eNAFKVgNS0xMbBXxwUQ2F5W
4PqpHB2EyBQKqjytLnJFc3QxQnNw2+dHdJlv/pRUSkQyo03wTa7EFSlz85ONW2BL
TNGMbWOTlvT/2EUmLczcfZ4lTGqUFp6hDog/k0sghWeqG8vlWfIe2w7KB8Qo7G0E
YWcnPk0jEsR17TfmcIv9iw8YxEp+l6tSk/7t1EY3Q2RunJCJktVKzk631ocCujmW
VHxni29HsYEarPJCVct0NgG9n9NFl5waqagifk37DXD4xeL8U266somUA6pXV5P/
xsO73aHuzK1HhicHDU8vGmJ1Pp00UkVUFKAq+5qj5EQNcWKM83S/eG5hM22FRPb7
nSPjAH+9oZARW5f/eafBlHrBk9UrtWP1w4dnrPFX1jXOyRZiMu4RGJr4hm7DctTX
HMsBjZ3h/LFcRzR7E/QYWDKSRBA9LmBag4gKGfuJ8pyhUbf7o6IFZ/ctuj+eWJPD
f+eaHgwNZ597j/54nmJwXNKYLGgU3x7Lp7HLP7vsSWmzUb11DL+wbfZGOcAyN3BL
nYeAZ3VriQq7RZsWpd5VAgeK15v2z/ttuu7ilBXeJvk2NApfN09nI3o0j0zyuFyW
BpgHv3fo8f6UcsGjj+8fABPUh0x+muaKiZToJmROhBmWU3lMPSGf8AOgKeCCD04/
hNGjdbB3AwXY3gAHQLHO0zYtCkGiGSaO5TjLhlGLsqJgxPxsu+mFnnhA8955XyQW
IdAY1eW4Xly4ElDrYimrb6C62N6MTSAECIE9Q5egPCRNT94lQzGac+8Nfw2J4j03
LK9KSAAjrm6KVTgYNvmQ0uIOnS9V4JDOZZRbxTiTA2iZmJ0/TPAXNTRc507f74Tx
0gIJa2L4UInJ4DIhmsXTOooQ2S23jsX5ugfCfmaIT/kOOmUCQhRK8NotbF1cD1EK
bX5Orqn/AINHhqYvg00ulW9PdTj5lndN2zKjjybE6O5SknE2O59tvX/i+5QyAWFv
COKxBvr8Jv1VOO79750CBiFAvtt7Ys+7F89eMe0qaxcjvhqdAs0z60ickP6ndz1o
QeGvXJGpp7TNi5IMUwznk8fe+x7PT3GpbidCO0VkB5zT+ayW9S/oPksgTsJoojzf
nnzMZWrmhNMTX3jYblh1xc3Opx08KzE8xTBHlj993+H8EyqqVhSLnuFA/WhT6FUZ
Cb7bP9nDzauDtD+PvPS6AynYXHxiAVjtouAwWDstdI6X+ftSK0Bep8Ut9jNCWbuC
bjAQX3HefOl1tpczvfTuK2XWaBbpwZ15YRF9dq2LYGnGp0f/9cASWDrkEdan71zB
SptieOFJt91XuTNc9skIXtU/FfJomAAK22TiZ0uI1pfdFLRZLulm1wHdWHn8Clip
CTypRykyUnLjU75wHpGUOi5kvukCQeni/Rsk7qpMXXKGyyaC+3ro+SZ2SdQM/iJU
FSa7c2SW7R9+QvzfWkQ6UKsfj5pzkNPrNNBypLCMoO+G1le1GRQVjMGJZ0xib0En
cIUio1r5w1WjsK0ZdaainK00QWwod7i2NaQa8Vud/xdqlAN/8R6JhRcKYOf6EXG1
cClUzAB8QW5B23ectEZaWLJiZ6GXa26Sf9iYanLMbCYD2deSQbyGIPwxrg+nkEa+
A38vxEYvUDDhpPtaMCPoopjARAk3x2dkvHpAsv2BCQE5OND6KhqUe8/Mn2R5f741
ihd5v0p5X6TBK7fnZ5pQBJCCeVOoaRP0TWDYZ1EQ+fdRwxR9+iKdOwPwaFApRADa
KQc+VLUR3UrW9w+fTdeSCfuVJeUeKL6feOUEyVInYnLNOUpKMyySNjZbPZVaxBo8
ZgNV1nYoU+tok2bveaNoyRoE2X+Ug0F5xsuZqGhEzHZjzi5Fp15yyg/k3EnAdGwh
f/h9a6LfCuQ8c6/eoRR68oQ4/sqykzQlzN27tKi/h/oC/4EnVyMKtZ9wj0AEimxv
eR64M4p4CUpY31YIhYmzeDSeLXUW6wEZchbcfFpaSHYeDt5BbCn3wiwNCvH8foa3
nj/efgBmNuRuDYB7eDlrqg250dswcpsU7xaV97pSYvGuSZMxu/F6LTqlPrOyarDM
4xp9ALW22afrnDPQQMbZKPo4O1fbdHRZkRkd8eSfPisS3syXVV5V2HvUL7aZUq2m
PvTKed3Rh+Qnwho7FroBfQ5utEik6LeqKzgBCCywhD2D4Hrv0hZ/Z3A947CxcGtG
mb/6A4wGJ5bSKQIpUEKk/kmLQWIPMwfR7caux8p3Ee5ALfbczTtmmRKrhkoY+RDI
jAYoRpWHKc9qiG34+IAP1YObW6xnmFUR+dpNlar8Gagc7Pq7x8huuex9SyOYdmEt
mn3UmEiuyWW4d0kG0Gk4gIFTPLi+wjj1tTdF4kam2x7myGoJmS6gVpjbLgMdJ0AM
6zVKRh3WYIhOeiQzyLKIKe25/pMuzcD7IWvP5G5AnnavChoVyik90jMVFtczmXkL
orcFQhbWiyanZbGEraqslIxsPiyax+1F6cB5Oz1anYGolrd1tI4khTzwN+hZ+5hd
q0rwJYMwh22Wcq+BsdjN3c90DwNBIc9pwdVeObrzKV2PH0KZhpqVEutU81P6lurS
nyccRAMEQbFykUw3swZDflIhr83ESxauH76fJ7SGRpazw3ApGicd9A9E0HpScdJu
Z3gdSsqh6A/egXD51ebr6XTo2JzAPNZu3CoBGzx6VfDbaCP4ITyzq4sO4UeI+iZH
/Ms6dbw8wYBkc3AJqdv4JQox/K34UuaCzBxQrtF9ATB6l8cmcObkI7NsvOeRWPcl
uOzWgUt0oHA1VXBAxYvHxDcw8rr1ALCtaCEJQz2NwerHoB5r1FPZX8RA9reRO+05
Qn1hrliBZI/stfA59roQtI9BKBR3n+14uyYJzbhJ7A59uXSmvrEkTXU2IsC/wFIS
Hp3DzO16iVrjPy11YuOU0WDVtVQkH6MzFiuZs3rVmBMviQLeCIR5s8rS/bDayXer
Sowv0DDK2HN4b0cV0zdpQ4E5RwnZACXpZ5bJVxmEA4Fy1cT+RkYcs9ravI2JwXsi
BwHnO22aHIr60G/EW2IEYo8xj/c9PRuP4e/7J0qtbX9QetbzfDD97R6lozYrLW4n
pqPHTCos5+aoQRMyLPY2eV5PoxBSPcza3MCr4hfz50DoqtxbHKwvbBMUaP0lQSxW
zgZHR21mf9PWwsGKl3/frgvv78oQizmljojJfMtzHXuNmzoaIg5plpOOXt9FI5kj
LkeaSduMkJc8k+sUuNGT0Ykys6PoVkLqcSNljkhEC6bPL/MO9e8sxrWijt9D9iHo
xgiY9fKgMAY8GXseXKTR2iWmOMgg9V4Tm0+qvOmUQy3BdhxENJDOp6oZUW7LmHeg
UjEBGcMJ6/GZQRQ4lUSkD44Wk6uLRc413zC5hdZpEV4EMd5FkvRmuD1pjwKoSO0x
mh6QV+4JDC9BWEwcYMNnSlryUkezC7pxMECEgPgZfEOr53eFKftz07Mscs8GRRHb
nWpZdiqvyr0v1/2yDVHGwJ+CuQwvIclCZsP6RmwG+GRtC74MscQgk7dAvSUQ2oKa
1kdNXkXteLrnmmlAbZ4FJBrvpNPqoOI6R62G2hyUXzJ3nIBXWtHULbWPR3snIvwQ
fXJ3lUiuPqra9QESNLmI3D4rpMSChbt2ETjR7fAamQR87xmuEj0KeJgef4C+UA+Y
iWK905Gwlhx+aLpAVS+JTwpuXyO4Bhjw414zB73vYHfqxaHLE7b60gOGaJVXrK6X
/OGfcYHqxF/uEBFWZh2CwjOMYUcF+vMDRKtcaMOn1VHpn2qla4WoQ9olzC8jafKx
ivFU9dKoaQOT0Bt/fB73801T9TGVTubLU9lsV/9pu5dhjtXnQp052EsK0wflN9Mf
zvdYVOOu2zte1cvy5PXmHX29+98vzSnN4cEZtd6U8nkxyeUPzS9rHm71ajBBNbEL
mCOqn47S6JJ1y6Qt0/hN5yjkO155qac/uVYJ8XFvmsi9wkqW88DodEJ/8mHrb7iO
wHQ3+zlwsMb0mLgRyFUaNsJjD3VbNtf/D/ADnE+4j53Kpk0hi8ZP33Htm06NB6VQ
AUAhWsKx1ZIOFTDsUwUOd2TOHWi1eDCgLgOBcmIrGPH6cl9zwDIxnRZlGv2IqvYU
Cq/FDvFoE7L9o3V3I1WOR6EGx3zZpuZvEarC+NcGn7BY8G6LAgfZf1EANQoDr0Go
9q/vyxdyyELA+uSvH6YaDMyUP59wR1f5nDWL4LMp+DNPqhy1WI+2c3HW4rwi9hT+
5i1eIuTnlPaO88+r1ls2t9RqvYcUGyBs98CRZxBR5mnRwo0BNjpNIXfAbJXB9lbA
mtpjHmESXMkuxzyvojBRr7em7tyGOVKuVgX6/Nhn2a8rqCvKMAhk/dspLcJKXpSE
vO4Jv+A17ZxBd5yG7+/GH3faAD9Yd7ZlAu1M6/6UKkHiJiILP6aaTuQFbo61mECZ
raLNh56eaM2bLDoV4FuELww1n7wkAphalKgT2Q09ZZeluJfsXGyaw2GInUo9EjOg
QCC0Yn6dlY5Vo2/TUV3QUfF4mR5BIEQkFuxKy98A65cNZxp4f24A8IjX+F1mC1lA
iPPL6UIgLCxbc+K8Htrhbfz2ZvpbyShpkY5sIU0SrIVrxbvaoHGXrQb5h1tSTSUh
Wji4imlcRzhdOHaYcQygXassPGOrLGUcTtxkn0OPJPY4EHJsp3M5HvPHVnlcRz3r
LwTmFUpRZfBPZkOsofy8kfB9Z49c3gbbCvWkqGVZEZEmy791zOxlFYElZ2rczvag
7gQ4NDyDkJdE9+PvaGv703qpi9qN0Gvvj2J/v3hYVD3RJeWaPMImYTQq/d+Z9URO
EYrw9J6OZ5i7JW5Qd2Ua7NG2rweo0TIeLUKWYeIDswtte7YikAE4ul5/P7dFi0MN
rhKcc770byAWQeDkVMfNP1isMbeBdivKxn/mcUcdc27f1xYLLpvWIaKM0QKBjJSb
EsrMtGMQSO/gyhFB7AM8+EuFbnS8g50gX7k+Y7n8qrPF+iLCQphde7XtxD+Zs812
clsUSyv1FDNy5rPQbecFDgiyFQa5glGSBCprOC+anf7uWBl9qRHZ9lOAXXL7JOC8
KLwsqSp/sshGD6yL9lL8DfpkkllZKPbNIwQyzwuh+i0M5iR2+9W2FwpsHD0luINw
uOJiSxwiOelyLwVzwYy6BY8dS7Z/D8PLdZ1EfBURww9vuohJwpmmg2mw8Tyy/aXs
DGyJm+HCgZUup/Gx3NUZ4v8OBPyqDBEImRLp/UZ7lQP85qm3kiLuM6CWaPE6LYDN
wqncDwgoqFeewk23/AWy1BSvibHQN36IdyWpqqHAHFW+fqnUamRjWbP/S4AcK7ZH
yqRqrsnBxkLiVpqO6t+dHJhgO910vno/65bHYbxPCpSU346zXzE7QMVTuWpEtG4h
1ura57PPSJ2W4t3QMPfFpX8G34omXOctkYELZgmxrx2WQj0PQ8kqpVOulGkS3kpr
bSpaXgdt78jdbVOPNBckrL5gjCpVdQ9w+T0OlWpTP5/LBAMt9/SeuptjjD2f6x8O
XFwROtBET4lOtQVXeU4OMgUReN50dR3IaofxZ6IuLenmGJ3SQeu4L7M2d0lV6G1s
eOd3JViCfg7HAZfP7IH22VuoJaUvL7sRNyZoJEGomKBMI0wcgXE41VAMvXzmX3Pn
M5pG0JfkWIxPfzY0G9Rth0TQ1YWKY0WWA24MwBCNINXAReQUhk/vcTY7kDM5McPa
jofiNLf42zzwWWDFdZ9r5K6uIR83CkvrEB0CDfUeQ78HWsE5TkjCW8rm2T/T7Izt
mSi4dBMFrJRQH36WHdsd84Y2kdX2/FRQ/bp4DBWS5FxFuaOxRzR3bxX8SwoDFaDX
OVZ5UyQF3BAkPJAc8Z48XUgGxDSOWOPMdsMgitUJrfDo87eH0dprktqcYgWzCqVL
F4nMPGKf+OXjwEdCNMBJS/wh0/9nIN/MiJl+GiX3RDgNMf8noBRehWSFdK69nvnA
vxGmwX8Lxvm2G/Iv627mqVJq/MyEJvRpp23w4ad3m1WZo6J9SToxtoMXPrh0/j08
rBvIMtN2fdwWzcP0W7Teykce8Rkg3oKIWtvUMYU/KrFujnQhByxgDNuWjpnUarJW
svGggAzvS2yBw4+X1MjrV4FYPGFb6AqIulOlEaVZ4iKkpPmLvWaH8qHTWgMoE3ZE
tE3H7lKc01zLlSnY3GvQ87u6gbz3kCSaRPw4tbgGMm0TSPkl7t1OnboDMhhO+wvu
sE6Qq5okS57imII6Zvhik/IQx3jaZ+dyV32TVxJRh6VO47v+R97FCkwvXsSpHvYC
oLzOmQxZ+RJbkzURpVAkT7E2LMJxBtuP39yy1RgpOPLjW4D+8CaDW6aILEMJwMem
t1ctRIgcyCA3Fz3fa1Tx/vpk7LdDQNfigNVla0WKBJAuLclYDYGeDuDtnz/7U8Tf
jmAnmaKrQFwBpyKRnTAx75FU3wxVz9SD1PoGKC7lZQP5/7964eCBJSB6+ML4I1hW
vUkpc0+VMvV3K+caHD3gDGyquWlV8qdUSX+51fkYHs2C894/Juua7WGAnFq5okgl
akxcXDakHOSjP2WDtNaEEYNYX4RTh8bLVKbS2FnTTlTrfuaoIOwX2FoWCu8Q7T9i
nTe+aTxuZxK9VAoLpQQvcnfbwUlOCVcwaqXTqBLq9wvKWMEGv35QUUW9Q30mwHAc
uCeVX0cuVrtSvqJl5su2Fg+J7QTWlBacsmwbPH0GVDvegyzYGrSDuSGEjT5t/YZa
C1SqsphFHdHGzGSVK//91aDi9q16SXplqmw+7LMKycjs/dVz+cLZfC9QyqOl6S+U
3/zO5RGDShE2dtYp6TC4wH3ftU6Xgz1e+og1CknA+q0GDAE8QppM/L+m2ynqPXfp
jjuq2b8hB9QGq6+BBU7NpBrWGxTCO8ZVMLR6v2WUKJ6BPw8IJoZ+TeeiysjfngmO
Di42tbySZl01TuI/1HA2+7LKW2xKi0WPRsQ+DzTHmX1/xUAlfSFtEqFA1qIo8FHI
7BR+qW2f3tEe2nqUXJWGPLHk46t0CAT63QwiUg2kySfxEE3mEhAWP82CiZ9N5oar
TGfXM3TirY0ol8AIPa1ejoVFtC1JAUiZdsuFG97P9obXAGYDg4Uv43xQiiXKZhdu
xkzZL9+gmI6PA8VtPvd8VIfgHQhXaS4pEKXr2UgAcPmU/29Gt69+W0rAo7yGRDB9
w5U7J2h+aha46SS+3kxbjwpVhGj0TA+Cm1zeE1+EBIUCG3dU1g1reSCF+r98Libr
`pragma protect end_protected
