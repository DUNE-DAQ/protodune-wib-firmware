// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DqI++NhErBKu+ol5LegHz94tq55xMwnxG8HYX8Int6iC7WCD9zYFvyhbXxmewDfs
uaTkpPpRwdvUp09bQpjnAYI4EhCx11L52sV7gHHw3vZlhBMnwoAGPmO9J9QvKpJ2
LNrjJCWiv6WJUzsspa0ltJGIxkLvu3pfPY5u0Td0v8E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 103472)
+SQO9GoxOaDjKwcP3eDN6OpL2RV8Churw1Ac3LTumHrqgZEtBDGkZgVRuco2MbWK
AFDzFfYSNjUTswwp+eSqvdlxETfxYVHFltg9O7Ce9zTf23bHnEXTirJ4p05Srzjk
JcLfUgdhy2LqO6XIEUOFpDC9thnhsqkfJdRXTFpVTAyvHQ3kb0lIu+/4V50M1hcm
pJRb1cA4C4Ui8CKHqHTZSDFsmu1uTLkB02me49yrvWQdL/jg2JprUGwPq761cpPt
MHhiMBEModfAJ+z74Lf36gpaI/MicnJk+PS8dbwkpNcOVbiEoKa05g//uIlQH8FM
2ONCXzVTWPzQ9yfteKwb+/Vszqatpig9yXTcmLErl2uyoKjPDbbsrWpiQOFzv5IF
jIk678vdBZNVhLNhNHxo15gtyugHyBcvx3j+f0Nx4H/slCJM1G1o224tben7/Njt
Bne17Ixkbs6OV2nRYi6QoyUbZsiV6tySiAY6Lt7iekNsKRw54jGQ6fIHxaCC5V8Z
+tsbPKfeTcAJ2HGjVnqD4+me4QYtC09rR3HEapJ35jDDBk5e61Zlplx5eqGpClU/
heV4houUkLol/yVWKlwFL5hh+0ltqUYut41gUFDMPdKgTXC6dIwJhDtKh0h/dvtC
URi9tKTnxiDIYhdOpYu/62bQp/q6IXnTRdz9EZ/yTtJHFTZX/m9PS2ZJI1zKTrCc
qKDr5Cgs0OPk3sxfNUBsKADC+ouvx9AumA0JxrzvMwRHloRUKLuUY0OywIALp7d2
+JkYnu5WdKwDklD/K+irY9n/YkWq3gYFAN1k88Br6zx7w2pZBPCCjGM/Os40XBsF
pdONwH/H4hSquZG6Dcz45VqPgrmRmNpUqXGwdQl/Ugmfd0oIjwekCYjYNVWuQmJq
GaaE1VeE/UM928gg8AXMO9aQZgtDqmGAE3hIUtRxVGJWnVDf674soa3/lihNQSX4
cZdtJrAghtASBGtPTQF6ncweM129YOrOnOxPiBpio4ZY7xJYXjuKiO4N6XJkvxEx
xlw+fr4d2qdiKp23JxGBdqnX5p9hZq1gP4Ajy2hVqy5jrGB0T7/S1d6GuW8P2akp
PEpIQXTyA3/FtPFDaZv7Nf7iN26gJ6CWqB9cTLaVoZz8ENuY41fjVFRh67b1swSt
IO3/6AKcwR41/bBSkCtjwOetaQA2ocJSLTYeq/o1k4PsHkOiMTbf1eczzTAjCKeT
3Poog6RG/im1/UjOV1O+KYUTR+YpJIyj63cNzJlIIrl9taJnC1P77kug7k2Rx27Q
fZfKogf6XrehzXbvx3buMIXqGnKs/PtNiBcldu/CpJ0kg0tLX0ILi3eLyu2aFX3p
Ghcr18426mqR+hwUWTdG2maSR1kyyPGRtEfLNVBVfrSjcWZ0KtkJeeWnKJUeh7ru
nZTDegomSmO3IHpO1J2Z3vuUI9jq3U8klbynbSgUuyN7jso0KcIIXRH+cbjeJfi9
SV5nOvKkrAF0nW2kxFHGAAbFE775kJjLJ19PxeE98bjI7B9oj3MEoM4+i7NijvK7
osQ92G2seU4JxqYf9gwiBh03RQWi+L6u0xv6InfTGkhfYhr30faWUrzJLhsEzd9/
ixqyJxSsoLGbhhsipibh//Z/M7mJIP1Guz8jHbYhRtnG3rlQsstV7buEx3xmz25o
3OZINMqkRNu6yT1kVpcCkrO1a7MrPeS2P63RBQCg+dY4sUZT5nWkMBki/98adnLz
aQwlYUToohF0nIyuCWM8LQIcRFq+ng4ICHqqBLwanqR8Ly2pVJJVdTBaA0j0SySv
mRmCFFWKnkz13yoR9fyRj4CXmMTH+DrILDQWHnDxY3RpgnvPcujX+3eBLzHgV/qP
eoAOVjIqJQaOd8FvaaeN/E5tiZ9b7224kmGll78TC5Q5vX/6hwUW/xAXl6CI8KaK
gdzVkErjdb8yNvDu9hWKh+aEBMHUcWodHalnfct3Lk58Q67EXtlC9+BdOtylllM9
WZ9ejDnJIDxrCwipEQj1yxz7BgxqE5ExmWONmt4l4O49pK6QTVutpCpHOKz63CNX
aEhkNZZ5x86tvDYVjBoRfeH4kp6Sd2us8noMdup7iQr11+LFMwLViUr65oA8ydI8
1ZIH7YaTlZguuqlKyMTlLjwKNh3h6bxatAuaeD3wwXqeL1wmnQGc4KLF3SczpeIi
biVv/IDpACR0uyfBaxJr4VlW+sDtME3atyZaZwHq6480S1qkHsn6v6Rr9PaXSSBs
3I9wbacKPr6jZVwWanSTk+5llzl6D7/mCIp8q6//r6haD+JnjzXvD6ivl5SF43Lo
t1ONBaKGaoi41Vf3SGWApLFydUCesC3Mfk0dJE39+fk+mwxS6T614eB85RDYnjYz
2Pu6he0HiBuZzX9QmmfJFzUEm/i0V+4vVznwf/4u8hV9XXtx06fU0dZ9UTuxp8Vg
Mqb/6V1Cl3F5+DDB9UoOFhH+M7zM6jCAbAokvglK2dGOa7XE+lwshetgxNmmo8UJ
cs2G3k9w2nrJUzdxowMwmzA87DFL89o8SMkZPQVsG/JOFwzx54TpNK50nfYhINS/
rEorpNwETswAG6r7zANncHE/RRGxfg5qd5gBnaexg10Rr0dHzqsJ7aUySgaq03Bo
gtJVfSKVMCrczXufttSXUguBRHhHNCfhyj25JdSsY9bRYiGJbNDlTtt/v/B/S/rj
uXyayCIVgBuVBUGawNF5ICoiPN0EgCmVEvOiBJr+3ETE2v6BdyX+0CJa+lXFG/ZW
NGQvdpLjmNB9iA5POblqfwn5dgrc9EvKPY+A4cmoc01wcHR+RvKjugmKC7DIw6fY
eVvYRG4oCedKutigTCUcuHTgxwrhP5fN+8rbcQ9LkzpUqe0tg00WvrM2FGs1t/v1
yF1TZGY6Qinz0ABVSgqYfgKH4lsiZcCyQMCM0Hlelt/3Rm+vJfCWxgQ3PgcpKaHz
4mEUbVIb2OrHCvTxZSozpD5gBUps+1NbKbcvH53TU38w5r33weW2GYt31/clh3kO
oOewluXYAhgCgl6L9xexpvDhMS5b6cRAZMA+kgoaTp0CbBywbu9brIXM7fggGyS/
5jTALB6mOjlNcKcTACqCsfuQyghEZYPTbxlieUH+s9tngdG+9NfaYI7uDYy4fDop
11iSKtAK2A27bz6NQ6rADD+uj+LBCtvxTTWieY7GJTzZfK6o7bjgs2n0Ps5ibawf
NRGriT3PE+fCeFO2g05aWQ5ntgefSviFfhPcIZYXVpCG8RYzpMJWzRl8YKkKkMj6
HPBjdDErYxsyopZxnwyNx7ggXtvbREhbtTDO8ktSmgduTphaJ8mnZIaq3bSoDiz8
a4u9/69fHd6OpZEbsCVhNC8lY8lAv4QGQSmnlz/x5CFoMOBLP1BjJrVLcOofGu9+
yXRXKu6dJGwHSWcr+L6aNlyCLh0j8R8i8nKcgp+LMvQkZqaquOLB7bPPMhCS8bWi
xQZhb45SbGnhs+AppJph//ffoAa1znXQcQDbhymmrS2Gg/LqzHdjWfJVEyTgZEXV
CH8rSuD1UBlfLkUC1YBQ0qZE7alT7bXkulS4eD92KALsOf38BTjudZMDC5WI2O6y
ZlaxPcWfxpXb4oFokDOU4d874JgLceEM3uMAZylLPhEfdFCRV+3KRAyZ6m0wyTjB
uJdkuQT6t+W54BUw/SYiFe1L41EHlt32tilLtU0ulzN/on/IbzONzyL72psv+FRg
1r9okRdjyIUaPCax0nuW3uBWlWFR5P9fHwh1KxsaOi5v/I0Ivwj5OodEwvJiAkBH
ZTylOEnr6U7htLcE2eM1IpdwWQ9Vk+c242lLC0L8oaZw+Jaj4IvfjcIimQ5P6W+C
B+hV7X37G/xqpcnzPNJuI7StCx7wUOPQyWb8XXwQBT2LlaophPMd8a5D4xgc5JUD
DjkA0EMnKu4DiR8TBcBuvAYXNzbAxXQJUYBglIMa1zU9xO4L/Wrz97Z49WlHkuVC
DWW0QLBr68qlgzf44e42gDg2mikaxfN/8lVPv3dqFHyLZzbYHUg+c42b4xoZpnQ1
jF02MYU4n6nP2SCltk/7TfkKJ2B4ReVrSFQG6lNdOdZHjQCVmM/58Z3+HVqvMZ5I
9PgLVuSpKIws9t4/i5dnHy5RbzJ/kRecivSNxXi9hizEof0Bk/HfWohU30BhxwfS
1AEN4XdIk6vbeFKc5RR43zDfCvMF3Gg3J6YejtvckaheFRECV4ZpU/rLj5o9KYvU
Zkk2lM7aoxaEJRys9j1vb0jdJN46LdOJBE8VyokXhlarmHeb/piw9+vwcG4K6wIc
o0EMRoTcESJtZfWA6TVFRfNc45lfwBl/XGCPh2h3leU9OMG0KLHXSK/y7KoEY5vj
M/GcpdIPP9/ahGvLIIupek41dGFt3avYEJaAl9FKphP16zYhgJ4qJn2qXqoFNVag
zRim6WRUPv7+jdPh45PZ3s90j6HCT64T9j4PVcDRRmm5mgXEGQOygnxRt0NSchFo
uWpmlCRwsLmURIwDIZ31r0ulgOdDbHkSB4fBN9DSE5iQ4XsxXnD03JIHpJrg0FDr
kq7e6VGmNBn6WTW0gF5f9tj14mmu1Un9HR3bNMARwlfrgcEPcVeMcH4pSwbo52Yy
Eiuv3sXI2wfOX6B5WiWmog3DLUoOn0CsmYrV8wJUbpmQxaHMmpHmRQ8A7s3IOjhr
ISTEJmu4PLPLwXxEUqhriRHxrl0c8Ewvft8GrEp0WytN2YQj0JBjpqPKf3MKQ3rk
7QGd5XkoPZJG8l/oOe1uSUfH+PdYDK7aNjtMqA5umDuAzME+ZE9DZNZZWpRPoqOq
o20K0vq1Us7iSc+lRFmQ0Equo9VRzr+ZgEeOpZFYoDH5Vr7DRDRxAP76FG/5k7Bj
gfDODBQUu3ZHi9cDGPXoB5Rg2wPc86e2rR+4TgFVDIhhaMFVuW62ixKuwXDlDc6l
QQEUngSQOtnzkeu1uUiayH3+5v0IRkolhWrjpeJeDKT5mSWJ9xUR+W6WQTztCe7n
zis9aAlqdeSTKp7oE6EtM6l2/dJyg/BM665XmX7nZePLdUquMC9IVzVh3gvQJH3e
k0mCicZtrbIVhklRmsT3OLqKRe5TAQ16awUxGByQw7w9jEsvZjxvCsWNM5IRoMkS
BGz9zmheGJviI7Q6mtUXMwMH271eGOz38SfR4sPKpDh8NW2ahHC12TFXWoeGRYPR
n7eB8JWjPsO5/0siPgk612uwvEb0UE3gFhKPDNTuIr9u5WgM4EB/bw6+Bh/5jL7h
xX3/cuvGLytVcDCE+2C1iLBbyrXp3OKfi+GTOTu8ie8aAETpkeZcWV/NvV7U+yqN
xovxGGcQ9gy/K9Y1GezJihxlpabkyI/iJxKRtHGgeGTQ3auAklthouNIEX7vQIR6
K0ETezMYbVikbBE/9mlDJ3Pi9TpGHAFXcc2g6xW4fCkpvQ7BkZQqzZQCLOlx/bqM
CyXP6oqtbfksoJcG0XgndID7FvO6/L3AE0zG1JB4GnSr/NN7AZMeM3LKRVCNdugo
mcnxG+bVpyUew3rWoksagwyzTwALZova2W4czCKR0tNGTgmhPfPVEaiaCfSXRTqe
lW6pKPtlYeOFVaxtBr4vw9Vm+psiTOj4QhuJfnBHIQsPSw1nzgYR8240S0Y0xwrJ
J/R2izW/3nUYTsuBUPeMzCgCXk3wHfElj+x2XUCQKQmB9ModfMSDvToi1kR5n7jT
LFF/WCkcfy5CC/CABJ6bF3CsmQc83fwH69A6yqxjOksMM7jZeU1MKF7bnPUKbTtO
UQnIg7ITHVKk9wUNYJhHd6iw8z7G5hAG7VEM3daP+PVhJdGBya6V1dOMx5G2NbMa
oUkF2pD69TQo4/CRkcXB+5SIAho4uVxjv61uA8FopCK6lXF8NoGJwOlweLaX9/yU
lqIE/0yx02PFpgGgiwTZyUyVawntoGEpWg8D1YgPKPckANsECP3I4V3MUKS9XTsk
Chc6UuSW3DCNxchidr/jEZXJo96A4BoWKPZjQseFDOEjHJnUncBYxpqxcV2H22Zd
eJ0Zuix0ENo3JvQurFfRLlXIj7awc7Sn/dh3PrpXviu3BW//UDrkCta8zGnK2UMg
tGlHBUCiPMfW7FzQrGpVCO8GV9ufCkkylFPq362v3dpoR8axJ/9/r6rOLGXghbCd
ZYt+7X9aF3sFPzklC7KtoMTMv/In0OzdDFmP9iS8oE5GRTfueMX5YpWgm5tuou0w
UdMR4TCua6oy157Y18K45a7fOX+Mi8wjICDWxWBr0/uLNhsEf7zPbQeCg60uf8Zp
8zx27A+dZlZCLQquW5/WFn0ydG5zYonnYyd+A9X8Yk84SClE4U7Vk2GE/YQeuTbZ
8r/Kzb4I/W07cyxnnw1kMI0qLcDWMRz3XEDzTbnpSYMxsBuAw4INDF3nb5dVB3f6
rSJ/tg71k0b4sbwaUK34L/IFHMdSdvwS6RHzUS4zCDLpS5BgLz2K4dm90qiO9gSP
Dlll3b2MHyGKey4JoTMgCXHqfyWatOL7OrXZENUMA+mDK+v4zDdo+SGr5ybvt1cc
+8cDpp+3ATY8bWSifq5nQE83VbzvLprhvWQPP7rx5DemN4/gQYfQ9F0ZHnJ4zF2T
Q+4LEYfi0cfZSImBJoz5ctxS87ZKoewgyQN5rB6o+OwfL1d9pVs0ixH5WneI1cP6
6XZun7nBp5O23JvGGkzK9PXYvjMXSHbxQSnAq1lr65kG9y1cQJygQTZwZKSzIn4X
vxmjjMPDzWvrrQWKomTLbNjsChUZdzVvIcTyNRfruY+ZODKXmJP1Fb346VjphC4I
MlgdjirFj2IdV5NSyMJRDZKHNqjhcZr3k6SGbF9ldVmjRi/FU++SkKi+VsD/hRmX
CGXPcfSNYss4VOSIPwsHDvym6mZC32NufiHVMOTu1KMP3i8pmpq6saJkvZcbphRM
jiZpKoF/3kCcYUWI+0K7Waxv13DUzOEZce715bHaayUMnBOi6pFVzIRiPoCFtTBi
fJuepm43n++GDOCvKmUKUkhLDjdbz7Y0SoSDwiXmv2GooTEZhdO1vcURUMZ6QVkY
9RUDhd+AI4rquuVJ7kCeLWxOtmlz8vzGRdbO1y+MkzJ8daqHcePy3N1XrbfsOfy2
GPMPLs6TKabZgixM5ueEX+Yx16AbIu8nvhTzd1IIGEm9u7GA6CX9U+v+9utLufK0
hRpJOkuG7o1SoafmdTuqd8iz6pe1GG7vjpV2giEVC8Ef84BMPgotC4BMlVQBsAzJ
+8bQeuEFq2PfXSwlQEOu9lpEsNmo2PXVbKwYYo99ZvgMj0mgc+bJBdGRPa7haU+A
dy/DqEaorCFXIeUyxMos0H7rs81rMkH1yEl0twrruXzj+e43mvoKkG8xNVd98aEC
Rp4LA8SZJBP8fd46NyltlRp62GzNXttWh4XnZFeS3+zNtyg9cf/WqvRpmxdt2rSD
oy+m/N2Uvdq6ezd226qOG8sYemSKgNWGoJWZugnjDTHRrnvbr62MqOW885nISgqM
SeDq4Cw1nux9BWeaoMJVGzJDVVWDSyzeoheSAHUp/npwR9UHiqZEI2PO9ulUHfng
VFhm9RS++LGCSauXMzbdU2YY1XtNkjo7b1hco3HWMuDrB12k1MPDbioXQFt8+Nm9
0URV7bBHh5CAsePW5TP//eH+ak5lpYPlWUA/vDvAnf+rHVTUYDXzyxhFRcRrFbwH
xE7Sj7HakjaUUcTCL5nMeZX3yVkrtpaev0nsYZQ/3zuPLej1Q5vr4VzHL3A06zJ5
BKxr6vnQosfuyd4AxDTfmniYfOV5LZHbboNPa0SLhMF/5JP7RMrDaVXjWX2/Dr1G
Z68xIE00xpsu64s8jIlkeSU1dz6hG7jLsKgJz+XkHF0VPNiZykFYITRyGU6iohcP
2bpDFoU4CryG2jrjXekr3+6BRR27Lt8UYYp5COpNmm5tjvzuH8b4k8m0UYmpekV4
f2Sj6ZleLdcT7v3cEQ22AlcaOg9EsZKpCYPlU+63t73+88SfMc018r+ia7RY7I2l
sEVchKY6uPY0jyZFl+MBZqUe0H4KwpeXmCuYaDzKCJRIoKMnRtPjxzjilMT18MiR
wJefEKmoOOHN/sIU5RAdxObMJcLSf8MtAQfZJhfR4oFbrS+eQluzdv6kZItGa6JT
ioKimp1whmkd27GtodW/MwQcaYH8Fd7UV6ynrw3GUsd2BiIgHEfGLE0svr7yZ+1r
18HeEwTcoSJLvYKzHAidxwF2qxSZW5ZF2S1T6Ev6LDkkFqx3qbeZ2N5MJiHSCV5J
wbQQu9AzIDfrqX2MgBCcbq7ECRUrTmIOFWBt1kEZ/MHinJTp+XMYjG5Gum787VDA
ZqiSrXw/yF8FsG36jj2R38+RQIvnJEL9M83FuM+o6iqe3oU8COFyZWxlY8hUgvt/
u+bgOCU7atv2cKNzzL3I2Mu4o7PIkDMC9gkJNOa766SNyFYbJvtRqHYDsYJoFHuV
5epj0yI/Oh5l3j+eocw+gUGF8FM57NOmPAw3RiAY+khkkRYycHL2s3Og9efqJm31
LQGbKIOwdEFXpPcqL5fShKEJ0rTydfApx9YW4hayfD2kYcU0jKBJXqmqiVXJX8Ai
l2q+Saj0x7HljlvjdhyD9/9u8M4TdtLBWPnLAU2Fa2Z9Te2sHnZC1DpuiBfdWcGu
6TPHVpYh7Mpkeb5UyOZE+qjvGe+9wZq8TED3EnkD6Xw9orIkOQefPgPpBD+ANYW7
nDNNPYmNRPkEEMuN6lS46Pjv12tWQfXFaBxwcHMb6xnKBNCyODewaUfsfBY78q6m
MOR3BExDfcul34RaXbToqOz7hfNB/aN5GmJuCa0q3Yx/FQyL58GppbdYypaqK4GZ
YNNlN8WaZD56S7e/XJ90ikdP1yw6KoEdMRfxlo/Pt3kYgU+eNML7OaJikPfqZbZH
nNuHFE7Nd/q+JKHNUnnTr0NMHwEANV7e9gPbnPv29KH4u2vaUIUgyUfEY0Xa6ZrM
onckYZnReLW+AykGI8Z7zUFO3/J60/uVteV95MBH6E6u7mSwT093HH+sxD8JkNSb
0gDhx1oQP/2+TGf22MZnYGUYnFwA8dkF7ZZLOm5U7Cz3HqeryvlVAVdOI5eJWc5g
0mjgDSpl/EUzYayJPXFuItTj3WXYNAX8cMFhKBl9A0IUuN0oYyg5Ka3sUYjAOBcs
UuUg6p2sz3kt8vUjgn2flC779xLV6CrKCocRNeeOzusK7DDFE9Gg2jQh5ZnVygd3
5+XsXqHYX+jTjq+9pdMmvMKMShWjhcNBtM4Waz34Mb43HaWiOrJ8SfCb+ZX3I2Ap
irtO+J6vvx8uKT5w5k/PNUtW4gaUO39DC174IBt6P/MBC8m1QTqBorK2wSrivZNE
OSjMAS5v41FR3MOLJCFPf7I9gE30IZt+ua/S7lGWfNCsCIEuapT2aPlxYEv8JeNO
b91TrhoRBGINrrB3E+EnmHEiY2HqiYdhxfA2lF+Z8f7iQUIqqcwcPwKcy9q5AWdw
ovcijBOtEkYFLDFfjx1foVZO3QxBBG2XOrtitjKbXibrl7dScPZCVux7RDxkHF8S
uA+apsFKlyN6lzAIJo6eAw7mGGlaXYsnPlQczMk9dSGQfo29N0QaSAfl+EHL6p6r
6R2Eh/whkNYauBXmSZlqIFiY7zL/YcvRyz9JIBW0Fc16T1aBVl2ykNeTdvjmYnhJ
zRIWvQi9hWRcTu6dputGkLzEur5q+e1r60H49csgo0xq9G3zqKhZeJPWufHYo4xx
74Ryr9WKUvtDS1XDwQNTnzg45TID9YG/D7yvjU64gHmBEoHk9/URMYbDJ121cwZV
JUjCgi5OrZJeC5uKQA1cy+U3tx5nPFOehfGgyHXc7vdbr3kxmR4L2W1M3cN0kOKB
yg96ZDCdLPZY5RTeAPct38cSAIVTSW400HX7kU8iyvL/4uthjxpIAR5WFHq8XVeP
0N8KpmHl9JgbaYT5nvhNyPTbfpVGJjZX/EIVjPItS5E1EBsd1ez8y9y/vb1H5TrU
s60oR/SJJzcfrpXZRBM1RsF1ponnWCqUUNdIWfhFdpIemj7cuKOC0E3xuOn670Fs
dDCQH2kT3BmZJCcxypulMmq7s9nZEyxxJyPmNbvx/f8nizSSpQsj0WvKXtoaIFQA
gUN8A1wyn0D3pin6E2QvlejBqYb4gxS/ooFXjUIFBLl7jKtlscVSm9As6FiUet+2
iJIMz2A0Abum2lesIVBaHbnUAz4eyKb4pKgM7Tqpd7zRGj4wfnjX1rqlGyDB8jlR
rb13nigtHmHCzLtvF15TPnqf9s0jeQmKaGzjHKmKyMhULvvwHA7l7/GnMcQImluG
9EQCFNO1ukEg4mCSmqFvkXr1Z2pgXB0E+nNuAGO6bReoeU/xF/Ua0iSI+qHvIrgw
U1jAGeMiYbjqj9NUeEQS7rmfCFE2R5NEmSrgDD10QxtJ7qQiXugAVZ01YNqw2s9a
NqKvTYfoAvrppdVga7IpsWtmbpHebk3UqYZKd+Ew+2+Yub1ai6S7JnJ8FMPp5HlL
BIEB4Wga/3fVQBw7BSSTOqktJzB4K/8rW827EvN4ep9Pu54n5gc7gujdsNzvL9n7
V417FmK7L9HufgFhe652kVpaSZu3ePY8ctQJZ4eiANFpwpu3l8XpfsNsvvFZBl4q
LD+/CIdTr3WEfnHGPEqWOU714H6g6e8/u/SHggBOXbRg6npzjpQiR859nSGe1C++
R/rp9z0bMMxIEyjwzzUPttoeLVH2jAaYhex9QZNxrJzzxMnFZepn9oL0Yg0eWNzv
Q3UdHTpo1lhQDSUlnh3TmIy6xurRrMyGxDBepJgLGq4EqC+H+W9cQ9BvyGpNR4aX
Z8VHbzhuX9ntwIcqxArME9n6WZ78htarcki6QOvLu5txwNvlHLk0Vbs1kkwujxNo
KFqy/o9fnzNBWeDKLx2ObbxzcyKipVXMG3oFKkJ6GWZDdu87wG95vVV2OuinsxOT
gjs8PlJcfN+IlEsNnrgzJ20LLaKN0SgnUKyh2IFmj0JNXI4gdNqazYEo0qqTlX/n
ocMH9DCPuYVOyWjjabWieYakWVSQVaNBZiYY7QK6RGb0wXFmwNrlM6WyeKzNzY7N
I89hGbkWKPZ831Eu3SlvTGQzFcytNkg9P4gUsqqs2kscP1kbGMNCiwXxPfgdS1sp
rVo76ZiMdzpRxRDNLI6YjuAn/MBanX4Zt8NPOrZyGg6+tnA4lZ1ESIzIrfPdKY+r
RMVjQYHmnisxV71ZuDPM9Kkpkq/zcZF4760j1EtR798hkl+S9Qza4/4D+BCyEzYB
pO7trovPS2fSfkmqX1oLauXUaE0RuuUzHUUUVXcYrGqq+5r14tauh/rWEdaEwfxT
TCBcrAhPABXKaDOlYcPb277LP22kKCzs9x3n42bf/ozN9LCoV5x6T05Vka0u9LW0
p6PZmhsRc2Lwo4RNMd28+YdxodwFzmWr/2eZDLVqXuZGZ25WMYYWFB4KeCeP60G+
lvtcO9/KMf/jylwp8OjpDO+SP90O4sJjTXDJaqFqN4pJLHFfRDpOa3kgtAZSZ/dz
EXXRMg6p95vN8BrBaBhvJzEMCLr+YINcpp4bjqdjUtcJ09wjNekydw1j0DEQ2eOQ
di7mJuTnbRBNhc1KwH2lwJ5QRS0iGq7/4k2kXMgeYrJnqAMhmrMiN7L5SSXpIfVw
eGFFTdNGRxD8o/ywSvC6h47Nv8sfjYoZhaHTsWynEQaRoAeNDHrl/soR/dHN/tRR
+inlLRcQ/ZZBU+1r5cfTU51qtfBKo0vb5E8e7u5tyDW978NlawxRXJXe44Tt3OWh
KoJidylCDbwus/WkASkz3xsEmxP0NczW+Pkl9459BjOwN+kImP8mpaBV/3H2wt2C
sY8WDwhuL9JaEDO3do7Yebnjz0OsY0qCMjd6d0lGVWZc0YwEliBRqmNsL1tS75wL
FQ/xrf37UntfNuR3m6x6jDwk98UsphKsfJlLtMQ9o1lwkQ3PzdMv8o+e4c7MIhlj
YoParxMPVi0xHMHM1FhTJtzk6lo4hS+SG9YfuCeQtZVVKKFNbF0nYNJFiF5xA8tN
qNXrS2Bar5ksFmxG7M5Pq2Wqq8dhmHmjF27xluqKmkKzHp2LLVeM5Md6EBjVjs7H
MbDZu88/AiKKk3uuCntU7LFRqZy8ENWbQ5NWchT4omwZwALR2bMQ9H6ZBwY1db9X
acZanx/v7r678Fm0c6OWfBpRrAHqRU+3DAFgpIUt10nrChxfFlyOt8X0HHJFStyK
6/n4bOezcqIa90cKE+7iEVxUIuFVt+fiH44g3yZCTVaoD8qQFaI6O84xH/ZDJHhT
Ux3gBVtHA3HnkhLVIyrMcy+WMFO9xQv4BG7E2Kd/ALAOJvgkxL1wLG+LIfa50uRu
bgTaxt/v9uul1kQ/fuK5nU9B9grcUG8SGJyl0jcIcB6nkbYf2Pg5BtYx1vcFqjDL
jSvoUqzcLvjwllzSVgItXHGtOa69ZY4Ddn0UenXQSUpYSht5e1XR0Lm/RbYGWRZL
uApxuVfnBbn79ZvBa4PVvMT64TbdG5EMVq4xqrDHufbHiko3rDdfvuzf9WDr5mLd
UvXcxVaTdQiwhxeodVX32xepuysbhM2n6zmxUbmyC7MXvmAYSGn5Ny1jp4hOK4dW
Nau3LdrV4INtskJOtacu77rCIxSCEwzwu8bt+Qmnj9bsw90mv/4uZa4EcJDnO1ud
/RfJziE46siZccP9v8gTbHXIgltNsT5nSaJpJ7j8bzb3eMrdkmiKl6oHsxWOKVKX
5x86IvWPh2AmsGMgfSnein9I8nrYD5RaX6zK4zh3wIyJAbM3ZCvcuPRgXSYomEbc
hpkQB5NJXoZEwUkt220BkjEBLoXMQlt0JCaMTsgT4omrdAvTjkyRNZrg3Xvqfq9X
2rvI6W08lrsXTfJjiXE7mafHl27XU+0cxYc/C8fcBK8iRZgqcrI1EHxjAJqDP48H
IGKQ9rWglNF55N0ccLSU0D0jJg8SV/65b0/jx4qzqKML2+qhKadhoxwdUWL91JwS
RLOLloML+YDmxoq6Ek74+1mIOznNwNZFllGcue3dHOaA6XP7kHG/fFxSudzeHt7Q
baBjGDqVNWySWw/8jZHpycIqidjubx13G5aUx9OnAnYFoatklGlxhk99pdXPQsV5
LoZXgjxAhXji8kB4EJllN/caZOEsJ4hLEbc8oRSMglPIeqUxQwBIHwSbRw7/ZT1m
kMxsoEKWqKHmjL7svnUfyQUWmfmb5fAmt4iqD5zAy38CZex0Q5bkCiLlK+gdhPV2
WQH6xtDsdnEBxtwWgAsZjCHvT+L/6RaVrbDeVhSM7qqpaLurZjrL2wzKeTDd+KEP
P++BVRFCSJ2wvOUn3NFIAtZPHiO0EWufCanp+ccRkAoriQrrQ4lH2gzWuh8XBFna
HdXB6jTVmDhaIRVjv9f1sc/HcuKs7UWGswQM1hxRAz0aIy5745ohJ7OrVP+qHur8
abG22PijhTO7/Nr5oyXh5fEiGpmnZmxQYmIi38cq6XnvC6QHj6dVoyR7xAOxJY6Z
aC82ZAzBHsx3/U5csJzTbb4OWyLWJ0IWdCBLPKM1sgRhjoGrJrsk6i+fF4NTdRbX
zRxdDWLzjvqCy1UUhfkR6po9zUesjmtr041bS+rhmnb1YZXV83Rs/iTbTibQPxid
EcX6wtU/3w8aT5NgwEj3AFcJekm2R6zObYospXBmp7ApzUqGo0jHM4eXoluD1tH+
WhOUsmjwdU68KVQIJKUyH5CvEkLtJkhIM4DU1s6qCGtxZ/kKhy7cfVgzIV39y9fV
KSJyIxWq74U3y2R53COGm2mhTZaejvYD1B8g4/Pk4Ggz54+EW4rzIaPudJwfQros
EheVloV8eVpWiCVYUSTa9fp6A6/JG5VA3ejzb4bE2jMFN+/3GooSYLqcAXqz3i7T
WVeHIr/wVBivGhjVvlj1Hkmuj7bdaAjwPMTobLoSXWb3F4euUYq3HzRV2qh4UeFt
fpQoE5H9za9/EUN9WCbk4liOXJzjQg4zVeq4B27YlOcRGLzet9f5WcU2NTiV3s+a
e/ElIky88x/f5wzIbwq6Iplo/rkkLf+cCX1WkCJPoYd9gWsMIqEqsicCgPBjYvr4
/WUyTUV02UWHID8joy3M5k/rb2Sa0mUOzi5SJpeUtGg34P5BCL1YcUljz9icdJVK
F05aFds6col+R847TAb6y3Bnhp8NpcaHpGNww66Z2vQCcWPgwi50Euu0wUFfz3P9
VUJ2fuzNCe7hv4ChyJOC8WElz+JyS7tMLuQSBqIFNTsro0tbaM6K4GLmudx3idSD
MJuuFS8WpiWZWjadcvYRxA2lqZbBersSurWSGo03s4alRFITnzk2K90Al+BMxMxs
xHIddHyThE9Gw2KsdO7vg6V70DwF2OSM9EV/oFlfpQjP7VFZ2DNzCwnx2QCqFyDU
J9LSIzyQw61hPN+R0UcHiHZbKuggOKde3TBBrOx2RqQiGJK6oEpDhlmFcOkVnaxn
3PKXQW9usnazXhoJZe75XePcYDD+SMNfXs6En2L6NqgYa0GLf6rPY4zcXFVdfjmA
gQ2rwlCr0mIoIqOEx2tkRivml3fE0umzQl7E0ALAc8Jg0HN5syEkiHSWKX8A/1zF
E99AasKdANV4RpvF2lDsV0pj8C5sZ8Ws5wvS1X4fnkuzou1TBnqhAs3brF3QQ11M
4tS04S+Hn7VrAtfshMkCZquzO3kvHlVrTzHR2fSMIGkbzfH66xF2Xhd9n43X1vhl
7Ku8CGOpHOY6muCQsh445XwKHHwL6W+z6+8rfWvQV2uZuCqkQ+y0XuVB93+EbBy0
6ldLryBYTw+vT4k6ID9lgqjot60szai0VzIOZVtEn7DudBhY6GEQiMkSyrICqo04
bEsr7jVugspi2dT7SKYvaGXFCw0XwPgZL+hDRRvwvuUFK+NYWZ4b/L2oePWB/dq5
MBIG5JQULL9i0joC+p4aACkfFsjkVeR/l45yLdJRKHt6mwU6S9H9N3J8JGFJR8f9
4IDKkGmB4FAtnIaxwC8fOCbug1DGJA7f8NN53qoCKvVezpquW7zMJZyeU1ectvg1
7SrzFOBkUcjP3LZfUaeLHpGfwXRbRrmx5O/AvoaBg5STmgBoQNTDDLZAnPwycZFA
wgSJKyqzXJBI4yyVO6MvDKF326kF1GZma8ZP3b3hdPgEtvFXFZc89Ksxzkazz+VN
6di2sh6r2WHL6OUfShbwga3xlBHsnZy+Ky21wEEQS8X/bNknl7RLyxn5YrYnT6mK
FxHHYLTeAvBl3Zuo90yhrnIaCnsN3YJ0yOODuANn7abQSHUbGmeCqYt1RQoqoK0a
jrIo4AFcbgYh7YkfdTLM1CLcQXjBHE+gFw1jkwTRY5hUVNsKU1qHmman+0vJbNdv
yCIBsup+fL1JEuBErWsw/456CRz7Ah9yP4dUwbArIOCdPhUlw17UOlEAJ3Y52+DL
FDJ+VOvL8MhSF4cSGjZ1Pd7DtJ/uLOJltpgm+dQKH8ir41z8EKQO4zbuj6boNiWt
WhE9ujIk+BRFRtcVVWHCh7QM0C66trt1Vcd4XZOJM4aPEVCUTG0M2v6MOpZ/VWhL
+bHKlxa78IwQN2IELOMOQ1fP2VAOOzKhrXm3U5d5yw0X8PmBXZlPvdb1IFxWgHCH
+/uuiXiCPiwZ8EMAsUFVVr0hwobfDgDnAB0uxxQOuAht9UZBtPb1W3ldNl70UyK7
xycAMBfCB+PUW+ZmlrKROKvnZ7fuh2IcTelv9SV2pSStBdzR3Dsv2UhwvvbUHXFc
r6Yho/a3eM2JvNWaxbGDTwqzu4UAFom2oMt6qk19pCjldAhJuHKHMK3/G7IezaHS
uaGmwz3O5XPHFh7TlvJWKoHO9uLmhIXJaDsz+dSoGXHLYxPx05jQP8R5IRGvNX4z
rkSf870N9BYAL5kElNphw+9dw+VZRAE9i4QYxbsF/Cuyogh6/VXDx8LHPYYC0ZRS
tIgZ04yUMcxMnnVCEOaBkNkSzouPx/QGEaFRL4TGuuwryyCLkAHbt63usuUpYzRx
+FPEsvnlkYB26JyNaCh7hKhPL8Y9UvardDAdZ+EauaDUQMO5Ks1tEWLO0JwpDGvh
ehBrxQpcWM4swBvYg+XhyXMYHDejVKkCi1S768l4t1hvzmsDieG4O5jGWRe8CU25
KnMylFkRIRWucTQOnSFl6wZWez2rA/zT74Jv7qbt4kotSA7X3uvTh/FX/0zBOInh
Z7EdoWWKRlcdGGHvbYsMEKH3pUQWxhyZOdq43DqH4r8D7y9LNl8GIE2b3ySlvp1V
Bisb+t99IVEHBBqVOUc6PudDG5GWd7pqiZDVR9crZOtxLKrwtSFea8rlpaJMxNQY
rNhK7qhGhkvbrNwMFuBKqUBI36e7KdAEvonBQkfkBC5VkNeUPcI760w1io6ZykEZ
ARiEaNFBFRjxKH8Wt97WzGxE+7HtvlebA+4Fy7+QVw3t9678rDfABlCqe6uNs5u5
O+WiTuVDV+Nvkszcwn/3sUjMvQh6Jb/hZtGppJaJLdtkpGxpFPZPZs6FailAusSE
0fZ3rrgcuxcaiLHb6o9KPUolqVSwvtwhaCU36mmaU+JPFYcc45n5q+U2Mdx/WPJu
J8qWD3k8lLsIgrBKQEd+RIekrn+54jLnMhoPTijrqSycvIhiiZtVBNYqrJuAzA3S
wGjBABc05+zYEuaxjg8gO1hRVgcnLhIv+5/dwWpY5JXJo/P9y1181QmJbCSNBkJd
GPbI/WebvMkUoMrLA7i8OvKTGTZ4iwYEF2r3fcXu0Xv6nrGdlpNlaQW9pYh4PJAD
CAEmBTbvl8xoTVhveJmpqyYKvyW5vDDbJuwlHZjRIe2K+zqlELyx8nB9oFo9kfWt
yxTcKL9XvY5uvyyC7OnhubQ8/7/A/yNllATx71dGR7gyS2yoHx94WH4XUACt66MO
Q+Sp65bEmUwuV+Sucro1n75GHRGWD4BSUXApXdEfN9G3B/z0NrIVUkfJ2Ssodb3G
tJ4yyd/R5HUYQgFG4vYRBFPMsuZkwiZGi2Qa9dXxpn1a/SrrpF52uKk6103OY2ws
qVhpFNU4A5wY1n47byCJJtdHGRc/ouWQ4tjyfeabaMFhO/G2Ly1UoK1asI38oxEO
CjJsNgHD1OxbJtWFa9G1rh0Khbwe9bmPdXS7NybtKkRHJSSk1ewnaw4LC9t9w8Me
YyfH6kW+DXAzrukKqX3qbLKtZqe3DjCOaV4W0w5cdd5nS2s0v7pBdJVAIBe66awb
RNOe7GcE+JvOQ4aqqkIMmzrDUsaZpjrnQ22K0sc2z8aYn9bVdoseqzfefUk3Rpi6
XdQ6MVFEpWU6nXAD5jSqw58a+2afQUEURDlZB7GX3xAEOIX6kR9JCn/2G13geCB/
FGZ6y0eREBTMOjhupaf9UacmTYZvGT7CugVRxZlyLl5MxaGe+5dB/SDrqp4Mhqdu
Oo9nQmGXHVs5xg03rwPXOPNheNGUnRHGyQWfJF+x0okOv+rsExKlCVbdZCPvp7p4
wYXQ6Yabz0sW99Ew+izHiOwNE8BIAgzvW6Cvs4E8v5AynaVHGFpRZGJUfPM/oCp9
unEh278LkyvIlZYlgI2F8D92PgKmSxthDrkdNQ65Q1ZrxnhDSRPKH0d83He7NuXE
sqOiTNfCrvcVYvlfeKrfbQoWwMb9p+h/WM89TGrkEVTy2TZVJZQTxE6XkQoqOMZB
3WUv434hrmb8rX4zBCgt1sNP0pFQbMf6ordL+XIvSQVYueE7W4lc3paa7S0wwKjD
L1HUaopdcjDQ7f2/abo2JW2jw+8Puj8i8+clskmco5TL7fvNDvweAD3jP3t9PiaY
eL2BMGRn95FBXuWNeB7JO1Tf13Vqaq3pGsSGav/j/LKQKj1dYTEFY3RxqVSKvCED
U76cPjT7UwaGyYA3LwV+AXffk0kjh5CZpBp9kJ8YpUn/sglKdwx8Plf23jCJGKPC
TRDPPBvHrN84riiEipWH/47p6fdWRzm1a8S3B5Mh4+GellmI+sllnnHJe3D2oY30
Qy7mg6BmBD9vMa1RRILVk9BKS3WsF7FoqedGcrKvhqBYzPPKvteb9DiOwo8hYq3A
fulaMNNAabWW9QMsQsTs1eLYA9zIyrPFiHUvG98JmD5t8WVgCMe8LnOVfVY5Batx
3RWzBMNSqlz7+iV72xP+Uhvv8vJgR7QAZdLMNi5CVOTlIQYl/Pqh5MBJTRtqoE+Q
1p8JLF2TvWrKeMv3d5GSh9fBJdtu1oJ3bvuqvAUwlDafD5RJiHCxs8NP8KSqeTxU
ZVEEyIe8ouLkyCyOO9Wqf7KS9xmdg3/566vRCTpuOhNNBEltfoU4nXPNhvW+gIGm
IlA6AXMxMjZcwhm66ZQTFUtdMN1WDZIMQoSl3VF5pApYQhEAJ7Bkkpb0mitv+7KE
fnAG2MMcDZi8ABRQhyyacTtf61U5jE1bN0mRE/1ruTzWILAqKwaLwY2XMF55RLc2
/DXxAat9nNFsETbTEukWXkvZjfreNwfBrER/G/tEL7koa3g3PlZMIql9m2d3nQq/
+uxaahApmW/MLljJ6h+BqwuVa/ucpnnqGJy69GUfUq0gmrp+fp7mLjBHJdEjLDnu
s3zFN+G8/MOoL4tGY0FeUdYiEQCUTWke0Crmxc4M7UBSA16Gz0E4TE4Ld+2kL2gt
+lZK6lbIq4M5N1u1nQ8JYY92sMVFWLW9cu9/STUYFSLj38Q/HI8jLpwiEU7iKvvP
5EuG5I5EkNp1D4PC/DxiGIsRk1TDkXpio1tsnExwpXzRHCiW+kyzU+OFFcl3V6O1
+0P7VlA0//C7p4RsPi/juWWGbIRnwvvcWCg9HmwlHwaZtTi9rsb7qSxtmKgvoFdk
MWS16V0vCGOx+YxqaCBD3SeC5FCQH0lr+3bGqI/dEsE1ExG5GKO46J0sY33h785v
DYCWUhjf5ZWg6xs5kEtJwsjuxYZDuxYLS1/oWU0LuiH1obtG3pew6qAmTVfDODw3
aq+WzMy+bto2k8/r+X7QpYGUodYXxNo+aWznDuyH9i9Bbr26+KT4R+l7nqfPqDWT
fu159gERmC5AaFWlBK7y3L6ms0emDvl69cwwczfeN4e8LGZckzTnFlNMns1QXP7N
hbxPwZTbN9jDCnavCs6iMCV1Nn4VrfhPfZwbdvLmd1P5BbnkVaP9vZRVcYVyTqY4
7sPSikcrpRoVKRXFnDgppTwIFDkrLjQoz1Vx9ImhvZA5g3mO0hXM87J1L1gqLlwS
R11iLFg4iTUcjcMsjtnNdQFn5go78T5CuOEN3kZpiJqjicg8QoMsys7smwPpiyU2
3gjpxaSY7dTnxZfUOk3kJW8srQRNQcQNZ+QANlQ2LNX3tiw/eZRBkXZLG+cekxHf
tZl92kAOvU6FckAQWNHhuZf6y+oPdFp8ClGv9gr/ZTDilUIGk4FLsBdbC1zoVIbM
HA68Sj3O6qu1leRSmXEwJwLrM309XAyRqmubk/jMfXLUQyWVInVH67BDapStFJOC
hkyg4o8B/WLZKXvqES24qAKrBzwZ8v0jv7F1rHjKGXWMmY6pBTwQzqdUVsYmdsZn
WgGLrISbHo/4HmICCu0FZnWehqI9SCTrvoktk9efdu1fx8+XDDFMpbZ0lLiw6R4y
fWO63XJk2boC03CI/6ejRvkf1gFSrD6DMtfQf88HfaAcPwxXYorOAqOPfPgpZd79
W1qVt/jYsg+Q+G1gJnUdvDaKD1H7/Su4keLhDiHxSu5W/mkb2Cs55j5TPkIftZUb
kcDyW01VMSY9wwwVOi40ANhk5H4EJfMansRGSf5M5Ky5dRj4/Gqzi3Eq7C8JN7NQ
AjZO8j6FQxWi5Mm/peuLq2rDzh114CSSOd3ah4QoTNBWkf4Ue9QG2IWqj5rtLveg
F1pjtDBGTIZkqu+qk+BTPnCEUABxsQ5aEuLVRXoTmHbhucQmhqStcoNy4a7H0G2G
ysk2H6ncC/mLJjGIgT/mOz6xFBESJyh2P5kv/JYl8M1zPXopPjjl25LwAyt1NPy/
IITLO1oJqo9rW3d+nBDiBDMQgcG93zp4uW73tHZoSfh7sNOCVg49bdx4Zpgixd8a
YmvxyPEeC1KE3Es78MrPI1vpMPtdJwNhwpJKfEXg7Sjrwhx3xnCZwNtIBP6qSSVm
LymB0BA9SyQV4oQQglIFDBDJrZzPUmE7Sc7SSUFT0WdbQSMmUyU0mPkkWyR6hAop
f0ZjfHbtuBx83IjLMP2MZLQADppkg1q/yj2LJSAEINxZT51trdMUXNSOz3ImsoZp
rcGrD7XErw9ESXBvt0ZWcHs5HjWMAYA2wWoR5x9ziBQRs0qvy6P1Y1NU7jcL2H+m
zKlnI9/uGPdBHwdz/d+H64VjH+vPlwSc67Y83CtdNCtevDK5CDc+maQf1U6cpEOd
tvR3Ljp0CYJe7/fD3lrEYWc3RLoJSnj+oQ7slgGJ9g/9OqeqeokHPF3KtHwaFh8T
AZeWGlegoMaMa76EnpigUa3Vc32cEEW9gVflMOcWmvtmZBg3KyXmvNHPgO4a1G6J
A4T3WcFfFqgPEknSbxOX5vXnKqpx9WmzwQ8Inj4ERT3BZbAMYuVG1BpQZT1QztC7
ZAzgqwEqSU3J7TmrUECny9wAOdyg+Rt9TWDWgm1j32pPOJNz8KQmYEd5/M1uSyEs
3KrlumQTxjDy/BPWfnu5qH4AhO6Ptrf2qhYPd5ijQJZ6xFJ4ga9ijDVhqGRZr5B8
B/woJ2BoYoilESIEs8RcUpCjtizwCgsisXqckuf2lNz9cDL2IjmmY2OqwCnxiKRI
FJDjP1ECoMGBaG/6VeuXEDXuwdK3sfwP376tlUpOsLGgvbbGguEOLmCGVRMVLgHn
EIWky9ffiuynAcT5Rc2XcmN+okLvje74bJtdiHc+MBIxj/IMRras2eMaaSdMCgAB
LFb38jTxovet2H8BE6qHkQ/Z8f3OdmKcKEBkt06311GBXnfwOUJOsVUYJ/0buGPm
JkXVkN9t0NR9ASR9iofc3QMCHEz85xzwhD+SWAYCvrMwgibHA+e3vRvI1sF7kEXm
rocLuF2qeapR2VyOJcA0Hqf37ar8eamTwJUzEukZ0i++w8nLpxYPl3Py3pZFtXZ2
6vqbenUkmNmhz9WVQ3RbddrA1mqb/+KD8I3A61KR2KAW/Dkcbe8+lLyeQKtFsLgW
jSSqSDCPW+KpS9CGUj70NfpIVqqMB8HNplpzePDcLo15RgoZLeJbLOrnvv3aodPh
tofHfrMo7XC5pmOaXEU3mNi1nAZvFADf1z3TM+OLAxf+lwv/P7beIhUKBMgHgwu3
+7/LBwsqnJsNou7cUd4I1oHw36Yo5hwxyb3lfn3IrNjrj85DjDXNfj992JOv0al6
If66xajUToHKhGZzKycuoF2prPVfHoKzPYkTiluUOKZaJcNi1+u+poBKWlq92MYq
tdVFLKjUOl2Ve1ORBiZMOVTcZYlSA1RBCpIfPw/d2fjihZ2CX5XsomOpN1BKlp2M
GmQ31eeCfvPtoPYDndHJsNu+nsq524WdlBhGamOTWw1CjiHVaGN5RkLLHIEIKUfO
fzRX/xM7XBs3r4WlQqETsI996qLrOKM84KIZcgW1o40m9cZP7kS+R+BYnRKowxM7
F71velEpwP6LBM6ue9svXTYQrk1zDcswXiRrAW5sXGPQX0n57LP10LxGlwNaXSwK
3+Q9GJNv9pHd8/NQG43TCX0pdi/o1ZlXm7c+xlrUggdutlIhwP8FFmKTRxy5qMV8
75H5HcfBewH1yTJ4PBEb5czGvxUO35J1HfyJ56T8+4c0NT7Vrd3+0uBhU92hK0wQ
60ScUs0SIKuaVxS9oZKudwcqOxNWUmvKgUS6kP2ppQEIky/8B2G0q/jkluwlkwpJ
Dy9h7pDrChBIs5jtK/kW4f/KsHzDtvlLmUVr6i9Eir8v3kLC8tocJZ+ma0mi6Jv+
aBAHIKFaq5OjkOLzlqk7//lA3AzA/o6F00zujJLT5b6sTDSHqFeL16WiHLCIe929
AdWNT7NOu4CtY5jB1P/KBrjcI+62h8+EXdB7W8/ICA9S54RSGezrIYdkKuuseHja
Y2C+FjlZ3bSWNWzMf8MBnqOheGQynTxDiNKYuhCJ12XG0AZnm0B4dbh4/Wk8uk+Y
+PLmU2cL4HAIWBUV7r7ugwrixJEAPtGsD46z5a55aOPErfz22bLZ1dgJ8xMqOh49
g2xzcDFZ2hTHGd3TWRQOhBov1111ZLrwdfwqx1kpNadrL1iNj9GZJKHbK5n4Z4nL
eWh1SGvZqrEuckACoaJvPmEOMj4yeqihsGHPZUmmLIyC52L3cc+6AqMAYU2iM/7m
JmTF3xiQrlYwx8qIdbB4SXybPFddAMijgtvzp+EKYdZLDZOALM4GB0U3aDyi/3Pz
Dna4+i7KsnRONuaRROsgULdyYpyUZjp2WcppAlrHcYeN0IGdShIX0CH0GTt8C5su
Ri4nSjl3jxxY0b5mNfFjJmTHNRObqNQH1W/uHVyi/f2bAdiyQcIMzksQ55nBvx+l
vPLr4kXlkjM0t/L6z0kUyAOta+xY0ND6fgMPoMPe8J15Nax19zzP/ojC8LRJ8eHs
iHChgvNeki1uGnx8gAH5tgjm7B+RoZN2iV1MnjFyPJVQjiUqxbXfLFVAozUH8gJC
6DI+xjCU2Q+wFh0X5UxYyTLlNRs5L6xFaPegie3IDXgwKAU0U1lRlo+6SUC2zt7d
GmJ3RKFqBOrzMMCozeVNz6nlMWqJjdzg3uMPMLyNXvxZn/fV1eWnI6GwogP0EI+h
Pua2RVgUdC59h0cH5pCGzQInVusVjjWrmx3w6ZoZHdsd+OTMuBG9LZaTqEqLAiLk
vTZoJ7iusjKx+LLTN+hrA7RXzZbIjcMYDqCBz1HatXp097PLl3IUvT3l6InhKFqY
S58bVlHIAgrEPcLR6xUboF/2WdJxZmOh9gv/fN5P8EL34oQncU3CNqduIWB5pMyx
8uVjn91zK7S0pNyKynORhyUrnjJ+RoDRYk82M/EmbsIkl4v8mFihYvxlIXRCx348
r+1mAMRb1pxtcEdG4bNEfmTqdPBlVj29ae9fKJqLO4/zs05C0KLm8XSDWJy8+G+V
ILxztqjIItJJ8/zxJuL0jUahU16Ky2qBW3aOuHNLJB7DbXuUZwJ+RPREgwmagFi4
lELMp9ZodrjBFrb6cSyEK6IpoBOIJfqwapQkSimMwsAn/0VhljLXrpcbBvuOpOn1
oyE/LxTEyWchwqEvLoO+OfnOO56hF1sK3Ry913SNaAb5U5Jx+u0OZ9Ag7uzuvsKD
3Sc+lRyFQtBTu5f6yeKVtkkrofffiEoE/Vk1azLEtWeoBubTGPz2CCy5WFsYeS9h
yeQcMsUGRv7dQ9+uYFhel/sKHg5G3IDksVwEYaScQBO6SRMXv6TG4VXFLflb+pXw
sT0Zbifiq1yVIYGZe1dJeMsyqVtqEBHzmm4o4UU2G+1vaVSVXEz7pSmt12tGhPMe
scWLlKqPDyFJ1LClvbZeB2dBZAy46TezlFVCrXE8Lq6nfWVuPk3hszHe/AOSnZij
aHx5h79KWJqX7k3DOmUyUenQbn4BThHDJctCyV4ZVPc7BimF/rbwIoFbbhsjYAw0
pi/KqgnrI7kMq3i5YIIsx1jFnyTXprj6gVW9zNux45/fdtUIVjqo7S9WHKDnJhF4
f+2LiODJpztTSzDa009IN8rys4bHmumF6aMmeDCuTeOWtG4ktDtnammA0QQ7qP/N
I1hZVU6w34dXNPmSF00oixrXxaKa6l2sW6vOWmOGc+Qmikz1THhvBS1M0puiR1+f
SNZbVGyRge6w2doj+7ovtTXyUBpXfrrw6aIDcnzCX1CQgv3mq2CZpQ//6RPIUyYl
Tuq+QSLOH9fOXQZTkiRXLzZRptjHveVBuNCwNblZiSOVBs3qIUN/Z1Q0lCAqYmCv
BotsFrRjNoQWS96qAqEzrxTHK4P5CXEvjkqOFJPcn9hGo15yirly6Y+OPCOPo7nh
psSpA7JbOXTq/NkFd+PeSNs+w6mpCkvnMnEGHkaPqal8oQ6RDtE73Uer6VqyFzIu
6MGVBoGUSxHtFMGGQipsPMmAJ10dMg+CpdohkPCEnrykFIYGQAHI+SGtFZVkvPAF
5yzb2cmZAxfMT6AkHSBIr5shFx7v2jXcWt6Heu93zChQGnOnjFaBulEneYf5iBjp
AiDI7EHZYHvRKn5/CfhrifI6lS5TyMXKb/WQtKsX2RoEJFLk9Wg5eX5EZkqbdJu3
ELA9CNnt3qAnfHdi2cax6l7rFzEr3YKBvNhS09yeMl34Fwz812YnoQQ2YSqYrVRR
Acf3NLzuTHkDIo/OR/GYPxXckpR48QwGbA1s68fM9FPa/21BLuF7AQbTIGhBN2Tx
lkAZhqSfArSFZH7zHOPUb00g/c7d/U/RTfn9f4PzyVQCa/qcXEqubM4hWAKRskF/
8eZJWwl31XTaESMDvkJDKdOr4XREdFUejalybWUDMC9+he9LFkoFpP4brzb5iz9K
4DEkonGCCX/sHThKnysBGcEqs5p9WILTzcIl9Q1RweDuydS1JPWPW8bqg7Hj2T2y
JMazIA0GBP7EyU8cx4RNONZguWjEWe23zHmv9StllN/nDnLuAo4UVaHX3N9IKNxr
hvV+DrF1M6S6a1T8RI+n+saZw4ypXnFqsCgpKSHGMXbQ0k2dO/th/g4laaASHYji
XIJDHy9Nf0vhEAbz4LOy8WSyNINa5MOwX4CV4b4ab0+WEwRPsUVmjWe/5UlP1gl8
A7L+afV2Ala17XRhyiJ3g+LKrDFHrCyiKWH2arv+N2A8l2oTM9xxw3Es0wrpJLbQ
971gtzXxbdQ8ay8XLbCwKHIb4TPu+UZEJ3KjvyChAPOvkUcYLd8kLWp7+zfkdOmm
DhBDqKdUU6PVj/AOfYYtZdWZSh7qeTBZQzF5po8KzmzC2xWkFuZnC66Jx5W2qRUj
7k1dnvwWsiZpkycsHvwzXx2puzz7TnymPjEK59jUn5vBKqjbLoRphBd26A+mW3qZ
p6MH5q64rj8BID0Y8cvz6Pv1HT22bCjuU2t28zYzXlA+N8cJYA0mp3z4KSYMUNxb
v2EF/LchnIfZnJElFTEwpRq4U6f86ycvaFt1PtbT8Fz1EKKeBNvZ3yfqkHJld+9X
SNTEBn36BKT/rZ1HTAshYmwidjvfarT7BSMVulQtKPE9u4sEqSvDmyojJURrWFEv
ZgDEDATMO2Bv++PI+jUKYhBQCKZj+EtuKXiavIYVpjY60XV4WKJZ3y7olT+j2iMV
tU27+BMMQb3Vr/Z1zbLMT7qUsHGh6HQVvV4f6co+I1PM5dP16TJk8EW1JxEwCiWi
t1KRF31dXWvJtlecs2TyKLEDVt/ku0cFDYIHHAB8//bWj6BErm53TgXePNe4usOq
7S+BBsrXgRChgY9rAB/au2pu9QvOBdz/KEYRmBSANQ+QTJZgFH/MrYRaOiSb2zPB
ST9AG2wy8MD7RuiQMTvHodawPU6oegsrRaeA5KI7WdZLF7mydpEJZh5x/M7gL4BL
RbEMihfJhtJuBp3qbHKgVcezS8JXvJ+w5DKrMtbOjFM2LVUZMoKNCA0vnHZbnHYr
bjgfhFyQ40cKmsFFy+gTOjIpexM7+8/12wDKkj3EmeL6eWmDF15ypcukNzEzwMA/
qD30XphxOGcRjqJjc2MKNht3nI72MX+baWvIwHEe7ulVn3AZToug5qiRqZEP0rV4
Vu44FB7DWTQ8GxsxC6bdFJX4SFOJR/if6K6EHo8/s2xSkMYLootJMKzxr1VZXwBi
6NTYuomRqLQ0q8h4IDywRvNQKKFgPhgKdKC111FcvmW87GZdi084Xte8lqcafdFM
UDoVYat24lCgO5XBAyxZnCXatI4nZqZlV6dqp0iZ4lXPz4bxjLs1jzpAw9AgT4Nt
5XCRmJTIOHQXGl2x+NIOsOOCRIdFFk1qjVqorhY/6w7hbPjwNBqN3JyEDxWLw1LJ
m0Rjv2x3GSyQgVEuLs3DLGcrF8OSVs4lqUQnIz/rnkYvAK7HrMtBv7mgrbL7r9qW
1foZhkMLuQIXXrt0g3sNG03mq1zgT3tFFaxqymddmvyKDwJGPOjfcAKqoaQrx5Ug
xO4RGZ8JTtLUHW68V2lFfkpAxMh2QJA46V/DoGq+8pxeS46lNbc04taYLrdhQzlr
PaRqL5OzryEldt8hIg9jpEIOtw0j547J/m5A+xVxFpLYvdxyVE2Zy1oH0vjgE54T
MX0ouIEFO1X+KPlNiETvAAAiZBFCAuf0l9MSgfoyXvpLABlxIwhgrbN+ij5Pbv4t
ymC4SM7wtGKsEMsM5Cadp/cnAh6r7ivqW65uz+ILaRDDzXKjvBFJne5D3gTG7HIb
ETAbce+h8a4Romisy3DcogIens3UdpgJr+yHaeILMbQ/OvgEREuUbkix3DGtREf5
QGgTq/3IfCBEkzUIE7uWHH6zWUUq1gLIehwbGi0eLempxZ5OAtfUC44sDjxYpVNf
ziY5jLv46G652RQ1iTGTTKrpKxIXXlRzdJuzJ3eoP1e3wE32syiMyoN4rzwmr6uL
GXMASEYYPoEinYuGXk0sST5QnLE7MQ+UBSb8UuLW/9/FdBJV4p1FkImgCkssCfm1
H9d3pFh1p/PO9aGy1wbBCWKeyEfmMLFT6OMTsibAE4L4sIywTsqZvnQfTBsXd4PP
lFrwiXYwBl/1R77DBhvqsKZL58MEtm2J3axgNT09Yk85mbRR606qr7xvLqV+4v6P
W2gQ33O05McY0fdn3HlvGvOj0cm6sAxu9tsGXViww72drx6/sR3HA2KvxHvXprY8
1hW6Cjd7vQnJFSkOzxQ69XhoLyC+Trd/6OTWcGLDtqwe0MstglCBcyaJwkYhKLN5
HSi2xlQRhHErHWp6tm96z6YmhO/SEoic/4kieiUomzv6B5u+Hz3MI5QJbBRp3aS/
RlgFgmdwFlIHBYD0tTANysIVzF3LQLurHhO+WfBYan8jKeo+yOh51LyrZ1c++M1p
KmxrPHXIeVj2oXRCH4vpBxqwJ6ibKA/zV8PH2uRsz7eNHnK+4WuIf37ZEMSboJGP
1POUMsWtie58yCbXKhwjW2TQ5xrntfGQsfRj7d+ajARzi9Lblo4HCe/Xe7KOnPQB
z5kEqsl3kO7gTIyqzNkq416/QAzZfC2gH6W+1ElE7Al6VNBkGGe/X4S40WKKiaFs
Iq/WXRULecUslSULad9UVQXzm10YLdMyES5460uWem+lteZ6NxWBC0L1Kih4ykvj
G2ywo/i+LYDDDFcbDkxHQ4YI6aZ0/GjmpjKUvNKXxsJAzt3kxcPIJtAZO4tSeZaQ
iH9QKYIZuEIpV93hvV7+/Z7DgJ1lYOIri9d+Cc42nePr6zMGk79raiyKHYFSHmbQ
xpZ+awgI++tra9AB+5FNe9kfhIgnkbeF5ktndrrvLI2G2CMSIkCR2zs5L/v7s82g
j9TpnLdJVrRLwEO0ngAAvgm1Z9cJlsIHDCVo/8T6by5uYiR7TMtDTRLsz9bM1MvP
1HxQ56bH31zSQXKKjAdBlkreG+AbanIKs/1H8+kqL8e9JazclGdVYJtikQ7BZET+
q6ufIUjlrOZMUG6R6CzbVi1Z4gtSbs5fUzn1kI8cgxuJodRmxyF+7MUX7wVQa0Po
f8FEN5FY9kXrpHlbpwcoL5+AXP1hckFdR7PqVwJ5j8BbUGccqNHH4DjXuEgG39Ve
xnptc3zFVBFFStmw99C6c7RuJS3BSmqkH5FQpWM83Idd6UFQCbUPEBiuVMDSCBFt
jUQWd+WpQ5mbKKqWdD9gnu1kpbXVDQWAAMfwqRMcnmhTKyLHfU0ua6Pt1aWtJUxD
k4hQIRoSBm5B6XdLnISOYlUXabekbI3eJCDOgmr388WYe7bDLyH6L/AcWUP9Ua0/
EJ4pgQoudEjMNreBMqEnUihKChlLL8c7e4zOV5GYiEtY8g7tO0U9/oE12Ek3jUkL
nDbqzUtoF217eXwvxlyrYUybPrqPx+bGR9CME7QArMlefCJNkCAizZj1yf6XtVGS
On6Z2FmYIeouOuNrtAuu6XNGkhX9JJyhLqkBu3k936BFSqCqUDmgCq3sb4d7UqBb
U/meb/XEzqTI+SBewMKb5OB0mQLAFNXMPUkOLghNc5IQSE6ZsmBjXRgwQy2rY4gk
JTyEyUDgguPBZeH/pkIdIYyBw7c+IhJZ9VknMvVQEvG8aqFLhrXnc4zEgE+h5Ekp
JspBmYhDWqHrkXIoJzDE5RyZRtojySsjhAclZmq7ojKtF3qsim3L4kiOc+63OUjF
GMj7zpwnonT5XCqZdl0eIGLpQHAlOaOcdIHRbHMJ8gs3boU7Els+9RD8fd53ZRjn
MNW8BPMR6Bh6khOtYsRR9+NVSGZwen6KTOQkZRi2ElxDup7NDWfFXllEeMIhNMNu
57vVFSpfRyMs90espwX3q1wAWUtDMd4Vbaa9jUZ+Cu2ca28hTjg21gV4je40WTCA
5z7JNZX9ShsaKNiZm6y+UcXHUyELmO3PJ1TEicHpa+VcD6cfACeZCcKSFCF+7+xT
M3y0ETj+m+odz2dkZrSHxg9cngdUPtdhyWnja2MuydEkeFpljwF8c3kvOMDwk2WM
Azv/s0j3HfwxNI8uzehIoXUIw93XJSfEr8e5A8INceJfE6LETXZ8j1U7/2X4J3ss
76NUPx8PjoiLMBSTYI/sCn4AgorT5vc3ykQOiepWeiRubm9l5gPX+o+9mW/w07kI
eNEuoR5S0tbfG+T19lJJD27zeqkHURe+OlMdifF9ecnPLicvOSDDhrN4V/6aSEfQ
8AC7gdY4iNqmXBrMfMSGSxUTdIgKbuAxWXnxLPz4BXSr+XFV+NnsRwsX/ZKLEgFm
bxZ3jUgxSvJ5S3uThGg5TFXy7vakIHHF9R7cmnfQmGhJ82Km53BxyRCQ0nbSvlwP
xWf7Ci3BlwyNxZpwXAHPcCSfslobA4Tlo7cfwcMEKy/fM7YjbzcPdPIcXY66+Gop
q+va5XYuGvSvjXfI2hCw/1HlH/NE3FMGutSYVmixmMA5c52P2VqZ0sLnsO89rQOQ
mgK6orS3cUApk/qcCkzAwYvdFJRhD2aIU3dW1ps0gB68G+necHO7czeoUPiG5Dz7
Oj3bCfzARKuFUFGHGo5p1rEkcDCZWvJQOF0Rui2yzX88x3NNGlRagD3j5dMoXCo8
P84+rjH4hmaHSop1kt0xo/8zFiAZ+ST9qVyRZCFCrwRN1YdH+SZBvtFn9Zc6k8si
aTGhLYcLxC317epKil9XZce0LGn0Y7EqPOLm37w2ADVhtiy+AnPN995YEeAvr8fB
76YUFRSz3Y1BXAMyKEULWP03Y88lTg6/0Sc6Zxd0ch/AIiNi3SFF8w+1wc9qcE9x
y/oPGeipDHa0MIjw8FDiYdTmiqGWemdUvNah7Gz/WiZjK+6+C9v/HZ/hGcLwjtmN
Zw7aSxd00RQJ1RN390edMKIdZ8d7+lGnCG5HTklkbi0qpeIq1v3E7jHoYg6Umd80
Db5DydxblFG1j/kyUMxG8VEWcc8v/0tFd/F1bezqVY/G90LJYl+EJzyKCOOUwxwP
g74CkEuDbFMxF+Mw1g7wkSyiNd0v3rOjx7/XtBojMxppfxOfiT7j4RnZuVGGFpeQ
9+Z26acva0zxbje0cn1Etm0GD9/vbizXGDwdpGB27PhmvSjH+98Etu+SaKXOni3V
Yk/kNK0P2W3Vw9mnr2I1GKK9PBRAyFXomWPTXljCXilAV9rjGaGTdA4u0r7Nv4yE
0vyJZTu1KZWQL+/k+TdME9YP4R4tCJcbj5jfdicpDE75jSu1+KMYWWO54GYLEtQ7
5w71dU7TGK1mVGNFIjMPP3/Ec8WnNdPALVtGVECQSOZbobT5Ga0zAXPAmCOI5PcO
TMUdaItL8R0lF5EqoZoEt9moJmqmzI+GzGrJHAt+JHpB7rNu9YXRwRIdOkhka9Bz
bek9/DzUE7yYye5i5ff7WhiHmSAiBBqW79GW54tBbUqrcEdN9B4zIfPkyq3KoAIc
sBQgQFVj+SoaVq8W5yR/OI9yqywqDZvb3kGUBGqycNWXUi4Elw30wZ02I9yvX2AG
Z2QfX2LLhVG0Z1E4J6j6EN9a2LPk1XqMshaPkf03XD9R6hrFeztRryrJEaRnw5po
yCDq20KhzxMmvvjGsmcy1G3TO8jQr4t9dPRklWO5oo/H12P/ESWCPBFXSCy16AZj
1xyyRdOqNUvOyyffszrb6gjkI9JiCA2aw9ewew9ARy8OHfhSQAbjjm2wWGr7EZe5
0lt6D1+k4ogxdJ6FcTRUklcirEYoKNCpfXbkXrks1OlmpsW+c10uk2Xa80bZ7I4x
O7fGZGG9CswjwUJvz8zWgn9AFz0E54UxaBQi+SB0mfVvxx9gLCgFal0WiIu4sk/2
uyUpj+XbuJ7zZJEXF1+Hw3mHWAd7mMKVADka0xiz8k7o9MQUig8ARRienl3eNHzZ
MyiVL8qOPSqUuXEXtMwp2dVYHvBGPUJhUHypl/2+/s37IVDZgti3SHg/NwjcyJ+5
NuBQs1CNcUUvmqgT8YRIE/vwEuoZWh6VsrpsXL3DevNtLFG4CLPyQEwmLPa+fxmi
Z36nHoX0mCIPdNKDV99iWx9NRDe3KEjBp60Bnm/QZdD5OJMfiuWTYfzgD3LpvpXl
PuATK8NIF+bfEjHOLtW6u8eEKO0uMal6GVJ/QGYEysNgoQajx2RtTFI0Obk/qSb2
uKkGg5n0y82GLwBqM6nRvAuS9gqZFKSE4RbkekANLDyCHBKbUsockTLmgf3sEkeB
QKgwBQFuFvpRCOpf2psySJ9KrM6u3LQoYypoeIX0aG6Aj2Gq3Z+ISQ3GHRLnWbcZ
1BsTNts5zGCDh58RrOMtpGu/4rP3HbkqiJfmrdJmAUEgpVBac9PB5Dm7eW577/Za
XJnCjEDw4vZ0u/JMU3nezpDZoYjf1QrsChQs3EpeY8J5HzRFiYC1mKLGiGoW6s8X
ZjTBruFK9RlgufpgtSRf1lekjTu9qf0z/LS2vbwKjeL+NqsH/MRlJ6CYqSjFL8Gq
pbCBWFuslymiPyhEAC0CcUXKLsgsXpYrpQ6NO4M2uIVK2EtgGtuKlHlsjN6aTKVU
biKkS3bpgS2Ds9l2+xAXxSO+p30u797CArct5qPvBc2cbYEnQb5xJxBk/3g3HXFD
cbkh4RD5ftG0c/1ycC1ESSQak3t1RqFe9bQImbKCCWpz95ANIbA0ZYi2Auwm9uDL
XlGvQ9CFoZc0EQV2HOSidAEUMCxd7/YOH3hvLk0par1OhhoX+cNjUhkjhtVX8XuA
EsNH07Be2/yivbradUJLAvE5QaG3PoMhQNPCOUvQRRPeD/4urjn1m8ss0KeR6IcB
e8jGHQ7M5vSeEOWAQaFSTyIlAR0MSFtVVS5EjUgVCGqkcy16P4/ltdhr2vNgTnxS
o81YkUj8WN/IoIBACeKdlYM7OxfbyTy0XMEcF9NmUjbqZfMCZ58Rf+Bv0vhQg0wK
PCYTEZE4jmIdnEUaHKl43ZHfsKP9zEBao76j7phOUnoPbncj6pXDPZOXmp/3ZnYm
OEGGU2J5TTKZDbKADbAkQaO5om5WTLrwotPxQWFWw+JdV3dewcFZsAEe4y0cO0gp
KSQWFOZZ8dFu4JhVz1eVUYyxFDA3CavZEK66e66ZXq4XOVrnmB5P1gPLkzUGoGji
wwSOC36K9JrG1dOuxAXriUMvprbwJcUhyLPkRCZZrUu9IqByqXiQoQ1oChz1xYpW
EiaSoLWN+PP87zyMw9NY87CPRG0+c1KlurqSd1GhYMEjm1HZHKGnHwDSWNzlVrhw
IuL23h1mbJzGVPsnlTBXDJJ5sga9+U9surP0unQKsIonfwdJUXmA5U7dY+fnhfgG
LOT3pA5JUvn+TeDApAxUwTzkpmdxUNG1ncVsIdXDGf0RqlIvjKAC3TJ81BG3AJWI
SBnfBSZ6Xrng/e5qZWBOjSSevlTPaNaFrQGCElXYbQEJrUBJq2yC/XcfTGYxBsm/
eo9ZT71ATqYB9QrV9NvokPhjugPlqsEt8HwIWMVMetexx26KOh6zZJrAES8SgZFr
amC6gz5ZAWjmzh10hpPByOQifcN7b3ylOS9gHOUw/XvHpv5Nq2+ElKGeewBnPT6u
NWWHQjrjDKVNawaZ0wWsd0G48qNfZXEAekycxsh55Hkb/TGV/YEDlMYWAjoXqr5s
gd5sr/ZJvv+0fXnvI0W+T0ga4UcFNDbhjKccMkeGyQ2oBXgSlgTehXSML2v2g/6R
z9Y4NX3+sCL4LJEVNE5BEqgMaI5kgqoY3sny3XTWBj3V+9zhcCxAQY9pCsAYBnqx
9zNZEvfqr27OUT34ho+2wAPFBeMm8LWPc6DtvtJU6oJ9NyNvi7N5kja7ZXqjwhY4
M21G3qev9w/1IKEJEFrpfOOdJShAAelOCX6ba8AP6mjm/vIodhxCYHO6e1/bi8Y0
pUmvtC1MFFAmyzdv9ifyAGf0M1shORjZigRDakAwDeOD2fDZ7QGeTYReYnCFfarT
xg/anL5oLZ3z6lDdM+JmnQ+KE0e8Ga/8fAKRECDeAAA0oCCFgG9mkEAOZ5Xs61H1
It+p9x9G8l+HXwPfiZszhVvvrvJu1146B1ERu8V/dhsS73DnsGpP0/ib0h1/3q3v
vCnjFNRY/dC1H6PtcjQ3oCyfuTYr/qAlN+7nIH/c9jytIsLXuPRIhilQ2IbXXFmP
1w22H1OjW3LyVzhnnFRpS8PB7nDNLUalBzf8a6bnxVluBahr9AA+3tfDaO9Uotcd
54M+StJ7RvJMYDI/KNsf4kBgi0YIW0/nxgNCWg7L7oHgoM9d+mpz5q8K0KZV35Nr
YsVInzMn/1dT0eR6DuPastuv4aQMTqFloSobrLIAHSP9ANt72R1oA/t9+gi+eT46
b7sDyE8It8ig1Vg2Yd2t27Sc+nTtDGsWVcMJs0EAhtHv6bb+NRB2yR8qOQw/LwWP
btjCqK6/xSZxpVhdHon82c6oGyeAkn8IMM0HWzGn02N4L0aerIXO2EN6sGKEvAcp
/zsZpsVO7RX9cSuCLRnMqEi7B+iJia3EV78AjOGocyNp2n6r/1ZSXEBWC/g3kGmE
rsxO0TIzdVc0jO5u50PDG43y2KO4/CEWjYlmTt8GZU7JpenmHC9sUF2iOskrofAI
qnRCE4q8/GbJ7KyyQNaPtSgI0LtdneXPptyrpcbEblERG2rTl9hOTbUxB/X82PCe
qCd49hI8DVKQz511JYAzJ8zmMpXbx9UfAe+vdqNoJ0Qlg10KnS0/5qdng/8BrjXx
0p+NI1RNpv/gWmwMez7SqSaMThnfAwiGdU6XMtNrEZPJaI6xPL2fnNp81y4Q4/W2
MSkMD+Y7VZCFXwriy7X2jpBQKJ0t0Q3eFrqf+mRmHAT2pb41CqQ0yFclN4cylJzi
HTAshsEPMEfnZVtpbkse4KmJjDFbkJm0y3MzGEZtmkhzO0ra3HiFOJ9Z5Yk3ZwpI
HrMZ8+OLSld4QcB47ppdiEm44EyZ9PMzpDXUpnT18jpdMJsqvSinleUp3NAhfo5w
MtcB5wxt0HNU4KLQLtxKWfYqzcBUzoRu8KkB7fNzlPCJ0W7+CGItK0iQ1pAWWwN4
wRgeKyfsls6ZuPiIAgm5vSDDjptguFwvYAJqQpfqkzqlwbm9P6GKC21aapprdUzB
LadMNJE4yy1iEkgzXfBza5kLqY0pmdp8uuG+kztqGPr31G1RH3dpaSAjaSK0U6sO
CcCHdj0iWZOBQx/TpYJEIr6YvIO2sgLjaJqtosZpAHQpxc6EBLcTzFaAA/IIrSWS
G1YGrKVcnAq5qUP0cwHTGrHt6Tb67nZg1qf/ybweYFlLM5cpf4FaQM5PUcSgJvS0
9o8Z5spQmELX/mlki0y40Aul315ogPlZjFng0iB1ZSieAlcppVCODhC2gWR/co3F
ld63dkCxd/K5WAu/uRe7WoX3A/3fsNggXzWznHNjAfNTV7aMrICqMX/L73YtAqE8
RXja4oM0GqmJS23oUuh70R7MyM6hEdxlTB2ijLtLx7qjNjskkkmBU+/paWdIctkB
V7/NYsFPBrAJyp1/CpvA9j+GIL8+ZfBDcazVem1GNsADbb7TxoF1vrPYTVQDIDRD
50p9fQeR2EscDiOXXr7qeAxDpdLUFXO3Tb1Tx2akHfU4o5fuwrAbiYo3ueNc70r/
EqZBpu4EBHEs4OlI9n6ESTdcfiyI/cBlFarkkF6gbaHltVGUtPUTH0eSlM4KyJph
IPsAqFdrinDjNwvs4lt2qVPYHNdPO9h3pBH8jRbM0gTlj4cBf/AUH7SsNsgRoQdf
lq7G5tOF0J+XYuzpACV0Dr9K34MLnNfUsum0osRa8wSOUR2OPOMqDxJSZ39/8M9r
Wf2toTIsOdaCsp8pvjcOr1jDm+C2qbkwkA3sogRzsY1cUlLxC0T8RMzG03k0kYxQ
AgDXEKezy1Mm+Z8CHqgjArNfrxry7za7QuHf9RpxAnEfIcoHWnRtDB/v0rKjSdbh
f6TBR+fkWMOIgLEFSMPoctDvt4pNFZYEdaYeiXdaQvWTAORu3B0OfDs3Y3dJzOd2
JGBTmTTSqUwwEt+mEYDjW8GfW7IHA/yMTE+IL4FNauDhFwWApPNHBJs7TzJ0i2kR
/kNSksH7V/d2J7nf6tb8yVwyAVJkLYF5d+U19hIRUG0ScFnL/1U2ims2fiW2riJ7
y2NMPveZ5DekwbRFghz4qEVLIzYkZWtsCAerp+vFpcLrqtQp/Bs8nH78E1WAPyk5
iMMDRSJUd5jBJ4D2AYxWe7lUE/Xm1XAH7q+sInXvcC1aq9cm9JS75Jg6ywPPF0kJ
YqePjFUeOuLvK7tSyThZHpoP/Lg9xCIvpsatSQTWpMuCTqwag/ABds1AHEtr1b+5
08q1nAujjyFy/Ua/QV1dUxQhmxh5toR7Kav8nn2rC8qU1YmivCS4wzB1o08rP9J7
wSdpQ9F6gMymW9Ye/pQ5qsttg3ULDKBQL+ioIL8PG2THZ7Dg1tc6AVElseL4eO8n
4Ytvnm83OKyY082vfc5qkEnbl80bLPoHpZB1baMTcxEa1ONjMuGJaUP2idUBs8BT
S3osD7Zjj//Y40H8kzP8kwp59a96VceeTqiDxpkvgf4coJHbIZExtTGWeWjU2YtR
BmoJWIW/aJsKtEjpGsQSGoplcPWWaWsGCc5bmLBgJ98LJ2Q6orxjO/tjcPYVn7Z6
jhrBn3cjyo5ACpGCC2SG5hsHlLVoSQvHNeAhzvV7ENiJm4lP5XyCDycg7kWrZls2
KMrvcT0L1ndUjwzCDBknru9AW0sVJ/JAaJn/4OFgN+8VEE3+LW2ykaaTCdFJDVPP
HrsoSaUHZxIrqYGNlJfziXkfWMHGGN+3R8ALRzWykM3va1K9PWM1pf0r0kfG5Rg5
0q2jACDxS9VqKsLM5H4nrFA328Eizi8YG/s7hx/LgW+nZl50WlDgsBfumuoKLgD1
UvJ+eAGuoMQz/ThpZ9rfTF+ShDO20eZTrvTvQLgqCDJCrewME33WWjEMjb3HIzL5
zgIJJr775zMzcIwgkDrFExbWsJPlw4QgDk4R3WEL1dFwEkx52AvySuP/5b89i1kH
2fsefOV19mZXRZ+ChryXIEycP1bkm5kRYU1a+LFEi82A+AjwfeRVP/O6m5qfMejQ
aGn91sOV2sngsj585BWPnOap2MY7p5PJWJ2zA6dhDeWylT+cDUlofOTuY7oZ6X8e
We0E29NG+d1gJpqTTYxC++MBE74j88/K33F8t28Zhcqypm/Ofu0T1hgSQbJNK77X
brIFE65jri1kkr73uwdzJYyOafdI4eLGBCrcVkGCdPwnJtPmQpgZAzMqaxOB00Og
ZUiA+FdCtdr3uLmYgU9ttmu/YeBXvpjiQKOusCqW+y/afWpg9v1S4sjCYbObMOzE
phYSl6RQWYUmL8kYS5UVgEoetlswgHX9GyY9TyEfcjckXF1h59aNsvLDjSaKZOmz
Xr3eOp0Xmkdqjgb0SKoGJfLWv+w2jZd4dBY04Too4pGO04VOQIH0dBpPK9JZT9xW
Y1oK3938A++WqFQHWrxZbJ4+zYDINAxwHHrE9Cp9AtRF4WFgQULjPJFHSO9PS/36
3jQsCHtwA/xJuPmahf+lT4yFDjlby5u6xQENnZnySjxgZreFUYFCoK8SEFTedVfC
ysMI9mhJbrYXaWWJrhRmjLU032dE6CpPQkgt/UOteq5fX3rFMyQCoLvxwMXD6can
UT41r4UCkLd0YMoGU4/8wavx4iUjTjVAMyABLTvueJP7VvHmAOtK5qYo7FHiT21R
gOR51AhpWLCp4lfjGbfJp/G81qI0JZuANTAxgEJeZeMNbOWUCjQZGnuQ3pHToO4j
UqffHlwda9xedtQf3B0ZvI8k6h4RLnv3ezdQJSkYWE7nZSD19782M9vHIWTnVA6A
cceRdVhQ8aH+KfAMQ7oTaJBUk+sZ147TQxJv2pM36/Tb8305tQhyT5Lyh+4NPtHG
7a5egc9wylXVo4SFlBqvrjsVLENMg3bXxAFMumWmMMqB03eLHpic3Rc6Ke4kAobA
UrT3l+RxKwYFMaEquvY68CaLGKvRQJK/NBiiD2cogn+WRBjyBv8rJqt11iN5cwdB
aUGqKZeU3+d86RZe619MU5/M3ocd9sp1Q+S/2IbBl4h4KKoNktidBQrtQsw7grlS
Ey6ZF+B31gmNQUcGy1W+m7wXrtW1fdcRKtoYlYQmK7udWxx5mLOEvhb2/SY0JqTL
K4HRF+OWKvTRQVgSXK2eOAqRhzO+CLIyGSARGFSrUmpUh6b8LAr427KKAqnF7OKb
kN1HZK4B/D1TI40zrPlkfG5pPtVreyaApNGtdqvLoVM54XcA1vx0m37Iw/yJlxHV
ST3KRj3JORQsbBm3FVlix81c9Rlo7AvPZ9YUfHmNqkW7+MSnfJQ2o4VoW1shKF/e
j3jMpjwPeu8vSRTx3Z2Pa+AzQAGVOpEJm/GxKeX2orZga6JUXjiShtt0Yb/kCANc
i1K7M56yGlyGTo4bRHWeuCQ5C6+3wkTtOaPu7Zvm59F3tbTzW1P5FfF9reg9EJ2x
W3jzTlWU1XhxSeKVVsdbt/jabp0D3C0LGQ8zlvQqiSTe1v2S8K2p593HoXKO5HgE
COyH5gxSjDLC9C3Ir/i2NLu3iZDE8TrONUUFZ8JgFK/8tcucOXRnF2HTVTNPJwBr
vTIE/hWejUUxE6d4/vnzBWTH9fm6LTjGVqQt2g3AyonTZwbO2eyCT88H3nqlvt8d
+6ehdcUnP/WJNI3jWAKgrouVDiuqYZFhy8ILa8FsuJfWfz2V5Oyt4HRwfrI63WCB
KKO7AmpUjG3GeusYxrmURVb/4N0S8QGp0s/JAiu5rc4xr4zj1DpBIay1SldhUTjf
DE4XiAREbujxfUoLG2xAlLG5RIHmT0G9T9ijrLnHrXXzVHVrUv/b74PU0xmcgiXn
+feY7jSU81tYPtsR9H42RAbyfETWoqYazZVdfXiNZz/NgV2cp8lQOOFcqivrMM9E
G61iNW1cBhd6JOlTV3a7ODbMxlNA8Z5hMAQecBeE/2AuosENqkcEMhIj091/CdCU
WdKo0sGZfEjQ4hxMLvgMrX/9/Qj2T8EVkAGV7bk9xwq/Ye0c5PKZWEqbiQqBz1FJ
SC+ANFKPIgnWJj9AuTLImvOcBOuEDAusbF6gbK7TV9fkqQ1A5oTvmOxJUohregxm
x5C1+DfDfl7K4ThKVV4SV5QKhSynRFT+pm5QvHwVe//qfHDeiYviV3OmVmCd6HNR
t6jdqOYoKkFxkxjS3QGqrDf5n6FpXgCquUKFmZRPVpvblKNUHtqHCSHG5QA/YdQh
0daaA3u2sqZbLZshMf5XnzVoHsaLRbTWCZCOz1sQMjxW9rfjMdAhlrFfkwOXzI0f
DlWAOpRAp7Qfmunh7eHuaHoywv5Y5T7kfmuPDEEED+e4JMnnWPGmRY8E3tdpiBz8
ni27OFUGh4ETtCrFFskzPpPC3WYvlAyy3TcorEZm0EVm3kkSGGeWKccAtdEPpHL+
PH52g/P1NyRJ1wAafOfRLylWEqhmP+A4ia786wcwlGJ/bdO/LogxZW2OE0Etsqg4
2DeOwz6hCjrTwrxMOC+mZIw/3C5VO/bYSY9/48u3CMCV2Wu2OfETQWfvZVaZt04E
aUKgChMiN0x3P+mQhF7+1VBClEg/0ifNUzHCw+no3hnk1wLipij+nKTS1g7CfBwQ
X/Xtr4jEiv6n4MPfJbQM7KA9FnTGnHxyBPzjoGOGx6Gusy1fv+NhaFrdf9theXhw
40aN6pClaqbX0k5r+NIPS8yFaq+ydZRbmYnGphi5WL7E/kmIFbOZBYk9Pc+jd2Za
8Frya1jGcVGtg7a49iK4Ua7R8qvcwmc8c6o5viNqfPMNboyANr+paDECLwF/QNyQ
Q8FPuMVYg1AqDreelg92gVW7//15xNgarggnLnkGlhpeJePqe/lkzQBtiuiTpLj0
GikSebl0P6Pn5zJzXVPUJIAlb430SGz3dCQ2ojZSKNVvRW3AYQDSMzyL9E9xzYY8
EoU79YoBAGlK6E7vH138PRW2hmdTMwEa2Hoj5TgA4BztsNKbOw9HP28fCnwKtgcI
MtmRhOeMAv2HQBmRufGChsPp8HXzWSP+U2EboZ1x+sNOFTh/mZu0oJrIP96p35kX
5tQsTH2sCFGX56IzB34mEDILxZB1VBr1RYOxbRT73avSlxb1WrxGLJnFK9SL/ny0
V3eTX9j0j5J7jbY/gw/3vf3uizx5Gzn33VfiPnxioaD4XosD9iQ4ouuY3oQrPpVY
aA3AdNo96oc0TEOx6ZKH+WVm+R6r9smY49X2MGSC0KWwN6E0Q0HO52lk+TErAowc
8ea4q8n9XW+DrusOagqo9n19ytcJ0hf6zZ4f6Nf9cJW1qZUrqX71U+uqoiOi4qPE
6R9ju8BQql/tInSehm9v3B0OOju344hnGs5a+FLHRfrqcax2+zKm5b+M9rr3S7ry
y9tbMMNyj8lU09W8SeYII7xBv2taQkNhrwIiq+BvrQN2J+xPx38MtzQ2MntMIvo7
Z0RnuFfC95ZoBgViSUWULEuRpkzYljGxnYZoa2FOH1lpSzFexQgdLuWhTdQp9iub
PlQVpwU7qBt2GxSdTdp9qg4kuHvCdtDTP4jWV9RS0X9+ei1tQZXuh8FCnVLjNB1j
IxvVYz3jBEOPMZntO6OiLokXeM4wvX7Z/fXwDIIKxbPYlTSaLoO4tQ88S5uczQKV
TnCjsRKbFhJYRQ1XVt74JCLzTqekgkputfVsC11OT1wUFn21xFrwgEmoIr8C/LE5
xyfaKEWvH/JTX7ez+IhlLBQsvZl+uSxlaENyhIMsobgECoW9vAhgD9h+3WrQQJuU
9+EQKr0ikTp+xrnBySHNi0uRNyu8JvHkomT3UxJCzgPBxS+lBoscjywKeGvKyCFk
7fp8Ks16oRPEd59arT6pGVOWvLemSzdIilRZG7BqyBAXveu0a/fvXWQUovwJbpBs
qDx5Sh6aHRu5bppQgryWGMdpkXXOe3rBAtuuE0Id+nyx/rQdIv6GoK+/9J8qUdsC
SXdJy+RRgJzf36PXQ1fr/O8i1aICZtQvOedvEeV0aNAumGMDMhwQW/iplsn+dJrH
wOPBp3BoO09VqYPK10QynpV1+OmnNOIGbENjtc5YIuQfVAXoC4ALAtNY3YM070Z8
tsOyVOKJlKvl2H6SdLKnNjtGFZDp11ywtbndZ/gDDztE/ybpryvuIlyeZImMRsFB
XPCzfYrPwFgff3r/O6KwDzXnWbUJ+bDdnIGG9uP8JvzS0OeNsuYXgfoYFKM6PTNk
7Ll1hO5KpsY5wE/fhnub2Jq7D5EXuqeLvZ/mvNFMnUyzhgmHwlhcQMb1JpB4l6SG
L/lPKr76nYxuy6iJGQqy+fTb/3engharza61vklysRBop7JasQOBuIGX7uhy858a
i5He6Oej/FjShOyrurFxKBSQd+oRD4YwpwM5mcBZpnU+S/UipHdH80Tj7/Bxnv+Q
ElK3//DABbZPRkOx6Y7krs5YqmJ8e2T4VKlqqkurOosCKiy8xKv817dyMuemJLDD
1A9UJE5s3xv0YFjCHkFG0S5vhSMYv2tN5dTGau13V+9MjTPWVhsEoB/FAbrXTsSG
goYEzUOg35aY92gV7kCjOmmGGzxIc7US2WM1e29qWZFF1Nz2OPRpIvSF4oCAU2yi
2TGrdQauO5FRolRbUpVdpnxdOSD18zhKH7wGDtK0zPd8GT27Q3sL50PAX30v9Us+
lq700fHkXb0QB8iKuqUzuAZZqceFvJFitbNqQeyEoZrM+7UVtoLHTEDFbTbCf3jp
7ml84/Tz6rYXKYgye5Po9x0Af48CNuu4RxmMw4t1ftzjvxZh8dV3N0lNHDtkFTBn
eo9PWvqGd8oVvVKoCZRn7UPnwEljgSxlWQtF202aePL9A+b/jFj5lrlPiO/zxypT
rJxa4f+oaHIxbWERnlLEEfh7c6tvuHdQuQNhCifbpZZrwkNUMgFJf7b2LoscMHEg
8s5y//CEDYT9ICAI9cwPNdiDkJg4JSMSDexIqN/XtF8SjX9vtNjSyIEsXoI2FLYh
3CoopxBiNjvgYwT5+w3oQ72g3Q04chVOg0zXFH3EoF1Upja8bNkG5F2Axt9iFzv1
PtOcec9D/LJjEyYgcNHUa4DhfxpBjE+WYltXXEjJ0YBA5Gbrs2ThmjoQFR+aZdf4
YnNGCmiIUHF9pMk4Ez6y3DMfDeqJNuD+5f+Ts40KgitRrCLaLYY9alM6swTshisA
ZOGLU3U3hx4sjGNh/DUjuJt3twxuVcWa88tp8+QM+xs00JETOMk4RwSa3EsdCHRa
TNsX94Zx7rQ+sZlOi7IKHctbU7d3PF2utRkcT+V4xWUzvILwDU6WD9C0RYKtkqTr
zMx4nmQh+NZtQCyTvg5nWSKw6f5xD8VWy1EI0I88842OGTJ/cKW4wmxljYK60Aa3
4s6Y0sRfwvazreqICI80cnCbFNIDy+gn9Es5kbVJAFl24BgMQw7tigXKi2w7DqT9
H1bs9BELydMdCov52rNcjcAPQvefsG7vspXcWkahVK4mr6eXWLBPsRLGQbuseCfy
drgNgFDZ4ecEF87oJQDTENehC6ofZ77HcGFfR4Bl3U5qIOdjkoeiNJc/9JKpjxSH
s0JbG4X9wiHxg8+COwRXs8YmCVsJKq1MF6ithd+ZY7iDUDIknQN5DAO1EVyvmSDJ
yXPAkFb59VY1Cg6z3IGZ+rT6Mxl4d7Browx/H1qXkte4LFhRDCg5xTEcTODOmVm0
zcv6EMdyew9QCtf5auJ86ILLtDJGcvDF5NG1ofq7JMMu3GbMiJ37JOEqqmlqjegi
PWY+BLzFShTmf3ZpY9s/pFdeMGda6WeaJtDD2eKOh87HPjwBTA2gph/D1+TiJ4Ei
PIgOA4NeWc3e1+AQNkFh/e+zCnK3hS04erau9/FyVeFPy6J6bizVtBU+LsAmvIqn
1hRMW+iDwyvUfzZUsay3mi4QhQG7vfthzmukRG2wZf0dSSItRRBoBUgDeQsHncfO
CCPDcf1MtQ8oUyz+typ5pCR2Pb7cyGSJGttoAxjqbvbNGrCIa1Q+H0Smcf3fy/ir
pqWO3S6vnKjE5+yphY/cgPvODZHll8+OBR/hMp852SD4mCyebREsr0CAl4n1DmuS
6B8FNWiwnr19ffk6DP1pIYHoLtSNXrGo81wFbykB7gDdsBs7eHSFzDCiX4nC11G+
EYgZg/llhji3ASAcf2mcvpL5WNiDdpkf5bfBmHpUPKDfikBfhwqq8EpMYWs+gC0S
SGTINqm6XlTwWXP5umb7BGB/orbZ5oSt3vFZEpmWb5zx/LzN9PvkLUILYJOdKItQ
6Mo4gL8kyCsRJ23ydfL/kN6Nt6HP6mt6zCGL5GhmKRnbE9JW6nKuOM2tcgn/hoiJ
CtIpZIV7WH5mMmA/rjq/ezgUtoE1IyOwk4cb+oiNpH2rccIp+FmtgyBg4WPQMwV5
3lBKsF3mLcmfKIC4U+6XdZ5gpabAznyV4jDgJ80nxGQ2ceprtjAN7kZ32In01Q/k
DtMvRIS4E2GctrJbhlQQGYXOb2J59WzSH/BeUz0okM9nktubLZkmcYfNQ2cvMeoe
chJneymm1y2mbeWK2dv9JiL45DVvLDk+X+ue8/PUriGpYYQG9jOmNs0c0+FLgizS
X3FEphO7/TC/krJ82VQ+pGIcD9BplGRVvcWHxBXfEsm9K6RjGZue9u5VoU19Kd5t
2lxt8JQSNm8B8NbvUoU4kaUg5kqt6pifKjQDK/RCsRRLXfZTE4kDvYQpzW5Ko2zb
PKKUtTBgMZwrCvfxKtvBlfOjkiwIZFdSfBH+FUFvWdC7s6qrMlffut60nh9dh2r5
Bajf2OTSxyg1ukQ6Xj4hOswIff/fTCA79yEneuF2MF6Xw/VdgH1S1Fwv1JLdXY1P
tr933+F/Fn6U/J1pUjtlCzRbTaxgNzD2yrFZ40CeRJvKtprUIUKdITKWkIsSIVTc
VwzqmMWw29Macdn4w23zMygRhQbteT8Xsh5TMoR8kAAfHu3J3qgc4QnYTb/jaeW/
EzZGyF9oejSWf6O0TwcnAhkfUMwHqHNhXvRSf1mxWP11JwWqerWokgpJ6Qc/mfO0
8HkCRyZK/egDh/AMjQr+tLbudirTq1jyj0sTZT3iN5qLodlOQK2+1wwFba7MR7VY
cm+01eXk7if3EbA7CJQNQ1B24nxB6Uhq3jgZIFLn3pOt6eEdET6tmE0tdAI+sruP
MEu2OuF714qkjLqRvGm3ELHFbdIHRzJTwBPwvM+7L7uDJBLYbC95IRVwa9FOFkBj
urnp6+BCWEYlJpBUBuJSiLH7OeqyQ/nGjAcBBaleTeRbNUV1JeaH4dKMpyER5jrY
YFBaEq0C5rBAnMotXhrUElMTvcdesgah9FtWi0CKN53Vzgu0NyO2aVFxxSLDoYB8
bXogy+2YrfnrWMax/YKCacHN49140gwcMSNyvwnwJEDWAY5c9Li54ftoKUaXd6bc
0I4WQBDw1SKflxSxWXyLADwGMRO81ibvGE4198mA8jM1E6qo9m35y35uye99v1MB
Sa2iHdx8YaTTcrXENExIN8lAVg2Ew4p69sxmwnwOSOrU39RgVDf9m4AqwXmQ25EP
jhVwVrm9cjOa6BM+RqlY8GDt0TQUqvGqUPSB2YvSWMwKN3jPin71HzLNaGmafVpf
gu2LUjwlP59fvPcGWiig9nbUzYMY1BOLNEVS+osgoU9sDA5U/6KKnyfJW0EGr6Wx
uSzfwbX7VJbpewczSaLXlLTOkf7PQK5zHjzARQFzS06F4c/4Xl7pq7PECPrRKNKv
VEhzAta3XZGv4AI6ks8DOZkefNQlTk5INYLQRVHV0GR6TWD/YoqiISdJv/NRBuhi
AnGSydyPxu1kX0ZCb7XDkpsXi2hrp0wj0etV2EgjjI+GEqTsxb8RcyY9RKhgMcHZ
ZHw5cV23Zj1EtS3LJTuKHRT/rT4eQkDRAWpg3DDN1iSMw9T0qS7Bhuon1mv5j6nB
rut9UcFx8bHuSk7TBYqwcj8bDo/zY9kmWMdVOFwgL9J39Baa94ehNYiIgBK7imcv
kaSPrszC3BKIbQez+PgaKl125W+GeCubp9ZoyeUQJqNRzMu6TUAVh4JhK1QRy9Wy
T5kg0IT50cC9kTwZdnZvAutF9VpslMIDtxLgoQV8jIQkT2JrTX+yP6aU83jsWqR6
znhmvwcWc3GbGMqJMZVOarxTupPGIJ+b50KQ76PDSYsqXnDCPWNK3ZH2YFuJmaDt
cj03ap/2uFeWjghnxp6DKMlqiQldZOzkP6QZ6nJ/68EBneBT+5IQRqg4FdnTJ6Yx
3ZTxN0DgAqL/HAAbO2n3oypzpzSHBbAqo+YQ4NLN/VM1jLZ9VCSNHzvTkk1P109j
f7y50L62Proi2zzLI/lavnEq3sSlvbUgscB4IJJNrpts8aue6nEtYlXYSDFK+B1X
QV6lOZYRnHI7JCFt/RrB87P3YNnrTR5WEHcjSeh1lg8N71eAdik/BY8W9shCfet0
QmcikAEOcW7TASErPlcspHtor4CgWdo8B6cMCu0fwPusfP0Xup5HENA3/Uw0MjHk
4QHQ/Dq7hKC2pvMVw9QXBff25FafOsPfVRCH2MI238Ho0OBDtWvNd+yfLedAqm+z
K9tu+lwimHztuOfGdz82B6xz8T5K+9qFKRDONONYBhd6COff1Bsm1UJNSMQc8D+r
EUKshc++K53a11PNQopL0r4MSzHs/nHiHlfXPz9aOWqU9FH6I9VwieeXwOYvFJe4
bbHl1K3xeacxKwS2cCKK8WWeUkzcfe8ehnzVN2RQGuxIe/5Rvu969eTGMsl0hpaJ
UCl5mfPWjKRMTgUm5oJ98sn1giSeGYEhNfbmCM68827XN/CjoIV70GMqP+MMRdNB
4ZDsYIuLUeeYd1ZPaO2fJDfu9miH5s/lO6AhmgqgaPYUmPO0K8wgdkBlOfhCQE6u
b+DeIezh6bekrW9yMpdISOqHhqHYuNE9Ow4OQPJnuRwbxqK0QXLahb0xXcHKVISZ
k1vLFcuGDubkzyhH6g5nmbxQa/HKENyWM+TdJKzYzfPMt81rZOwQsbOfWRTn8btw
XggPIZ4ftmEDNCfGILAfVKYHSQg1cQgwHDG131xXDIHlXFWAo0nEGDd3l4IXSgCa
ZN1XLdmK4jUftMTjMWSUrLRijIgNjAwHRfTUGQtA2gowx/enYTXfCeRgahRCKidh
EPwV5gP9+dRoskjNqjZQDGlHLf/aFzOlz5qlABMEqQxV8NqKf3SOL/0OXR16fruH
MDM5PxwHIafHqBVoYH46bd38lTfDfJyGzKZxRiDq50762+jcjqBNHOdTSx1hCb1B
onNMk2anT83v9lTLRwFgaWGXNxE7yI7U69OPvCrwcfFswX2mo9caAvwaFbc8eV2q
iCeztpc2kRGbglDwyDDVSvAifLxBeuuay7aKqbKs/aZZ7guGMhrncE+FW22CsfG4
bt8yTS1DXxo94B4gRDDFg3B5fEvmKvuSgacdfvHhTCCEmgYVoxNiocRTToRjT7hh
qoO+NxmSsNpGXZcdk9Bjdhpzzm1zU/N1OVHMV1cLdY5syXsweitWvzaObpp/ipb9
UPMeA/ur7Z2psAVeTCpqRNxe2YcveTQPvQ5KX13UAkskwZf9dxstnuxg4pttLMz9
AG8ZsSsnsOqTbR3XGO9LaQdp9lxk5hVcu9AOADTVBqZCHDNIAySdgnUne9iAyVez
QqpM3IjEg9yH/RqQH+xYUBGJg8btEkIg4/9LBMhNQ8WTVOK5iw1yzdY+pof/SBLT
gCU0CESYLwWIzMl4OKAC/5GO4TxVvCMDKxNi5ie3k5Sdmzsavo6mTI+GJcnyolDL
CCpjr/Yqavbthyh5wIgEYeLMucifzbM8ltR807tAWppH3ztuSuZObalhnEthUcMg
LQOFiocxw1Kx4wfO4iWOG5YxNJQjBI0qajxMbOBZ+1g9RJtpjuWBIg5YeQFnkVmN
7HorFtmhtSDgl1WC0/A8q75B+blYxSRT/PCh9PssMLI6PXMCCF1d8DJXN9xyMvrp
wFt0oj7JocYjs29sx2HTLHXZPj8FF458800AoJP5N/5giTfYZk2R4fqh+6B7JliY
nHNXhdkdqOVxjt9Fq7HAPSr9OgpDtZNCvbujvkZKtwEhk9oZrA6yJvPGsLuWqRRe
YnKMS46krA/65ShxOFDUsSdSYYCmpwR2MwNyB8QWpHrm9vMiAIW/vPKWYx4Q8M8A
o27p6tu+BaMSR+1Y5kbTtgdrwjKEql2oYVdnLvnzgAxgeVVlvCtF3QZpEXFQJBnP
fVl7dXzhxwm9IGBVKXRFhes2m/MFX7lVaizg/8GX55PD2jrbCmMMOznRYZbjP5R5
5koKCrAUDbhFSELXwUAWj4DrzsDQYz3zF3NDnvy8KtimmNEe4yboryNszEClbKiq
D3Jpj4QKjyF+8XKNWCxpS9pzhAoUCxW3H1OOdw7lvhBvCB17V8z1d7j7VKf/SmYT
8/U4b1tk1OcDbuQU57eFlOHWA8qjqLkAMuUOMEaPZF6XGx1+kRAKDI8kTvmBLFL0
s6vnY0aOBrSQQUlIV/0nohXKyWC3+1rU0VTdKGtar3e4NReVLYOM5WTe8PaJ8BAb
8Yl5YbQveS9FidUy/1zqLMb7dyFTViGGlO5pr4lyEUh33hEToBaZ1C+yBQ1fx0+Y
3S2Pd0n+9iKLUF26WaqEWtZiBw90aNIEMLWjBplYDpJRTRTzw58RmJ4FVGKWr7UH
ApxXRuJA1sy8+4p7apQ29y3A9O4R2c7i5dwbgeKXbzjhxgPIvA+XidikkD07Z/b4
ffGpuNt13ualIqOJpAce8JM6aQChFVcUSZJwTbFhGqZ1oievyHgRBgCOPvulEliS
JkvEVPJ6E0VVqJl2VJ81SkKp09ZGaNz7PgjCNfUrYfKYMv3fhFE80pE+SWsFTWi3
KG4tgGTOXQTDC5m6kCu+hGYGR7LZZWSbGgUxIlR79PBL2mFwsuAS5/A8217/vXMN
cEiXLTvXvuow9Yb0mv1cRXQo91CR2LpSlfH5YuoBiCK2UShD9+Lyqjv1ydGp22Ah
DxLCLueonoiYBnEgDpdVKgeN8xJAMYBkkJMcXbzSSjXxeD3sSOFx6InP9A+cWARC
x9X6rIVEoyKVmub+sBbEICegQc8cx8t322KQva65rcvPv3bpuh1WMuI9/jPYHizY
vx/ppO24RGHtUvuf+/e856CaJSrzbCuMvE/zz5WVKMXO7meIlXyCjjY8+H9tzs1E
T3t2AahrPw4my6L7zpnNhw8S2oAZuXLs1wYLN9XyAoYIuvWtKI6YAl9uMUw2DEO/
GUgUTtkHK0fcoGZ4ZDR8+LGWZsD+Rjlj6NgDPdtxUlH1G2OhbBLzPAfJSyi6wckR
8Kku5U9C8Izv/AVijR83cTj6RpQKrbJdL6PlVbHkhBvhCC4Hb4lNbA+yqOQdvCxR
aSnhQx2x+Sh8kN20w3BZLWIiL8G+NaedC0Q/WWs+9OW0fQaNPuvqgkVG9ui5LqM5
daqJFPBMgkmDtB4M5tQXlvnTrsAY4i8gPRc8yYroYGGWgHqHeVLooEhwTeb/p5sW
eKRBLKxasEDBdjgGfSa0GO1nlN/RaTj3g6iB9AmFSgXI1LCJfc821+YQZ/M/jMfd
+sPHSyPcHU/miYxUtmxQ5Dnv1+LeVHCr11LrgeiJpx36HMv1tJxG97od7kTYSwWT
kTaucr97U41QuKANt4k9YgykDGcOkUftduCvV8ksep4ee4LcqhysRn6ko2kNHwiZ
9nvHWkEWT2IURe+3cncGeAd7gGaXPiqP+imLdIXV6VjfHfPJKkGvJzTZNtfg1WcH
RupiYksOGYm6tCD5ChEilcIaM1q2e0wIO2gyvxoOp9MD0NLmqgTz3zlGR8ikNqPH
N9MWkwV9LCGbMb1KxjNRrPN0zCrFagZqylYIK1gmby5NzbvHNtdJvwx7hDYxE+j0
UVAghaWFrvTyZJAqgqBDJ5nMtuLmRmOkwTUA7OMJC2Cx4+quXre8h6//ZDoF0TqA
OneRnG+R9XG/gdZEYeSC6K1fgm6H0jsUqe057KLE/0GvBriXgZeWBjn+hyHmyURG
/WimYBSYX3yay8ZuS8KONTm2KQXDf6mAJOSu+TlOriY7ILZ0V2Cv7jJycjdLY01y
QwIFNs3RH9kNZC9vYQhFXpy8YmQO30qhnlq5Ys1M9YOeftu3vR9SM7QKkadwGawN
aiLk0ww/9ZzKrNN5WbpS11C63QXB4EpWDst1k07FerbWm62AxdzqcYecDN5kLhUC
72N7a2mP6PX0IWGYQsjBjgZJ3FvCtjwmUe99WoDP3ZmVWQs+YRW69upghG1ERiF5
Zd85lRsC0s7VE+W2heDKcOzeVkGZy9oTXCvfVj2qGMIkV/459vURqlMkTBFTjsmF
J4DT67hs5O6QqTrZfIvxThsWNEampQkKi/VKT6TlJwjsXfd10kPi3YhZYLU2IXw7
KtuSxDsSEt7cqQ44LAshszLb8fa1uHSyJya31ZCT/nfcpP/BjDSWsBRTw0yOBqVI
IwKJ+qA9EoBQXb8t1QvH37GZN6XK6v6L4l0RgTAMj8KOw96V3p5FiQ7CbKNPcbd1
EI9pRViyf+ZRXHAczvzKtOS0oHS5uTEPUpfnhljBkp1eXa84O8pLz2QdOKYYFOxV
pTr93q65+5HUw0xvOeiedzcwVw5iHPDArDZLPxnkEnxXl4WOqUoghouphvFTemYb
4DXfepzWlOMdfUlmfIrXXP9aKNoIoohzB2QExyPEce7nKyrN307RnaKdq5hgEmeD
Qk9kbWI8V/AsamBh9yxGcNmqNrN/RfQYfFbMyZ57I/NxhQZy3kNHGCkAygfsp1hh
aIkJuCfBn4xkL/weJHorQ4rcpf9JzMBvuLI9UX8MWxDk2+IYSjX2yeHqNpLQLpTz
Fpsj/6wQNPqWTXCVAerzDWyeksb5b1mEtFmpPpN1Um/03P9eAJJMlsQj4kVYNfDZ
3kmsHblTfuw3TSMFXjxBYVLmnTFBfp31JbP0yTlUEN1HbHDmOrykcBQHVmMxlZQH
4wEbwHLfMpee2vfqQzOTeoYlOeEwLKp96rXgdsYkgCpWaH5ri0F1reMBccJGCHzv
DeVX1VgqcwH2WrOvXzbsoPEvvxdRxJl3lrn4EM97bswxEUU1KxX7C+gihX/G3jyX
jmTA33Uo0vg9mWgx1LUA4DP+lpqzaPFIkaZEzhE7OA6GP77RZdA3HBzM3Qn+IgI1
0UQRwJZk0dc/2z8H8gAtjnMTln8GSQbAYUoHNKg+c1GGu1X5es+nSbWPUMEO9omg
tLU+TM8iDvpLn+0sfkwuACqTEG30A5mMHjsAUq5r2N2kZLx1dlpugNZE0MYVN/+l
aPXjhieTvLLYLy3flD1neEehIas53700+UXOUCDnkUeNck1FIRwINThCINZ2WuGQ
bpYAVgLC0RomY1CRk9gJs3Geq81WYpqp+qq78Q0s2bsHDzAgdvvv1hhMv8ORirF1
23EMTxk9Yhln/KvYUiYN0xgghjl12MTwgCQgq5Eo6CblBE236AyUYbghHXgoIspC
wuq3a4LSw8TUnYsH2YRGIJhMQw+PhDfpr996JBBtLV4uGVzFXmegjW3lWqqwOX8G
1yNmyEhK6LC6KfgsOz8fEAom9OCgkMxQx9oBAlcyBWZUWyPfq/P5TE5JMl78eSdY
UnpgsFzJM1kJemOOng68EmCYJtzERxMhKislcNEUhq4znUDE3tP5DrrIASTubFDy
l1DFv6P0BQS/02N6vz8Rw6n9BmG2ZL1UeE5KBEWr4G+tg9Zfy0P+qvF14NjZmSTT
+qiBwGAjt0svdyOHsF4eBCUgugqrcUkJijWeU4ytBsndC+BxdJuBOcVdNN8lofaz
WSCS1rPmDbtGxUQpqfmzFXfAb7guPOepXOUxR9wZi97SYhWkm/B6EeM5lSpSOiht
dpXa6ttH64Tbf6frJtRhFIivpvJIYzqnX01de3Rcbsx5Aet18NkwbgMnNFSqUUmk
SzTFEdnwRGZAg5n5TFNtGG4mwMZkUmo/+/gx49YAOK+rU67J8f3XkhT7rQQqujlp
w80x15v0DIw0asbY0YsQ0G4CpYF33Cjz25rMtASLKFqgR8eruBYC6Uuwbnhumv4T
17dbnmGPHc1mcYuNwN+3SSCMVH62lYK3H/7zMrvD6Lyl4p3WFhzS3IeVJLOvAEiW
W9TSv9mKlpI0GhtKXKz9KBM8CtdG5ZNMejK2WEI8pcJ0/g4pKmqVwzLRoS9EMOa5
34Jnc4lXKCSjYgNFSXtmGdO7Q3QAAwAr2+Drb5qR+VXXMhe4UDt1bGcTH3hBlZLo
dPBt6GCxQBrDTmEJsAKU0tl/JHkmNMiGDbFgjgx3xMMEWreKdkU6TnRqtf+QBSKq
hYDNhUUZlLUPkZtuVhpvPhQri32hhWtf2hDmbjYfJAQQVDzqte5uVZWheeJ3Fp8R
MLQvqunU2pjgtzIGg7guqjSwyue5rrM/wEl1quc181iji4rizuK1bEy4uu1kZjwz
fIARy0lE0qdCZbEEftS9xo86ZA22NxA0NUvtMMcWyWL+ccIe4lihjYzzUO/kdGcD
9olbx+csDUYKDHgqMBs0kTbheRfYmSK9PsZVV38HXGPj8+IMCsv5K4RrbIfujayp
eo699Wl6kyWZTMpphrVM9H0hhi2sZ/0n2xJwzasekAwlRfoyGcp5Z/7cjWuTuEhJ
91O5D0wrjRBNeByyNM3wJ/NahTUzby8FUHzvxTMjCksJjHUDu+rOjFlTBW46tpMV
QL/BoDCNx+DRX/8nBEoQ2YgQYBgvtB9g1wmXxpoaJMXXWlQP6Oabqv9k4Ld+q11a
fnOwkF2hXhVE0FgYaBb2/YHYRmOSOSRip9Ez6coFb+MWC5nX443SPb9XOqB7ScJ9
U3LcrYU4vyIZZUTR4e1jOw1eJTvDyxUA1sOSGOB2xc9iTVmAiO0gMuUBTsR9mi5J
sinSjGeCY+Tmi9JffQsHnNUOeVBG2s+en8+uvROJdlpyv0SlvYHl0o1NAz3PFBnK
mxe0B0ErnKo3/GBE9aIX1cyG/p2Coqy9O7YuyT7Xcf33WXytmJukrnG4Wz1cGShv
GFf8AM2pvTx0tfb37QTthOxQjbnPzKZU+cSEQn3qdx67J9Vw2RuZ+DuYU3CSzSqa
OqXJQX3rkcVjtI5q9b1bgYwiTn/SEyWs5BWK/247qoj3fQ6+dzMCxcwT6UuZ/Z3W
7xgvb9OLydqX3UBU68UbNP1VDK1V4xIUdkePBxOT+yWgCsS8x5NciZvd6Zt4aHyv
jkY62k5n1yoKhha5301oy2R6WUTs8V2tQ2QHBfGevhXsxt+9Ea7cnVE6Ggrq/KIR
+cLfbssyws1UsoayMaL/+8s5dy6uXm2y0NzW65ZBnqUmveujW7CI5R6t8foQsbt0
kufCFd5GxvC3Cqmij3ps6eiLS5zov1SZNEV9jetuVYGMKGqUU4RQU264yNZJYB1X
GYQZQFTDV4v8nGyJ6jgkdBT8umsteMQ593uYqnJ93HN2GXI02iFt9mDcJCQ1T7IB
XoEqRmL3+vCdOM5sXUjz2f3iu9Rwd2HbOcmOvgUzfikP/l0AbOtvJZ4mWoe7hTXA
PRZHSxHqEAdT9iULR4SV0BwRxfPB8b2IfvRKp8mRh4R7E96Pbtq8rAR8JntuviKS
MeX1eksm3J4/cOYFSl7fX4p2jmNdoFqsHskfcuM0rQIZGHeoTbVP1ZYTea7nRmUa
xszU4WU4ZVyOAf/icXKS9JbOM0ggiaZjnECjAyLfoQXefxu7jj8CgJwlrn4W5mnE
5oep8HNQzWlCcOd6wPV0hnUvB5YH/ehn56bGW+nc9PRcOCFtmWxuEYN6OUaRuGMQ
/H8boJF5tA8BzAeszEOpAlOi1hPZvmCDeQ+toF2BBHr5aVlC7nY9tr7ce66mP8Iv
eWACnkJEdnBPZ1MkkoTGwuZdEq9RbILCMMBSUoNia1nIg5oSLgU2WhkO8mRskOqW
iUUrHSIbMY4sYivfSBAtbEbqjZZM0sRusuTOLFkTPCTlHH7NGlQPhIB3wgVIBuze
n6Ytb72bfOcdsEBTo/Su6mCPjjdXJ8qibl1iW2LHbw7OxBY7buKO3ttCGHiTWHXj
/TYQar4r1VOt7uC6wgZ1bDTrf2FXvRVb7iBpwnxz3wOS4Z+X9/DilowP8BxZdwMG
JLl6dOpY4LxtEPOoxutwxamkk4I+lNObf1mA95wMJW2EmAJnqR/E+7aHqzcKjDSG
DxeXb1YkJFuWUYLng7XEez9YMwwFf2LAM2288zYKy1GZSgO8QYIsmEwQ9bkFDmTn
W4OqAYGh8byRK5M8VxL250By+h2YKc3yherG4rf2Pr/GBbc8geUpUomfSWK5OYt8
SmrVUpcSR3LpcD/Qk40WoHOnGupZ2q8jQBtKw2s3HRPtjnlIfM1GqnV8X2LH0T6+
70SAYzljxl3Yao3Pil6s5wDNgFBLBOwQ4EK5cHA7YMHwMQ1YYVGX9XEctvEKyoG4
NCUemMmhH5oKg+5YiOgfaYtqa4U01T8toGSlpugKOdjAMBCkX7efTM6bW6gYrXir
UqanPzio/e/MVvxxmRGzmd+pia6L81sdiJzqtiCGziIWWlAkNBcGUoIYEc7vDgXf
Vslqh/Hndjd5bFXfMr3F6uzMtz8KLbtpE4/EgUE7NzGKqaWp5Cvs19wWTeXIhzB3
LTK1ZYFSh/MTBvJhYdOnwxl0XrEK9LIvJ+aH6Nb1ROxHmFPVJDgx2qg51CFNugV2
D1sULUpApbPscu/2Aq7JZR8eX6OsSaD86nBTzbp77ye8SDDDKEpGEAh5oyUhM3F+
exs5BWJY4Gn8QQwQFIqQx100qkXwtjA0TobAL9CxFqLcL9F9wj73e+g/RC73tFim
e8urCNxKcPqaXMm//3tcBZ2zeEs7P4XlZVonFt317DApeLRgh7yWoHzfEvb55Mqw
8/vg/WOK7y8FFdfw0+HHyBgPNGLjJGm5hnhDIpJrtakTpiPNsWa/weE3T7TiXqUN
32bQ52ya9/ZF3OVwKGGo+bQXzoGRXJApKjk4FX1W0PTrTqabE03/exdAgA00Fby9
NfeIWHSn/bFANwlqcj+Wx12OzM4BcVYBfOFWLxYoeneQczcR7uZMKvy/Jl9NQMSc
kMQwQsZBeQ8DTlJn7zSn84JVrzJgtobup9HbmAGqbDkB8/j8PhLjjaLsooNjcUV+
DFJsOdOuMhY7d7Bvii2G4sB82+ZkxOOxL2HmRMIC9UXHmHjpnm2gD9hn9VJb4Yxz
Et9otlG4UgvWTFNQ+fWe+JgSxSFqX8ZlNVcnax8rywTcIvJi/CmacPdkbn/1GZPe
Ac7MUoOwcOVKsjiHdBaejYIodzCiqqz+6fP9VoiCs8wNgc/ysILoN/FMZksVBG/3
qal+KvskO4sItbd2xwpFk4/LwWsfl/w3kWUvu12vgc/tRoyCef7B2tfUwPWy4ov+
bOPddcy0yM9GS+0EAWFGBG5j+MXpp7BBfQ3pdTkUBWHRt1AK0G7Z6yxC+rWTozBH
8pQogTaqg2pTflYKJzhx2rRg0U4Qm+UaVBvQU2jUhOycTZkiSzKVvpgXGvBiDBeL
5Hs6pwbhHwsD1CNFthF+ImHoef2E8r0tdhITqoUkBNW3d0TDBF4wE4+KEEGZ9dse
D9QFwOaLd31ke2bc78ppSci/iZISka+sMAYpHlR4NgYI2TxJeq5Kc5yGixW3MSRs
ta/PiS5W3EkYnuKZCLbq9whx4vnywT0C6BkXUegb6h2j1eyYMOlT/22tvz5+CIjx
LPwF4qWXrdvcXroKPg4QorPEO0S0YVkjSQ2WhTYEufyWOTkUjynNZbskCQlWwwq9
/pS3oE2+qsUkwhKSKKBQLaMxHUeaIyC39qlVq92byFa+pThESGynlTeIohnmMrYR
u92boCXyAahTSZE/1NusamTfKXJ5od5eSuLoUn1U9S6t8Qwwmv8Z0SZYJPNMHA/Q
h2i9BVlPbzBX1mCGv4fUnyb8OkT0t5A1QYILFYcEy6dDEur7vNhL2JeARxli7tzj
t9JW3fdzfcaN9yKuk2A7bC6bnSRrQTuSJ9zA6OZBu5OYNIzvqEwU3vUr4Gw2StFS
SKClAYAyGaUIUApYar8SGPC+ilKh6eW3jCg4Brudizquzc0S6fvb33dTm2Ws1WFb
TVPliLVsJ0ItDZI5W/66nOTO4KKcPyQ/bwohNBfpxFNBSq5X1oCOLGUNs02r6Ok+
ZD2VLS8qR6OmGUQborCVTTT+dYOOdoT/wNTM/MffIuF+8598qRukNv72+Ax/KK5+
T7tz9huJbP+Sph/UHHSfb6/eZ4EcNQnDgUpWUopsWpPBmv887b3kTdAjx6m/9aiJ
FZ5RqajGooIPzSSYcELewLA6pvMH8h9LSqZRC2rJj32K1nJAZDf+fCV/t957S3O0
egdVD1rCTBwB4ZMjPJDVAjX6G2XP2bCW25tGcUi0f7+1pQILPvlmW+5dTms6BnSM
vbGapHiwmUAD+0FEo9Xx/2i6eKurSiAPEUEO+5K04GhgkGy1lJZ+4jlBpaz+u9sY
k1LNV1+JxUgR4sM6gqpCLGQ/RGvu3gEWIfjzDQOnsMdPwUbVWxfB2UY1bOqZaweD
LTqdak29vAJEc0gDwWmaLfO+oXap9tEosq68MDlPev3zZ29nJzd2TqsPnqUncvss
UxbCQQU1ImDTW4j5dBZobV2ajQeakQUmrtUt0MKwDHh/htBap/py5rbX3JO3cNfw
kI0T7qnlOet2CeovVMbT1debxU0zalMNq8McrI+esxl2xs4IsHKpGYnbfmwn3Zcm
3qTHPUeJg6HPA52QDPKMHMzmRUR0TcdJaxzK+YG+JOtOJAH33Au51etTzAGcgvP1
6Nh0PJl493zLqqbk4MKqYS7sHqCVRuSHjiDf5Wnkj45Lccm8XxlgPs40ZFkHZIaL
oxFDkzG64Aq50Gf1uJqnKDS/t37HtwP9fb2bAgrM675aXLevh0w5fL1vKGexCTEP
TrHEighgC6gp3Csi7aWWu5B1cvR6Nj+S9fufU5O9e1+0ltiYuWTh8l1hgm2MkFlu
5Ts0O3suWzIblW426zeh2pdOUfLpLZOFkee4ILknXQsRiuv1c3afIGo+sikD7cUT
5Yy9JIQeCDHXbK1brGgIzPzxtJZXYGXttbINPIA46Y0scpTYeZjosHakXsvrBCDg
8JiI+objoWXpbCQbdVorYt5bQT311Lt7pq+fbfzS7uB0PJ1aVN4+gY2iNpS4wOUN
KiTV9T8tjryBRTLAaG2eSQS+RS1rJ5MNoWvQ5X7hcYFVf6Sw0JMqCMicU7T8+qnD
6e8VU4ebdSvTcPP1FGySnX/+dkkr4iXgEjmZphJC3fozCGJi2O8IMfXRN0WNqZXT
+TaU5YSZy+zvGLGaeuuvcGQJcTbrtReb/e7usUIpXlGMxigfsCxrT7E41kDznkKB
l0xIsn8WjkXGpTsuOES0R5ff5Gwjcc2nFZfABCnrplOCmklImlNVszeZUJJNazaC
Iqo+cGGHaZikUhUpriWid+GfVUS7d/vxIHA3TTJQuSzNM0iKzSNv4DT1OwieZzHw
3RTFVDceF9c3zc7cEWwojm0SEpRKVoawzz9CGq91daS9+RZsSaeymihVn41cYpz8
2nuFiGT1b89VaK4a6DcKab0ucdUGbYh7wH9ukgGMJw5zKow3oPJkfU0Qoz34yIQD
OqFweAMwX/jkJAGlGRDA/RPagmC6HdXqFoonTgnmNydAx0/Z0LibErJLOEj7izIB
7CHoYfGZeM+xvtXaObfq/Vkis/ZzJKCGn2o4AJtJEe3fZiPvhDDGYYx2beAJH6m5
cqAiy6apxQkP+E/1HAi587EBlzpxfB/0Idm/PxNJzaRMajkCdyrBCDd174kNF4UP
of+l8OxwxVWEg6ghngzPx0nNjPVkDh4Xdypu+sbX+ZcpC5yV6SjrUZ8ZHsouIyZv
2zTlQMZ2m59b6JgqABBiv6CN7V5j55z3YLnH5qhIvm5d71kuEoGL3oG6aOAv0J5P
IxEZZDHzZu+GAa+EhoDm56R98/WBs4ra3+A9pO0MRWfJZQPdj0dsDymW+Qvasksx
P4Mp2OUp24uGDyJrxQh1LrwzM88IqcvHKPVlu2cqA0O9UoLFCNf8FaQRmyCGp2bT
5JGcqMrUz0DdokX2KcQ6O5EGOD0eqQnYoNp8z++U5m5l+KnduMAMdyZVlx/AGSGa
61YRW/g15naX2elsk/wJDhAu4A2ns4RpPMFMk6TH/rtqMyQNcWk/44M1ptAnMTKz
KvSBnyvJjnnrnscZUgejJkEIWuzNmwYtzx41fw+9JKlZJQr1XUFl3lqb6XYWA2pv
WHtVhAb+Sk67T2bQ62f/0kyf0pZig9qOB655NaJpju2VhAxTcJyfLy2XzJf+4x2v
dkRVB1jw+zbztiTBEJtg0EPiufPbx5zXYBXG0jBsaO3evfK42DyTLj+1b6w3jc0L
FOnaON/yv+9dSIK0iu4zl80Fhi7rB/HxHrGy+n7rXxJnDjJatf4npWZkGF0Vqrnf
pOFFhjsK0+Q6ZhbZuI18MUKyuYgSlvd+QtivmWb6pKNjNpJAjtP8ndWuZjbip3k5
cPo91bhqaXbP0OmtBrUc9HJpnC+qIrJXerx9gH4DDymlm21anPJLekchYU8TiyrV
ebaNwtycZqFi+MmDaUcAOrmGzuWu7Fuos9ysxDm4zTMl6znzt5TuDO4ODn+2nZE3
oPUf2I0EEp9ErrYOqHyh/vk/9fa/28hw7DN16bIQ5hdzXas4lJLtuqbqfjzPR8P/
BE/FDb1QuEOtvKkDvK+Q32FTlWQeTHyYttU2tq7PgKxU5XKF8SDkwCGYfr9KyW67
8u0NcvYiENZc69uknj/cdhUZ24WlPChfjX3wxYnk9JBPcmBwr4slf1FrxYCLqLDe
KjYzFfBJqkqE8flR6dqq8Kq0igVnCfF2qZ2zglky6WETVVr49PMcIUd1hVKOTYG0
HPLOouVrDEgYQOXUew+Uoe7MsrYKjoFu4YfqVCmlhmqTzhq7w6+YRtb7jYkO0ibr
u/oGu8iLjXSJl9HYHAHWScXTVLAM83DH2lY7oSkWdKUeAgkOwfmkUgJQ+gGeMerk
+pqLrn+Fepfv0hGdHexKB5aA0WZ4lYdYqUpDeRRyZGVbCrPjqGveQvcGUFgp47Gy
O/AkmNZ7l5lnLlq7Z8xFsRfFemdAWEfv3VrYs1FTyB/G4WRT4Ajy6BJyuD4HLngE
PjZTE9t5k+d74kIR3CPtNqlMRo1IdqBHs0zRF4i1DNXCKJSBcqtKVUItrS7xqE8I
h7vZY7YZFDo65zfE5/xdbBX5o58f86duOI9nUsSzZeaPppq/jGQhaED+EUo/JCrS
7W+SMisVWD2Qy/E1P6Hg3M1nLX5dfvA3gdZDQK8j/V+uaX7sj/eHR76DVmPIh7kY
U+SJMJunQWWmiwZBzUrpdqZ33O4GkoDQvo/IOUY9hkjQZk1NilEgJCBsfmX/gUoo
vWNdfijU77xFsdWVxSAVkNFVs6/OtWd0bkG/VAu3v8ha3OJXmBlcg+tcEwAA+n0b
wyWCK7hicj673ZOAmuR0/h+zksJDLyPcXs8pDC/0RQZLNWCb3tvQP8Ap0fyJJWNr
h9CmfswdfK2I2iEgIrhFYN48W1g7X8NeE2SFLUvWhMFdCNU725mzgB5FjAUhFOdc
ad5Gwr5B6YH/2lB424jwfDr6SUe4HgR+A2al4Wt5CMeYa7U4qDEgphrTGXmgCt18
KIPiAFTG+Y9BhlOGC5qNfSydqAjQmHNOBCyuA36rjNxdE8E0bOoyOmg/aXl3dfkm
5lyHeQTyvOJDLu++R/ezr8QdCXzfO3k+s+QdPqGd1na27EYO7AVE0MLmo+M9bnBn
ctt49ouinvwXrD6eX2blpI9he7IZ9i1Txb5sycfldOcTGbyY4eUjY1puDv/doqF7
nfAtzP+NsVKqCBRbnvsw+bwz9PgsYsdaM8xXE/4Z1wy2P7sJwiLwGQMVA0T0N2km
hZn0mVhE/E7W7vrbLxThHtuU4UOixcl/KAVpmHfS6BmlA2ZcSdm21O7QdK5kUhw4
3cMNUvrYGU/K3PAetFoK8Ap2/C+NmFo6+r5FgqmLqnxbKLkl9Sg7CKRopY/xNzbN
qFI0BTBjvU7fdHUatN46VPCmN60ZH/NJzEGFKNG5bLrJjJ4oARu3zEL2CL4iN7NV
mtzjJp5wetgk7DygEg2qT59fbtEhCLtBoxbhywUdgb4sYfX7330XB3pDLBK2FE21
41q5syj39GGtu6rlLBYufE1aVrr5cIQgIWCxGCqUOWT0j4Z5FdzPdIYzoiW6O5Xl
ItCawhMxPcIZ+HPbmj4NZUbF1QbSPneeou+Sa03slqW+IqHfnGi4iBPKOpVVOx9j
8DlbQ/mIHMhWniSTIMHRxlqNI7+kz32Y97crBJR0H0sN7N9xrCVktsfV09XViYE7
YpmvXethJ1X+CHbmmXi/orVDvJYAuc+chOxqTkjA8kgEP1NYGpFuj2fXnGPvTzz4
pYyOJIURBQW9RnyJIygZ/VcIbD95qTxxMr3/cjxJOS8SjAw4EflQRCn4+hA8RveW
MD6j/AfqgLOzO4pQFjvhE9y6CzImQAZPvn0ugQytTWVcCG4QngddOA2KClvSt5fr
OOGR7QCL34MbmYTGAUhKPZCFyZYiAo96ak4RUjwMxGsoAQbDi5d7+tnLxfcT1Duy
MiD/zlM3/y+LM7IjTL+CQtwVOofh7k2BGxITICU8Boq8Y3OVnD4WJV9BBvzVJaS1
NOqAARodrZubRg+8fHAvWKrsAWoMauOeTygQLL0tkl5Gcx3N7IIaKUVAj7tUwtlj
EgjcGeHp0Tp/B7fBWIQNw/I2JDP3QpTGvjDqJ35+F0PFcatkBN6bYW7cJ5kns6tB
dNjDdtmeVP+2dlp4T+YJU63Wj6gwK3kcYUxm9yTReGATNacgH8MlwO5ra2TKL3mw
4Id5U2PSu6VdfqKyUoX7UURLB6iDLZzo6ZLanGyK52y68ggk9YfG7qSpotDN5kUJ
4z+Pzj5pjFmgWXl1canlXRoFXMcxkniXXyM20ss0ANIi/yT8Hfwn//lqUIgMcoYy
fttIqs3s59JkXROSuYjOcFDnjbqP4nLmylMc8mS3DT/WPF9uoBP6Cqs5U6ZDmkhw
2r/F5I/lvGmonRQJmC/ANEjRodYqE25DFLN7m4ffnv6W4K1LKbariQeGr4HQ8871
gzUqdCpstDDFu+qIoFqJ/eI0POtFtYZv+aEySn63avnRG7LviK26u4or0pEtx6aM
pTbHfo0ducbHVAThk7Mxn99Rq9qT6OKPs5ivZNTOTRIbL7CPt/rtY6WuE05Y6Qq2
jGXvZTH3/0m1+T48Wl+kk457fSvz42NGe7tUgSIViVeCtRUaS+fHhckOgVcNfeCj
D2Vdq05YHR0Iv6nFd1NQT2GD5T3+OW6+nPSsWLDk/vOSPob+D1wZr8eaSVyEP7K1
lQGSh2Pxwc8520xvjaftP3386OEPPm9bEzTtObfMNdxB1w3H+hcz0wDX5rg32WTI
zKWgXCKkNYYHHY+XcQJuqSS/Lx1x+db/E2WKPLEcxt1iC3026KU52WtR2c6B9mW6
BjOs+OpjA0uy734WHqg0PvRpgZXSmWvVqD93QWKEINdfY++aVrVr5wRbGbApgZ3v
NE6T3Djt1kbihfQ/muGA0b6OcnMO0f/JrCqyOEUQQdcMDJqLEXjzBI2IdhDGtJn3
Bz8T1hVGD23QLTu2nBVMG03lTcmvBPXRedDjANX5oPjursiJAZtHKfEzfo+c0j5o
9D1VVtzGojirJaDMPfXdnfqzW//8EWJFn5ZP97j3uAOzkhWsiAGqRPBYtSc7OtcY
fukzl1F+0o6lW1sjkQW3tR1Zf+eskdTCTV9a0YE9WYTsR2yILpzpTh5ZfFHzZ7YF
yOyf/SEM+l4e4nb8uFonofwEoSpQMtDpffMfesGPzfuEtqlDxnyKP0pyfG+g5EtL
ssee1jHMZDFREifU2iRqVHsGcnF55OX/rEF7s7kI2xD8uh95NuNzh2VzFMEg68Hm
CixU4LjBnUb/oau8Iiu5UES6tvj6lGDAbQtHiKz+baq/lSj4EEbb8hAruY0PcHax
0NnWx9HxYdM/Aw0tnRZFj3K7+ADh6cWpMR8zbyR8Jcf+IwuTgGg/5ORXFf+Gep2W
PJGRamxonb7Aqfm5Zj+6QoN33iD9Hd6RvTRrErA5z+JiurWVorLEOlWqw6y5lE1+
Nm36gGvrwJ/SMd/dZBHswdfiM9WCw5ETbWnf+nptHaDUZDAp+V1jxIpoGw9w2Lxv
3XEBY3CY0Kh8eIi5xrzUiPPJ+lIb9ts9bq7CtnAAAhIF26HSWzgto/CJE9MEx1pX
4tkJqZ+fupp1iPfGb0WbumujfAgWlPemFAeTt2gTwN/8rXEH9BzEP2hnjJASOE9g
jSmGSvrk0fLteRloe7oIWWhPxcjwNojLjQ4zI6qkxyWFzwSg6xyY6hiIOPoFHr+y
Q0qJKozShH2oWVRbD73fyV//qxC4AgRdIOcNzKRk9jreIu1lqPjNjbdtY184DiEa
RptWs1oflc0pTJdrNnAaBem+kc6m/PVexaC17s25vizUTi/vSrb0IvV1bMy7jQij
A46Vk8Bg7oszobWU1pNjE7yNFmDtxSrkNeuaZacoqJ8S0o8lYbdaKvBx+FAw/boO
F7+0Gxfl+DcI7h5UI47cbmFbiQ5HPuVtR4B/PlHyVN5yT+3V3k5+Jp6qtW3VcCVz
4nqN+w6TYMqEhThJ/Z4pbwqkeT6ZLcmgGPb0PVcQNSYeOmYlQqf3itZVxX83m/Tc
gFLM3DlpoVQmHJtCb61B6edequR26aPzxCIUHmedWG0ga3pjdxrMJcvp+vZbymkf
etgVyyt+3C6m4Mpq3m2/j5ayBkCNCct9+Gt0m4dsuh+t0PsTPE4Nr2yNh7fgF8hB
xRWjRSfv9z2E+vdiA2j1ngE5bGzm9mFERmdUjD/QoGTszFmBHGwI1z+4p7CGOLrg
A3tDGuKY662bEh3HHNdTJ4xPKxDRODETOcdsXo+uZWWKZIEeFDGdMzqC+78VK0xd
q0h1OYERsdYToIrzaNiwZ4/T/dUVjkMvtXdpdw9blZYy6DUuGXK/AcEhFvPophQy
ohXvMbK840B6eMPvouJM3JZOo6CQSSPfI8G8BiTjkNoIuTme+9WeG1P4U1MhNZas
LAWkBgayELW/mKzg0at1WKkQSmk0IZuprfHll/19tmvQaoYAGUCt1b7d9UzJJyMG
3SpfkyvWa8Z7JWcXshQvTu5zqZd88lpxrcCe6B6EyzFzTJcIX0KxLT72DEtjlaW9
1LyIsDuMdV42L1xWpEQ5bced/uchOcUSOp3TzBh9aO3yD7lWpmBlfd+Kku/ne8Ii
U5Fj142mUaleUOvzMWNhx0caeesSvBVMn5I8rxEJGSiQthz0mjcTEnfVSRKun5Q7
STBK8gDbRwUXTSN2U2Rv19wVodn80oeHs3ZFCqPp3jh/4MzHuCW7wHgLyHrbEp0v
i8lffXPEvBHa/CIGSxX2/D8GgIfUnnzJT3cWzmVGvfRcV0bruhcRAglve8SUseQR
9UR4ZE14VM2Xs+vZVyQ1IEXOS6uKpUH6PbQNK0vusRSE9U+5nSyKkXZsGGrB6U+F
liyE9Ue8eAQQDj9AGQKugF2P9vsqhBKqRN/DlL2zYwJNsfWAt+fTQM9TzR4zSSRv
1uk8Va8I6W08cMmQBSAWna/nptiVhcUFVcMINyXfEVyZOK9EKhc3hbz6ZnkFWtZz
LIa2GAoypIQ/hu7gOuwhV8R0Zm5p5by2BtC5/BzdPrByXmYKUoJrsc5mKlH0HYq7
XKY6mvQrF+bExSwouE0DLM968r4R4z2iP8aX2KZydCf1FkSNc7LFzerF3uq0tbeT
WrpfUlpUYSNGJJwIzpSU53HFJu/+525LhOc/v4gOTTd2H8lqA6BJCXkwnn1ZdZYw
Vl7Q2Aqz3CMNrz+LfiditKEaprgrob2O0x6Nz9Q/p9VknKbFCtn4jsNMgomt0EGs
axplwuocfJoqZhJfSQD91DMrps6H9jxUNpxb5OxrIy+qGcLHvGa2JBBhbNtcSAZm
KXv3yD59mHt3ujTndJr0lpF7Cq3/pIHwgJmwgYtO2K/Q4xPmBRpXKrZolajcknZl
QBTTZgyhYyfp5x7iDxnXmsGJyKXxPk+GwtB18pfFQYEYjIzUCMVebDeggtZZOKh3
wC3DlFKHrSRCbaQXkTPfc6FeNoz2k6c9SdQZIqK5QmHdlTLh1eTC3SleLRtMluF0
nOQO09gP9waDwXozhPzAAV/S5ThV30FhJZZSloIof5m38czTWrvWGUJBIxjGRnWj
6CBo/3O3x8x1bSsEwC/fCNEV19iu4ypxdMhP2kSoteh9+US47qobbDpxm98kD3S8
lhEeGQl3WvW8JsHcnFIIHzi2vjo5X98lsBw9oPEW6rSvDzgSsMF2A7Cxtu2N0VCT
xC6edlJfmc14f2lFXNGLSPdfd+aL83eR72ThCa0KqdLAUG3F8bCqDi/VroilKQGJ
F9WQPliBjPW8pIr2al4Ss8BkQDIs6CrvRxbdoVGyrhe/MYXM3+IOkQLIvODGOkeI
5JeZyR9stwQAV8O9XzGNb+KiJCmvKYN/zZOf9vylM2TSLmIiAQacXmHZJ9v5wR8N
HJpje8iGk+iX/qEelSrsuiRmmPbFcRf14fDP3v6a8J9mPsIuPxAIY4M38HzmbaNh
ARsbHozWxH3i4m+8xqaYi5WqFAMSHDZ388HiO3n6AF9RV66edijDlqA9xT7oasip
XEdU6j2Q5ha0tH2PdDUccU0HwHbXvPY3Kj11Dh+PTgm6R6acoE3S7/3vVP5PCG8N
YtwcGd+sLmzSoKMclbMIjAuj6pfpJNotkA/0DHtfa1OLliKTzG55IKFFCPOkgjME
AgYPtPLW5XVDDB0ZcJprTvwaWuyzCzToWfXtWhJpnzjvhlLFmh5OK1FNfpO2Yws3
bqhsqdt1P8tp/XpKADM0NgAyJWYmfmbDrQbpNi7a8ySV/RiOB4teTAIpL/WNtKXF
e7X4R4LaekASu+hHKz9kyewAXiwlwVuxuJFvu+VQwNtZY605L7NmKka+81+jwMyW
7d8zPp3u+rrV/wFT5hdjiiEdlkr33ed3wcHesGst43wnJuZ9XuKKKSz36UD58Ykl
GxVsoLCLVvtBweQKbEIYe77vGTuv6Wbf1YHZtH56/0jaxVafGL3RyjzufXS3Xjw0
h2mk+Ggz5n/ECmYtTmBG9gyHz/wzSqOsZYU1f+T+U8oTYP3X7UgsUg+MbZNeaYlz
klbmO99+Xt3Y1mPsfwSbw4n9Xx8mwiAkfSgkOi4xGdfjPqhsELEsadPbUoHVPH+7
SItyObKB6DG6YSWPX8XSwH1y/Udo+GiDm3i1zrv8djCdYJtXjo+LKYqxSLFU1EC4
8LVIA9aMiwGa5F/azhOOyeMdg3wyxt/in0HvRlLeVWai9bbaJbQNs+j7t2CDqoH4
XpGXyDw1MS0BC2kpgtapAUSqmTgRDWi262B7uxwHCdy5KwdN3+bYVzct64sgOfW/
ilR3+RK1zVL2Rz2L2Hlu4fWSPEWKs5NUD/1s7/ZTJCG5SHHxsuCJrj7VF6YIna/2
F0ej9ycOZXqVK+mfnJxLQ8VWV5gr729VsQGabz43WGEHGV/mHS0QP6G1+hz1QX5p
pQmFz57iU7UKqzsjj1HpqOBhGyjFZCBV255OuXV3kzcvKBBWskcZB1TS2HDUoTJJ
Ar0D2fybzIjwyei1jFZ+8vLvV/majuP7wCqPVFjoKkBxNgpNRBN+BrCGld77eWlc
sxmd+Z1J4OD7u0CZA8ff68C6+6GmdE7e430NoA8E43qk2ED/hJuQ0cAbYfEOym9e
UAl7V3BbX7nAw/13dPE90+ifWk94UFx+N6l6PAA/wvXNlv6xhUJlxPFoSXPte4wC
7R7eYIKJeL0/retUABLtICaI6/VzjvxzEmS8CRLS7nJliajtxbitOLNm21itAR5E
T2/NnW197vTsZMzl+06df262QFHB6C+VjyyF1xFsWzano/karSSbmcLtW1Ftg9+y
GV+5zoIBYLsUjcx6zHgTGjQf2VuWdNJXamSE3cgM/QFsmxr6oQ556dOen/+m6ar7
nnf5MD/aktw9no3RVRU0QkFtxal7RVM0oWJ5gEWBvPTBy6hgnHzgtF9p9fkp8Rll
XGIbUFt2CzFllIvyvHdSFCuCiAkS4sT8+eX+POYcd+lI+dHSwnDzxnACQ8R1ZbCU
u+aRbzQ1aXNcfJT7irjl9X8IwmQROe5HJdTxywCg133ZBZOyh8ZryfyW++vRT2a8
onv8/gPjtL9PW9r/JQ1v4AbXEy3/14NZC70lIkRkny47ncydzIwc13jkjLNesxjj
DrlL6jO0Ub0AoBpadM8ibEzi7OpcMSIM3zs7r4B4XzPWVrE05zF+IHwzXf6Z8P+W
9upxWgRhIxG3TPwuqVssBEyitPBoLvxlZtWnQqt2bzyoRry1lcEM16DFXTle/5hn
Bf34qMz+YnMJOool2dw6DU2OossCM5+0WLs4aItCVgFIFdadK0Iq8acQl536wGPK
87oy9g0PS4Ni7hZJahSWIngh6w8zjVovvZLuwOPhSNakjgtPMLWx12bAgbHEmrko
bjtF2IaCS5N4m+uC1FIsga1r164CreJNEq+tv7hnST1HwAbEqRJaTw9uthmaYJbG
8d/SdNP7Fjgkm0QPr9UngiupKbH8rnm76i3JhbXts35yNUfK4lTQ9x7hOi7ho/aw
EWCkWC8JZrKR8rMwhpXhsFMSp8bNuntc3XVsEAvtqLQ4zZMO84H8LlP8XRvLH3m6
Pw8afL5IduZeefBrCOgm8HUAno7HkXoQCxOYuU58Yd+QcYBNkI20lyHgeztEGgNA
g/7NY+7oIDspwaOAsMV1Pwz9gaJQHceV+wx0kKy5GR+N/6hT6CYLRlwQ0sZi56dk
o84VBvfrTsPpFQMnkFJVq5lChIz7AOA+VJyS5G3ain+th9RZtouIi3Hz0E0GCqR6
BkhwLfjeul8iPrx7YyGUvGvwi9sg79/7+IREW3qzJ4MuRLVPoxyTz1PxJGxXSAlW
K3YpWzxCq//L3CeYbE38EJ/5JYatc+rBWjNPmxofvSAv23s6BxKkzQ4lKS/i/5rx
EjPzwKASoAGdFwkaaqd8eic4jQ1wdIPK/WSBGUQrZepYJBSHQPSxErtQeE4co1LL
g6F9Xq4vEOapJ1stDG006TMebGx1boue+6ACS6i5+pkv4K2pL2VyBXIDRzwwBA2z
LGmRzRgUIuTLwB49xfdud3VCzaY2PyTxnnlNvoK5V+1FyZrzB43eWiPooriLX5av
fU45AVna2oqOcXtim4B0UVkTF34RRxcGd8ZW/e728M/gaMutLQmXWb1qlEeEwZfD
lH4l6rl1dB8VsMAFYBaobFR44HsfvXme1GdQO6PstHVQhNXdZ2grHalukCL3GnuE
Ca7te9TXmM2fxe0Ydryfk82+MwplEYVVwiWfos21sZ24GoWgKMq2CJoq3v4pbUzT
4TtvV5ZMzRwxYgChOHLaQ3RT2HH1FlSJsPG14qWuMQufKgQvZA5VBuKQCcWqIk5z
lx4ZBoffe3Xfrn/XzO+NbIU5xNMjxAqmoNiqh+ZQaugYYk2rTT0CcW2qnfqGJMa0
cQSip/DvedH2KdsXU5DWxO6Kx7fRpLQHAB8xUumrQ7pRcFGvOHbVFXu0LrYqFN4p
1S9/3v/XWIDb+EdDKBZwVfa/cTHFr0cjZpWh/gD831kjfSQyxcc5KlcAZ/SZoOM9
hAQXGDq+pgZVFcxjAeGQ+8JY1atBdx+AszEy8s6TUSWCw/aPfo2Em2XvwUc/XVZ+
UJxyb5yoOkbD8Y5sO19KaR84G/t3TGoQqj+J2uOQMbyS6qKZRiV8LS/T9SGOicOm
lC0xl9sRZ+bYA/WXZ+9oRDXQ3rSt+yoRC/yoZe/FnlIhJ41x1h+tlbDiK0vySO9G
iAWHpyJMidtdBVyVDWCEazOzYCpalhy5OldLVbRWwSrUI/lltIDGpg8hvTOULcgX
bb0awDzmNcKKYrO5hqO0HhbHPHbzvylbl23KKFXSFwEDdlknf/tolo4HmDNy8qWO
WeXzzULEc57ScvI/Yg46ynib7NyccD2ZLp7TCbZvOGAZAEOHYtr63AWbEmVlenAL
4HS8EiN3NiAs4B1ylLv63XLw4N+UGjOQN9+8DYDbCqZOJSZENGFmIHGZQY+DI8Hm
8vzYTRacY3wrr+DXlXVrh4cLqk+BxR2iwd3zM6lRwWg6OYDTs4gJgHgEKFdBxzFx
MTczuYvBLZAYG9lmdtqhiQx5GsW1pRNoiJiRE4PrSW9AEPeBfDMowGKlD/ZkXIE+
mhV05kO5HQo5MAXd0pSq7l1+D9Yfpr8j7mCYJ6282XBJwr8XT/E6yDTnXliNJaKw
DBkwN9YT3Oivfc5qG8cqX9MItM4EbyAlPEV1cz5ZuRH1RM2KmFDNN9rdRRBJr7FI
A1RH+/l0d2CxFgAOF+vyjDxVrP4CheH/ac3si5WU2TvUizoBZTQGTUiDn2baaHcZ
skNyJN5D6FLG7p6Q6aPzZvhg1aWTpJgBwNhzgaXmoZTXicKfStRydREogFSH3KMm
5SLwU0ib3IE+ZLU++5Ge7NkGw5LZYOWkdTxeSQSPMyR3filNQOiJnYp3/jctzLxH
XIWxNuTnviR+91m3LUYXkEwnsA1jzzeqk4j2lxiHL8gP06Lj+M3+dhj3vwakvjV2
6aTe+i34m6oozlb3nQPe+THSeV2jcXAMCSbLCDIDMymUJqvrMI7S2utlCoQn8BAU
P3augHL67lXNRAtTF4Px+euLLJpNOcgDFwqkSsUE8D78ksjl17DPXk31qwKXQGUA
BDCriKMpUFf5k1ueTTHUnnZlf8tKWKG0+WkN1snXcsKUCwoX7nd0I9XeEnObPX9X
8qP7AjZ0kgrVCFKXDytKX8R0R2JcCFyFqLNjG10tNT+hXrQXK7ApS73Y3CT9wMNj
RWJ8Ow4e8MECUDKLhd5NkGUVGN2xC8yUV0kHpAke5mOMpFA9bEWMC4wD4coVBDXJ
L7JsC+3jXV8nk0KeRqVOHUBk4jsokjVkGcVJbGefEKWvFh0uiB0dqVVszkVbQ0DO
N44/I67WsCTh+vklDJ0/R+IlSNA6xOD5p2QGfLWpiainaSdOOQaUp7MVarEL0VPP
Ukj8jJahuwsGjJMmxfirop7D12Z5ahzwPkUxvG5/62Fe19auHgbwaFYO41xda502
+s0zQP4ldXwKvF4s9yC/OoiS8vue04Cpfp/86IdaI70/LEWuTtRr/DaeeaDYL0pL
5jd5V39kQwZ8GfGuU+2EfMg7cZJ8auszg6bszkPDVnpeYAfWxg3ea51tpZuPJ8k+
wsq8458+CYeCpS7B23AXWB+JsPNp5f9OF68YyB9USHdw0aDRU7+j6S6InA8dXg33
BIP+S8tNlPeZGg0hJ1C4Y36efueBb16sJ0hwawqTIcAvX5baahDs0KsqOiCIX+KG
BXYYW+M2G+dKoubMapXalS/oSJRVR69BIkn0p7Qp25ov4lUnFsMbQgjh/siKcPzA
7CqhiC6jggKAM/y5aYggoZ7a12YcE3hDIX7aVXA314gfBpFbRn0UaUDK4JrJ9KKB
4MOMaILBtBFkT2z5hjQXZM6H/QkOAio8UHefipTQjFbxrWeLPPb71cYHFHC1Po2J
l154vOa0hJgnjMaa1AdYKlGejriNT6mpXoS1k7508zWuGqDXURMDA8JBOxosAsI5
UrQ5VcoZMDNgbYEzzSGxfp4rTFDQh05a+X+BX3NGQyirafIUui56YLbk7GdY8yho
02V5QjQN01yxzcoJ2Msxsz3RuKtLRU9UZ2qw4MTavUxaQeH7xjxh6bMONc1dnBHh
JOily67osmAmUKKlmYNfd3qpEAJLAktfuc9LDe+fgYhb45GkGktBiyfhK27aNVrB
K8eU67FufelyCLL9evhpdaAVAsSPOyn5vGaTaleQ+C4xO7bNpwzumisP2tJI8iIY
bKKABcJr+kWazZwblQoH+4tKhZTmmxjmPtMjg1Hx0vnbV3QKXEqt55ZZK8gadqlB
GljpLAWY/5L3qAswe9PPvQqYrX/+tivRypWWapN24RcESqDe/7Bmnz1geTCthHJk
4pyRFDrK6NFRaR4j72+4zhYM8llULl5lAwhybLRL8n/dBRsHQqTND49Rkl5mpTxK
bIKvmmgRRMR/qgs3pm7oshabinkax9MuKsFRARdzFJx50R4zH42hfsuGeRQcHUUx
Ihyugnraj7m2gzhXEfqQ6juYwANNBHo7rhVR+3QQLuRoY3lVW0Scrt8pIdoMNrRB
HNqr9K6Vx3yDj3cuzpYrj70m1whVmQm2ljzv+v+G7dCa0rrS+AfH0PIR/f4g73GW
FhZ+S/gkf0wNCE6OondY8uchqKZSWnuK7wnYgBvFP53ZFV59tvOuXKMxO57nNk1M
JK7CruTXCsHdmnMZkDBWE/VGMkgVOYI6t8jkHNVVPtzIrQUQeR0y5aTfknYOZfwi
bG5QvGTTIRr6xQwLKOvo6/An11Zg0uFvQu4PRYNs+JM0qWBZswzZNW/CvgSVN8Nn
+AhpOON/6nBGiMPEjWFDtJTFBMaeS311r9TxbdAykyZsO1daANcGuyAB8IpL+nPi
s0fZUFqYk3NaNXeDOwo3GK4gyXSfiRwwqPJfZ35luf2aqA9IfyVgo5a59JE6iR+K
k2MYXNfTKn3cTySg2zOnpNeSyfWV9P3tG0g+o4vfpe9Vuo0yzMv4WgdtmYLYULzk
IY5YlDhs8aDdKI2v/b3JYptQ4mlafItZpDUIHn5B92/a4FDu7WlmKXvRqyxPYyhP
Or2Mg1pISoICA5w0YrnMTL+bXmznZ431vApf6Rs+EVIEPw++m6uCEynEBfl2QDD0
8YNzrCRir1BaNX4Sxx7kKxGIpLmwLV/S4qHnuhJ0TTlNE0tSDqqpnxRSOawG3zY+
+InB9XTFRviCukrerlo3SsGCTzmFv/SjTWZYkfwa0rdY1152PupSjOJppUrfF8NY
+9F0O7w4tuDQpQRAFcIOENR48jVualWGnYMA/L83FBr44t9B9KckreS1Ilo8TBTB
VEs3X0OvVldg60lOgUIISHz+LPY/TCJ3Br2V11wUbItaZePWxzAgZF1JUQigh4cZ
AZEIdh9yv/dEjMPX5LPaoJR6KRw4gI7LjvmS0JD2CTuUJau+CR5xpPYPG8XrqvCg
LE3Ujsno817J/sGjwI1ueZLCjRA9iYXuKXCbLP1pxyu6iPLEsYMOwxBrXlmlsBC9
SiXbK7w7yW1LsUTuMotATRCrmkrHZHS+LxT6UpMU61HxaQ6DvxFtAElWOGLgm7xc
FAojs7tVH/MWUX3YeKCRKKw1iRu10aD4SDV8yJm15Cjz/iPJe3ndNBwOQzeT9atS
lEDPRGydRgLOa/Tpy52lscrfwVjOF1OC3WR9q+1BPpI+kSkY4kHwR+81RlzypXaU
vPVBcpWURTCU/B4fj+jIJq1IeiJNw1xgXbnzHT9gyEUNbARsNZwm/r5pN6wrbg8K
u4w7RUlbYBnqU6svk0koeEB74BssR7pgQCqAePxOaSgNc11+EvCebmFcKhHykk5O
+DUKKEMLotgyWYDCKzj9Ci+9xxssDe54EJ0JsRaboWO0VtF1J+ty0SZDWnNJ5OHT
pXOC5WX4cg4LJi6SD7/BfvieDgWZxS0LVI2EHXvDtY+G6RfXk98cca/qAr+SVFcB
PFH6jpYEkZAtcfDCWqJEI0LyvsbL5vJxZ4zUa54mn7wNZtBKyt0KDlHHHvng5Xau
FzaDa9Ygg+x8MTB1FsSyT10OhptF1Bu6LV+C4b0juDSCaDrpBVvSQ84P+OUUT25b
rVBG6QLCsbzlFPE/p18dIlHEj9qSeCChUWwgkvFZ99MQQ2B4wOUzXNUf1kpwWmoR
Y1dp3DynQAg93vjV5onOgBSPwby+o/N4whvIKlRHcKemvDNWrYOGJs45aqSNi8S+
YzsggxdqHuEov4JZHIb9Wf/o9LNGGTCAqRoIsfLHSXrdV/d3fBKEX5blga0bA1/3
kZ45Bxyk4vMIe5u69WZOJntCgbuau2QXSML6+YADb2J7z6Pp9v7rxZb4llRS+/jd
IrLq3Gxr7xmebXakyRb9LnqI1PAQpXXxllqQrZvFRE3ogkY7j15GpucxiHx2n0pa
bBBboPsWL0YayFHjf6O7hvwT6+DzlRaFvZ+qRzZxWBJhZFej1+9iE3eCiUdCHXsh
3BK+6hqWUJQSERTslouDKuOEKu1SK80EQPLTJCYUcktQVyFXb0OEUURabU/MaZ24
j0MqpN0bjp3ZB2BtqDvjhtXBDhLAlgKkKCcK9JrSiHS1kyHKw3bSxy2z8aF6ghke
c/vK5wyFE9Qiuas4wcArEMHTsvILsS+L3k+8ejLrvVyFylsSs6tyRZBAx1di+hmz
Ia6Ic2O7v2NM76NwhmbeQ/s875EMCwyx8Q3ilhqqlGDWOGWIVedQNTfG9w4sdOP0
LMM60SEDrO+m+wHGJjm019UXAXly7cv0GYJVBx0ZIzR1IkH37vcBbQI8GPxaKN/C
jNqkC0Qo/k0fsv2OGpp10FmkClbGUdD0Gb+2Cye2DBNOxFJ7cQjVpZyk/qCIiVDZ
1Ry5uqJIboTka/Gvk1YruZrknGrd0Z9XTsHthFPykKiUw/BsnqmVoMZr05NLfg74
//NASaKXskQAcYfUiVJbfJ+lZoEGbqYWrsZPwrbsxuuAtdH4LmFYJu5W0NWgqEV/
DQuEVC7HGXtSO+bKKO9jpXd5suuwyUe7aVzmmyGy761qWkPxigcLVrKttsnG8tjB
obJEms+uWM8X+fCz33XBLvAPUaKk1UP540EXT7z4+Am9xdzL0PlgfzzNMzvzaodI
CrSpf4VyobVvvzI22tftjr1UM2ylbxrPfAlHoVnwQ9ZHbMjLfPOM6rNEzIyPS4lW
cdi4uJUUmtnDw8umb+f0ihUPzsK7FZ7fuTiVQzjiI85MbEp0BGKIY7y7m7XPmA/Z
di8+ZY3gFadZEeeJ5aOiOT9WfjSzMR6L0i3n6HhNFzshbuJQFiu8mcXm6V9/oJEM
Pifob5i+1jszBsLU4D40a1/+n9K+wFfh0sMW3fzLvrsqbelRbeFzkMbVTAGcadCJ
tZFqJpOfXJAeIlYXqKUDhokk6iJA/mZswCQAglx6Zd9c82C6eqzqzN7z9qQEqTNT
dmw7PrTEuL2vpqkTHHvmeQUt4viF3idse4OSK4xw6RCc/kf+FpaaP/fvhbfUbYzu
2A736RSQntmFcoDrpL7hSQ4LtxlQjPnsN8q2quUjZJ4S57+y/4HUsCXRf+hmOZG6
mjaxPK+fqHwc/wnA8+gY/5bCy52Nq7uEn6jQWimeWi6f4bcaPTLtBRMUV6WeMMjE
A+bE4n8iMtPoVDl3b8p0wZfUND2JYzGeJGggOPCMIL6ptO1g1v6TBOddJLrXnZPe
TMBVMrmvM4UVISrQLnqnUxTUMCTua9k5kPxTaq0tZhKj0Hdtn4maNfKW3Xx39vMy
uQkOQUu567GLqo0EFswdsL4aPTl+zaEiQodHyxzAs2OYAn5dezIIrgsmbH3TMxxg
Y22EU/8tuCWJOqHEKoD1nqCQosjEYhRkUYgSvFVrnUh71UdBflTldMNLm7VqT+Uq
k1BCOZokn9PMwRp7X+YB70hkZKR/mqsX2LhlaFX2Oxh7AbiMLWwrKTTMxQZqHjCD
Dq2qmL2cipEL6/CsF0HgqIVwOsUM8KzbG0Q1gHMGyVnydP75y8o95d1CRO1elu9G
TVEsJOgPYb4OnTfmwG6GERs8aLVApd/UM0YzD0jVCjGuSCmtQVNPSv1x+VDEeEwf
qTM7GQZOlQGCB9xoEup/ywoqo6T4DC6dg6tC6Pzo7lC+5dAh5a5yPVWlD0ysuuMA
DiAlSHJhBLpIgrYD7GTfB0zCKTIAsHA0DXmwL3BPSB9yArT2lMxMV/hY10hfxB3y
m1J464Vr7LrjHyHefyInb2aftlG+bPGmBGLLY0FWGk0As7I+tZ2umfserpjNMrAl
Ni2dYrfF3KY5uYql5wFFBkTyU8YNgf8IjSrLrbhkEVLux6OhZVjeNAre2TdCtZYH
Y3v8M8aVwRxRkiL4FXu7AFpolgOLZTveZANwszyZlCBdW1FcrFjEzLdgB6h47y1+
MfTP514eHR3uOLaLCj4OmU6nOXJwxnaIojsDQmbHgI2GtS6PIxN6cO/E3j5yV9j7
IMLU6qnDHOD2GMjX7/hRhWPGrp0h5G0/elWyEnzPth+9c1WtoBwp0N7viHpA1ycr
mpiCEuI7lUOAZqsKgmP3maC9v3ax/4Y5aNRiGMqVGNLbYn9NJArC0bDmkzqVyR+v
vc7wV09AEw2nEZFzd/PDACAt480e4HOtKA7BCx6zyXPpBWAHXiDG2v7HDoAyB7Hj
TvH0C+wtK0zX90n0zQvV1GtEWXXitULxOsUBzSB2QAU0B56A4oA7OKMGFN5Abn4L
nSUjIQ7iLGZVd2sHazD8xH8fzRX9C7Tqy/LXO5InmBGSGSXTQ3V7inosOP3naubI
S7Ygdp/o18IZcjXT4srGQ3BdSZxiLixltXrC3x3iYX8SWHVnPev9nGa9dKqvA32d
js1Kj5S6hrpBlH0lXVazi1h3/sCqVjP6AyojMgmvIcHRfSYwcXv8nYpXEVwTmwm/
Xvt/o2z/bJboRXTVgdoU+sdKt6x1UnWurOSANAPhpDHTTDWgmlHiFWpTTVibJkA4
XlXQpGxVjQ8tbdg9YtYhPEdOhb1G9QXIwwt+U/qgWBK56+YWog3MS+vqRE9wsN3C
BGe2dVvG5xAZ54Vh1ciwvHnunn4hho/TKFim0hm35OeGfZTsoFHR2TUzZ53ujbeA
WPhoao+1PwauT5olxsf9DUwO5cQhxZJs5gh01p6dyFtqyXtSfkqM0RkkiqMhxLMT
fRJCpC/cpKu+QZUoFo0omrRtciu8p4lGT0XkOduW/P0EZ4jbdLYfcasdFmXwnkf7
qjz4UOqj5b3EgRvTIcDrSYCvspJ1WpyIz5bBmZedmR3QNLSDbV3PaeRib17uy6B9
0s77isHS2tVG51rohVkiMfLPqnL5mzIGMjnUPidXjfr7G++8X+eIMcU4vNGmfaNw
hdk4zyX2xiaKt48TPP9cl3R1IzGAa60+sOatfiTHGBNSVnQwFofhwA5GMOGOZMDV
weUT2Kw35zrdporDSWo+FqUenSUK0uXFYmj5vKENZ82FQMePLuEcHYJy9LYYz4Dr
34Q6t6LwWWBFm6p06mzzEULL20H38VPrYx7kLRNoIhoHS/rRPiPAkrQ+oe674fib
LZquc0feG0LC9oWd6Xw7Z8K3oky7EJrp66YDSg9+URuabbaRVWWRpfMrqMA/xwV8
ILQBgWuHzXJNylqUEqifSx3OcrsIy/gpO7U8RIZFSyMVEDwJBGVlsxrykweIdX/p
v4WvfSmF2ZUMax0H2FGyl0w2MLkFvjzQCEukbEsJYii678i4bFWDHkImfKo5Q9QW
WcTz6MaDm9MhWZ1E/ZDCm13elr+BCaEXppmAeXXqeS1bqaRgF9e1yCa+TyaBFDvK
X+4kFtqGDFCg4BK7MxT1N0NAEwh4Etj5wt3oz6J3oSRL1puowW2AmaKzZWNC6HQu
/7vmHZH3kl5Rjrc1OuQAWV0KdFQ5GuxkzCQkTa34AaPWlUqFKVok/dka+c8cGoPD
qdnOORJ+EdQK2gbz0BwcYnUgyX/Iy+GecopRX6aWQIet2d0bSWiqV+UpPYLxaHSi
AvgGxnjHfTh3pKKYTgV2OGSzIqW3d1RtVRmUoo/1ABBd34vOHfVkPOercTXwAskk
SvmkJK9tfcWxayKlj4SuqTuF4fLxkIPzQTHSkkgIStnE8XAL78CSx+SbWoKDV4BK
oaQCicfj+8D9E01Ns9FpDdqZmQ/FYCApXjSDxK6GvHp+I5lMHFYezuVX5pstfGlY
Z52m/1lX+VVcTKsX1J6WaGWhlkQZeOkYka8otFsFTM4lj4oi8aoF94DkkgCJPW02
kIPh6nJFwxASG3biJMJ534c1Fd4/WA66RdHP3es5HeI4WBikgPMeiFlHRAPESzr3
CgZGfaL5/16LDsDNsK+L/+ecC2MLz2unYjLnDhytUTN7oDe5vBUwvWPR3exNAtgf
0+f166Ebnyhtfq77SkLj4Lh57fTOzosdVoxmXtgfLSWvNjDKlV/sxRut2i1nfg+E
on8nsZ817ceqVI9ictLF3MXv0SrKMLBkQLGp286G/f+SFlrqIbOht613jIW8uYcr
vAhyDu4DFeOgyR2sPRp9Y7rZJ/mnVVx5bjgTflAbjF/W1KLTSl/9MTHe/Rwcz3QU
wz6GonhmAnVzquF0Gvn/zSvSmjW0Gz7BlV5pLrM18Ha9sIxKbeynZi314RWHsnQW
2VQmANc3E8SgXnUqiBdTGRNp5hrgg93FGsqGNODiNCS9kVeom+RcZDFpJA9mgj0n
XlXPjy3m+H7GFJO1dG5SDEAdbOJ+CAuozsiwTaqGjbPXX5S2aXN++4ty+cEMqRWA
h12jzvtpA+AjSH1aVFPLdISym6hpA/mMbUQtTmq45sVmVMgsdcgSNgANnL9tGPa1
wH2D2A/Ic7y4gBtMJ01K0wXfie+HGjqTV4i6jZcXqF9gcrjAqriF9BHu1hDMjtUN
MZfhDCHRDAClNuyeyBN21WKh6Gj/qDpIwKV+nsxmj4kfCB1048zdpR6KneJYVe8p
kYAmYTg4ty+fajyrze+f/Cl0CcBImK2EsfntiZ7oeoPGtrEUkRvT7TPp+VpiIFgD
lawtND/xCBkugeJoOKyUzlB+RMo2CbhvYOlhf4N215cG1JpiGSWpyxa4vuy1hCHY
rz1/de4YAiVEgAI17grfjt7ZnCqLeSlSfGfblbaMtYG8tgPIUdvyhfE5kQM/YO1B
/f+bTci6f+mISerMMNfGmX9oa7vjVNmqAbk4tjaCQAM8DrX3iQ5HGHnDQQ4PiZO8
17jRgEkRWBcq1nuR8qAMpxKIU9iSuxlLHtc7+sXPXxpOjOhRGOWl6E7mu1YaSB+v
QBTfVCMiDG8xJc/9zTZ3FNE9wSAWLMhqBghBG2dny/mCEoGHkjQFt2yuHgZleqWe
VOHOz3RgP7cniuDS5CzFNOe7w6YAZ7V2usBcL6jIq15cfDIgXie4gjXQz9Y3Z4Ur
WxMfA6oS+dytJJzA1KaLhU2+mlRehLvjLOPctJfCPJwnM5r1eJcdARBvqXP+VNhJ
LP/MGL56l8ch8ZcG7Y64Zb4aFjG6u+TrWti7IKARH+NbOyRku3uPdb0R5kZhRuH5
OuV9ALoHRxSrM9829mjRWTeU3wbNR9qfSWaIi5qRXSeeH1mpyezLC9w3Bk03zBTW
86SUmR3RfxmZTRVXrhc9oaNUh9s/MZ/YtENay3Jwqyjel7YkWJSQXTy0eFsHzgi9
esjfBp3wM35+fIMTWJdWViWdg/V4L5i8q0eK4ajI7h5hZzSE3HBx819vFs3ZZzww
v58rUMisJn2G9HnfBn7PToUWXcjZ900h05JLZcIouFgF0a2YPta6JvsYXUJ0lNjb
wNnMQ+Wn3NsegWt8YotpLZSXfFi4zmLcw4WPxW9K4dmu7m+5zUaSYIhUH3/vT/mJ
8f2Lw5Lnjj6W4rcsB3ozHjZ9pwmw/Ki7sAITONp/SzTtg9XZltFv/KnO21g/HSo8
uvY8IN8QT86RgcNmeEBYDfZh8MOpQPj6ZHDwzYBf5ZopSpeynonronFHQA+EK+6S
TEkIw4QLpHjFHMUvwpP7xWuCVQ6h4S4oFPfY5QcrQOQylObRBDsDmqNOnnS9b/6J
PUYdit4PZn/7iwJ5muEHobIO0JU6PeCLC3a0iviDQUJgxNYkMEuZiNBB85fEsInw
eyHhmftdfD+keNe8o5vRjHKo7VcOwtvhhP41GHKF3AFpraU165MFzhRY6fDkDBtz
heuKEV3tI5xQA/vbaKgwqBAuBvztMfWuGyQycgpZkkpTeSuXNueJ9ICtjONezons
CVbKxMKQhVjedzDxX8iOsjxrNYHi3b0Nu8HFuEqhJYkMeDKKUkoVDaI+ZaHlwPsI
AOAA1gH6iqLFvGgVHKl5VwsVz/nPJTHfvhIv4gwACXDN2djOdBT+DS5epP/OyHeF
dDtVprbBvFcwik3E+tJv+Y71TBzI1nQJPj89TWFiHgoedBJeaXW5yVtU9evNwcWk
NzxDkHSIbQ7aWQGbEzJHLrScr12dsY/GCZLWwGDEgyswH6hxJL9L/muaVFJfS66G
Lj1JGkPKpg7nskZf92p0C/NHzwsY+i+vqqArmemilunKEW1gmns8Evxc+SeHYwk4
sSxRCaJYySaE2zKZtndGRDKArpmu+gmzTVHbohfSI+FDBoGFo/UOM65MHM5DiwSN
jfwkgBlFxpf4x4g1gxxEFVaUD5+6tnEonbd6YqW8EXfOhu51tDpNvOoohb2fei5q
b+72/fUXcLCEI4K2pqHlKTSWVlG/k3231PTspYavMRy/jex3htFSM1ia5WvoyXM9
3VRhrKuBN5CoswXV9ppo4kmPGYY+CKowpbOc3Vi3AcIWh9jpI+2VkKWHJahlTACh
Tjhz4SULTHd1nZkM0cUl7yTgykfe3G9fLJayIdnLASZfrWpYe6gTzfzQGUMs1M6f
/N7AaBIO9SwldPq0+xDDosyhZ1sn3Fq/rBdNGDKEQ19hctrfcSR+WoBGOhCBwhdQ
sJ3iEhIkfxWaCsMPcrzsS2DWs6AXTOF9JmmaKnmWzhSe/Q4ZejD067d3J61rQzX6
wy22nTtB0TJxibIZDcZtZAFsC6Ow3u/+yKTY099KGHOsmDPWVabuocJvPi3UCUtK
mmzg3WeW+ee/E76zl6ej6TmYwTG7pBnX9wvRV+MB9GYLjwArBlx0yRtxB+KUOhPB
Shd9sxDDRk8nOeJODRGKpaPNYCEizLKC2W9bhG4+xIvOsmfP6hrB/ujBBAGEKV1K
53nrZjdVt8SKjBHu4DoqyIzFVrhUBgyxXg88ftOLymDVdF/XVGEAFqLnqod16O4z
P84Pzx4sOWrgm9pl/Oankf++j120eSZJvTYDbXmw3zPlDDSQJxmkdqlezIwYJHor
qxsKon0TtOi7pv/YsHiNlFPU5bnZNYFExQlhiGhwGNT55DRbg6HPBB68v8I6NQI1
XGF5rtJzghKoBhQhQQSHwtC9LQjegIUBPBKdZUKeGCvQihmEVe4XGYcTNYO0Z2+Z
1UBc7YwiWNYyYSaNPPwJnb4GSUjBm33tKMFPMJ7WDm8JMxdJJwjwJ69qpTHmjxqq
go2AOr1PRI40Epl9onOdeDcnmrQ7Yhq1o2hb/fSockPePlMInckK6wb0WDjH2ZvX
fT9D1M/rOPeeyFAP/c4hCOB54JVj8T9ymqxd2XegkjD5EXPgGDcZ7DDgoErkuGOL
AvBVUsO+wnsutPGjoYR+YOn7m1zUPl7PvEhHCMKAPCusasXQhgQGgMtQCbcmj/Gx
b9m12qdpbMZFPU0nIsyxiJERG2TICLCpycrhjDKuAmVfujQq3UC0Zq+94v3HB2oe
aZlswXHw+omyieM05/qeE6kji0VbtZdzz7KWZY6FE/wT/LUuzgSu6qVJitYFbaD8
BY6iHOajKB2Z0FQfoJsbY58mxgctuORqdX5yoJ9oBL2HIRUZwjGpyqXMLSx4cTtH
TanC+SwUK4VbFiI1U8q+iJpYBr7z9/NOu1Ms5batJGExOatSGFz/EtE0USiTnsrY
2Oc3T6NsDGgPQhS38ua0L0HicleWJarMgnln/Lri+vulPR1UsrUrrniXW5GfjeDz
WzfG9RvuN2yD/RsU3EKYzKqhAcdSgwUaJ3S1wXlgy3CSWO2ajhAWq4Y4PFOu9wRy
2f2WRYUHFTJDWQqd+HJ8k664nqidLl+mpI2fk8NpwMxKooq4D00i31PLF+fffCn0
UJt6k9FpkZXVXg3kZ36/IKbGt8TOEr4ZcnEv6HfCRueR+JgEivrCPa1uR6ClCYai
vbYzLGH04dfMSOgTnUwYOWknYPbLFEm1ZmLCYUgLli3rGL20q071He4FKC/i8yIw
tdRfkCUlPgRuk/uDFed7EMlCWQOu3GIROlUqBG4hF5VJD49ZXJaz6PXec+2z96KY
NRqR7o++tWftsANsHNzEK2DpVSfMU92uu1ruRY8eDH+Chm8Gcagqjazoo+QrIPSq
mBYPj09AJ47q1PgQnKP6KDsHlcSRtq7Kv/Wu6U2/o/Q9ex0131P7gzE6XX1v7SuW
kRgwK7OXEjo2advMtNt6udVorW2ZdkYhld+eUtWxsAQNx+kyyYj86YRYcBbx3ohW
fioV3Qi/yIIYH8wkBFt1i64vnT111IgOaVuxY+TaLXppr0ZnQBHOiPXVKgivfJWV
zRyMSLl5Z0QWZ34h71Lf7VwHwVhOR461/mftWBU9gOy7b6IM8xxJbkwuzKeev7Dt
Z9VQrj642klYopXK/N85VBWT2L488BFtO4j6sEeDk9DC52evB6O/in/qiPowdKXG
tM6E5UByARfTxAeOkMj6xG2JTXvqUM+2GPpdjymVgaaQYtpYvlBDJxbhUsFgLPxU
iYP0PtFOHelx1hqyU1XwRWefL4ZE7IDhgyvPUoiLLiNDtw9Dy1kk0Kz7sU+nmD/S
+JznVO69wTwx04VbNJUtejIatmQzRDXlmPvPIVhm/4vVJTz6JB/HMAc0xxoUMUhC
sq0JRVLlhomRM2GTTu7elIUujWFb1tr+mqMCXOdaXnXSHRTo48Aha0gCoS7LQFLk
AIgYgbtskGm+OqaVfvKB++FUWmQ/dchN2aoWhaEW2NntLbTguWYhyI17HdffjNNN
x0gMuX//1IoHb95oppQDG/SN03AHDAelmmopBkc9mOoM+awX7DQQQIIYvku0zJO6
bPdxp2SQAEf213pNuUluuEhdB7Y+Ix67q9ePnRNRzp0nRLmOJ8FtXHAcbgBbn5QU
NWOPXDOm9u8nhIjRs0+6NUZyAurZgvwx5fUDva9RKFDqfy2IV/eDZWs9ISVNg3Wi
Sf172FkvMKaX/AnIKgPR2yVcKEqB+poLICohDQA3DdLRaVoB6pM9nnSwsnucnnLD
eIGv5EEMUHN1+FKosMOuC5hfe0oX59FbO/l0XmEJxaCqo3Yl9H+XyzLuNK6A2xul
himGl1BeRcc6zIlbvIYZrO1unfBIWzjCMwviCykn/ohXACo0O24vZiRIhQ58r6tT
KYGQQxbyxN9zTxrXbL5Yzz6ohNoT6w2rYD3E720Dl9rb/8pujN7bmQRpqoknoEoi
SINNxsKO45IMp8t783CbKlD0+uFtUhCqz8ZGf1Z8bx0RzHLvoTYJXkTXu6HXao1L
GzyImOi05Tf8chGneM+B+sdCOFCFce0qX/UX0nCbSYUJa+ohaNm78t4AJ3SAWh1n
iiVdOSA7h3Zk/V8r/1BYBTlH8AbuFrgxz9mvBeYxACAdIPHNV4myovsIB/iSc6Ps
ThGSjg99Tz07a1EWm6ZdoFw88GRYspApYTfVdObCOZdXR0Vd5OJjYw5xgJZzjy7D
D9R0N5ZRk80O5m60adjR3WEi78Bv8UWC/cUBG6ov+KGiFGsFr0wcIBuqPhb9HWyr
G2ucPthPZzk63c8OAGgSyn09lYBrjRnScoGwqhMjKMIEKVUugLUzSPy9UCS0qeIs
m/sFHL2H3uExc1iMUzux0XklukvrP2fFKE0UWsH7UW7hyFAm1nz0W/8hWFV9rLY5
ObkwEW9nczzPf2Lg4oF/mE9hAA2nN6okxhFIRHxfH4BGgozap6fUosAV68m/3hp7
RtXuKMOjKx+lCO5I39AW4fCxYEyR9w/6771uoMje0/azZhxnotkvGYQzKDuXU+Qh
qtzj7B/NFwc3kHwoWzYYVC73T+4RxQS6+3io73nZNX6QXzbJHubUpvGuArDDaRDb
Stu4ISHil7tXmzidW8BUhMDeSN0FgMaKzu1uXD94Pm2S4Ps/V3CQTN3whfrNRlZm
/lryRH/zTGUFp1u8pQKI+dzzsMfG9tdm7qZcNlK/M3dFhqeTclZ3U/0tbSijG5fb
EiVxRmmFGKvNdTeKhwOpx46HXOwG3eqNwSNYbxlaqT6huyDcwaNjEIO56hX2Cbi2
cOEOeOhbRQfsiXYc7sgufcS3w67uMBi1W/MynLUg/YSTeMMnu075jdBswrdI1wwl
eAnN5Tul7RViVEDvfPd4ugNHdLgQd88cokAB4eGib63JvUtc/XZKcWlD4ESNe1ZS
uK94rTCTSNxZIgYEJPsVdQtJR3/+0Kn9mEiDR08bkck5uksP7wBh4yJeLKLssEWs
C9Tui2DmcT2LFc08FirIhvo87MeoLH+/b6v8ZaiLsHSSpBOnuvGGe/m029hgJVw3
hswNhukkAfU3NkwrUdxjmiG70O1xayCVKs2/pC3sUIuVeOfqtLevb9te6Ksw/3ix
I8K1ANxIpgwofabN9P/OB6uLzA9bZ7g2rd34yO9S1aNItyRdFoH8yG/SoxWVl32J
6f8tru+qmXDvmslSmnmg5mxUt7Dwv/vW/jwuc31pXm3IMEfLLXgg0D7HFYEVCPfL
wGheIc91XKzcm3xtFtsPTbgMPl/crv8x9ZwDWDq36b4caWZAdEeWHw6MBfHPFqka
ZWUE0FTwUxwahgVEknFOSiXwf9r/HASnXimKvSlvnVf/u7kafy0zsf4wmG4zQkKA
RY8etLKhrt37z6tkqguoc+tgVQrX1sH0jxD4r/bzdZ/FHzqEeieA714n6OAklZyZ
NwGSWKmyNCA/q9m0AEovcqwRamgj+vTdfkzJ9qQtMS+qCXWq3Gisf6EaxrKN0nyc
7jfHFDGX99/9VCgpG+ZX73F6LQjso3lTiFFGYg/rilvvvOFbHEQzgZaY7kw9kEV9
72m/dQdMS+7tzzQf/zPID6uZqCX0isy0z+8eKSBE8kieOyjqN73ZtVL6/AFto87J
IwQDtxSQ/YoHrQHFXaqfuHhtYDh4qmaXW554InszRD0NkFANXYabznyF/ZIXqiZf
cIQcJopMkycDRwbwCna5tcbbczQBPxhhFh6qt1YSCklBhOlMcb537nCd6UPiQ7fn
4tQee/TLbvMEefLPv4Ne/uwViWlLKu2nZPLPAkei73y4HY6iJLIVFETwcr5CKhPa
rveN4FZ+keIWPkh3ws+Kat6hfpZfqFoxTBQ18BbSN5xbHsp4A/LfT/pz+srKXpqd
7wAmw5LLaCduIo3nxbThyIXfyJ7aCMJaG7adJDUR6Cw/wGVKQ/T4YzTtHwm9MkZp
5MxDUlG1EQbFl39hETANVPYjUlc174dBgagcLbwBJoXdg6fhK5BOPovcFV7yqWv4
WEndoBbqEbwzQ3kuhhtLhnbFxkI7jIDpdAYxk1FTWxoruccO4HKGMDq2Rbr24Kuz
b40Ibf4LSOl/DoOc0U7adUGQda7JWYdNRXzhW4WQWnDk7rGzLtJAy/Y0XBhjSRgP
gWiNfO1ZfkBYYjudb80YK5vb+KIwEdJN4lotfBBuPV01V3vS35sqXLZbV1+cDDRR
u53jQ5yN/B7wANI4ORDiyvYOb+/UcemlRe1YDkJve2T8VFY5CbdjkQL9gjcAGsXl
AD86TGJhdW3PK7HvTdY++UViWIwzs6R1NnWb3Sy0O1Y43osiupHOelBa3C/lfPgB
DXakTYCk53W7uHRQ8q6VT/rluUJ51d3vY1y1C801RYoQSDdp5KlxxriG1Y0Kj3XY
kcOLq1Z4i482EZVCPJji6KXgpBIQqhIHNH8rhXUCIbMFeMXH2KQjIv2/v/4qHVJS
7pwWg5kdiMFHEEoaQIBXHRvSMpnlMms30Ucg8oJGJXMQw99rM9cSBtiG+b5iZprK
ycPAye4qPelryg0yrCR3Hmzaig3BTtd+xe2g+OtgDlGDJgWZWaEanstRvxeD3gRL
0ncIQE6ucDnDHhK8TE554RotgSLhaa49Kgfryvu/wMikEjcCGeL4s/H0kjf/+P8v
7hFBpyj2WCu9kHSUYBxqVjLxh/pXHf96FNwjy0W54Oi5sRvwrHb1HPXVolJIYBu+
y1MPnMezWGue/04NEX+fPOo6QYHCsw+TIcBobE+6PsZ03DVBi+1VkbzA+781jYF3
CYbPquNfRHgp/B5BJz5Gn340ef5LOALKWlZPW8z8xevmhx1qKx17fAB6lmQR1G2T
naDEeXQYWfbSeRMigH7FayXC49OvUW6mO8GTmmgEXyijtdbqFX/Jz4oggQPtSFTZ
V2EjCkJ9k0d3xR1iGeByuNuIfsaHOSeQjS3k71fAowYxCzDot9ci7PxtkkD9rQBW
Cuo72IooChi0sYnISVBFQ6lHJAgiNcQ156iAgCNk4RL4wOs6WSmeeEKsRGGfxbRg
k7ZtsGDKTY19+SLEoyWeIPChkoEn2dGlAW0ofF2JM+k0IMrxWOBbtBsiwo9L9svD
v3wTNj0Ha/lQ4+g0l8QEksjYUssYwUytFK3PwVflOsyhuzhygb6JQXSMZFS4af1e
+UWddhxzFgsbM6uSxIF5f5+9WyTcNwFdObPr/4zm/MvG2XCU5Nq+a99perl/WbJY
c5qC94FKkU7NQoghf+BRkK2s18esVIrhMiBw6oAlkg7D5d1uXC6Kev+c4w7w3hs/
a4wX5a4LQzzpI2rNfLzewGlHAMYYVEdo72UhsMiwTqPDx0sF6CqsMOd/2I0MVXp4
eUQA297MjKU1NK0IfKbkhLcsodrrgvmEzT5L3mJZDzZb6OqEIHFIxGFZoOl/+9+U
CIL8aW9/cM1Nb85Q70M2R8v8XM4E7A4LkskjqzjhDxJPkjSoGzJt8E1i4Eh2SrNT
4Wysgk6RxlWARgLqwT4sTP2UlcnKF7CgBJxwCiL2gytNu4y2IA6+fYmIQfLooxLH
sjmLYaqzW0wnb+1dWwwwfP4dkUKegPuGj+4kRmnJW8dXbeJzjKqr5pUE90+q4rxs
bWjLE2XXZy+0/+eR+jvOoIM6PEkI9cPRwQOIrgAJpXSTOPT8TayuxUayvbARFfhZ
96krGJ+p6sOJkVzwIyitudsMDeL384FJkVUXqpQgj3oghz7nuz+Z9i8gYqMhJNCN
27fHEsB4VLLPTicgTlWfUPzcARbuInYutIMNugOxTdZVrkGJPpTCrq/gM6xvNcLP
M0Bg+x0DrG7tq7Xdf3VU8xUdp7ScJEt+PlwU3ldD3TQZpXawUtehV5h0QvNrYS7w
QgO4N3R0mX2XSRU1Nuaz2vvN5/LkjB7kpNBlR7Mq4cR9kFzhmAnQZ5yNGY3uie+O
y7F3FeO5T2z0fbiLKF9h8yLnu5y2fpps30I8Jik8/Xq/UN7LHOK570olT6NWHnj5
vl6UdnwATrGUHV7E6wAdTDEYGfRPnt52EQnqvjDKZHJWeaa+QTFYHj1NG9nRtH8K
P6Gxu9JbCiljxL82c+vNY1hMv6vARAtSXy+GRda8eAIQMP7GkGxfxtLl+A9r3dgi
yFgmwpLOGFzsNqY8l8mgsUdqM50j3PAosf3sMknFALLJURndXZyJ70glBM4i+KE2
JYLEMr3S0tCNshfA1nSvsdky6OLbzUPLQIiJkfjTxFQSUkTDTPep1NL6TN8W1PuO
YHTKII0QZJDLcuWvSeQwuq0lSQ2G2O800MC9ZCIRN0N+HA11L2C4f95f73lLnBFf
ABz/4p5PoE+pawgTbqOwPI5oaLTtjdSMSmLhTJETPCqJyaR3C1BTakYiOkorWT4B
fVEhjcm+/EdBR/9GBy4UXr06hV4M2bsLRDVLTdUG4E0WLD8k1nA3JNThDuQVYjVO
yUZwNL7OS7RIjXTODAk1Bpg4h3uD8z6zgYojpaoYoCAmvxDZ8ElStMKh2Ps7t+sQ
A6bncxhvLSjOy6H8+8DAxAzL54e4f1lOhT00nZPTQXvaH5/kVjcFM4I3RQnOTAkG
u718vU4GyvNLuc4uIMsL/CwLRnkbuBZfh9V+5gRFIQnO7LSAzBLibfGwVOJdAGF1
ycpEvUzb3SC0qu+Rx6IS8DK1SDT2uz7i73hWgvi9jY9J2uoDOQs27Myy8gLCkEfh
wtBE5YLCLpbJki1HRoWTGirlOB/sOIJ++KxXvsX0OYP+5wOaKcN2PW/1E63gI6dA
b6Lr8ZvRbj31D9C+o538BOueYXSfLJJh9T9o8wL05EU9/qgaHEqjDhLRcWQ6TYTw
XAQRTdKzcJi8zIiuKHSWbSDfNM5F15ej+OI3Y2JwiuXzef5UqMbjUBNj8CUrBmE9
dpJn8wSi9X5F8oeYeXzIQ/+oJOOZaEyXIoFeArMO7l7JpQV5Y6c9+rtVsydUyFLH
EG8FZIlq1ziIS0p33z02HEWNdT7QYmdALfB4vLXfPlNz8cf0C/vBqJd83kXkRQq5
qyOo+QnGwfXZu+89M3HAQ1h/qfYFYuTivjayUjVftjY3ZZd0VAfOOZ1X4xRK72qh
zcpAiyi9Td5iLDETEcZtFeXv038QTVCs+YJD1zo/440vr/RDrVe+xP0uhZufnHf5
O73Kc3EVo0oyYwp10gzvR7yjVtjnUAs6Soa6Z/cB3vwZE8baJ8sJ1C9sJwYJobcD
0Fmc9pp3itggNrK3UHr7gHqR5DGy8r3qxqRJ9Cu8KtiSFIXZLR0Kc3lc8QEBsx2y
cuYjS1mTrcqrY4UKHNAKYjY843NCXY6gpEUlKf5P81SsPOKySuzRF7zmKxoZ/PBj
q4Txt9xcX4jm17oZ4LBtuugwOEoTRk8wjIQvp4s26kavdXnQMShA/jGap7bRSwTX
FyGpz7qqR0xmcL7QYiVnJ/4HGkeFvBw/curX1UCSMAsrRFa6JyoY6PGB0HPy1OfK
VSl5LJmurzUbHdpxzryO9TeluPN+i8W/HhuJqk0Ck6aVACDzSlvegFYHf04Bdn/B
HoGqFmoKnkFx02cobilI6tq4WYHnWisFn2tCqEf6BF2bbkVhKqMaKyEFF2bI/qF+
MqRNu729xnFQnGbldEeiC8SmBio6vYP6u1Qo3fKWIxgqjELS3tkYXF9cmr18WsgI
dgQTjrQO8OmxAaXCD/FB5QAK++/8t2BBd5cyQ9+QYoP+YtvG5tJ5unOq4fNGvFj+
ElFMAcEpz17EWR/ptuN7v/d+vFXzgEA2ua+R+XReKChLeKYKQvNO4GG7fEANkukE
VixPl24YNJDS2/Ukse+6Fy3sbhc0CZuI9O5Mu+GgNnFSs4eSoRo9akGUPhjoWm8r
QHJEp1MLqA1br+7epSE4uy8fLTr4iNFZnThycogv+j5O6RmS0wjTB/wnB4sdRwib
pPtyGaCiI7n9kUfCfyqFoed0JVjrsQpSK99OlvlIutoxyDTraCtMQUCx7teNOUzj
EZxEv1d+E/KIZA974bYaO2uTs+lZ1GCZCZCNjnruPh3KjDPpDwZar/UIeeYSdLBN
T37c71cNAGt9mNeYZseJijorFeCNfdiEG34cncy38klQMQCyOwGvG62TL+tQ/w/+
3AjB5+9cYds9AVP9uFh8qFBjrM95s/s12bfx6dV5oScjSM2on3UHK0avSVd967So
nBRE3qh5kWlBY3R+VgfrF28qjmDkwYtLVX93VyINpRAARyXEewOZVs+VS0scA+fH
uMrF0a401stFiTleqbwaKqFG8bJ8+qy1kwU8G0bGnPRetNYEj3mGSCZnQ6spkDW1
X3Fz3IS4snajXE5K/x+VDoQPFCoXQTRT08Pat6d+0rTWp63NtSji8I+AqJQfqPqv
MHaE+pMrXOBBwU3CiNYq0ZqGjtMaSkc6Mf9ocGrSHt9QuW8ldAlLb25G3EKO3adt
xZvbeFhLKqUsTrysdOt2pkw9KrEzmWx7mDiDpBviJRtph1DEESGiM56OwVid0PvI
OwV+rtWHIkKVdhcY4ewIy2oknmA6UCNBg8tNUh3Yx0cpKt1GKXZWn8Z36FVX/AJT
B59TV3SBWSvw+PMmKoJwooKMijV3RtdOqIA8i2pjga3tya+JNsEwyVI+LCE9mptd
cHjJT2agDXcUcDmsamJeZ8qN+p+rnRNBqkz33OOxI9GpuQMmYDNHGFvXhUne58r/
/fNNobzd6sNbKIS++qMIwLlyRO2AIDwuonqOkYxF60YQyL3weHZf++39MhTSekJI
jn5w6MquwuS9YGYSr/PPdUsonQvovpKzGN5ApM70COiSbyqskLY2jj906Xbdcuos
dcJ73IIdHifc11mhOWt3/diVnK4rSQIU+YGZ5vnNVFCUZf4/66X5MJFOxnYc1m4T
ZvcbCAYd7hUFc4SYj+F2goHStMh6dsRrrxDwcZJt9NZWO2HIN9tPnsxzmboFAWgN
Oi40MqcWrl97lwRWJ/YenLXw7A0SJlwc1cTY+4aN7Sd8Ln0JCgr51p04yYMhAKer
pCRtpZ7Qa64UVWnpsSWrnQYOadxhfiqx8uiHeYTFVp4XDymXRRGa5T2/Zc21yysG
2Y1Z/l4+AXxgZKVprCMx0Q5+yFgzSc0SOZpFigkwKSd6abSUw/zS44/f9fkMVc0m
cU2tKJRPLCqSjV0Lton1q15LzjC22HKCgO6Z1HzC/sKcNSuAxLp9QimRNLQ3DNzt
1Gthm0RuKSVrNejqvlcq+z6MswwPvfZ+OqGijo+99gyF7+hXcamYjO4Xso07ThSP
G1PiTLcvo73Z3/FDlxJrmYkgk52HkNFJtNbtCyP0VZRBcOppTAwUBHXxEruqtLC4
PnqpqkKIr7bk+iA77a+MxAcMtMsaoRdfSJpx8AtSYTzRckat9ckoYccU4i+JPmSG
06CtHdY+vgH6CcjcU8MVz8R8J2qE1PvrpBiF5SIAl8s6fmv15+J9ZTgTf2sl9Xv5
c4IT7cGiPMUD8THBUM6VTfdO4re4EpTSfs63ZtZNRz3D+l9Je1KpjFXq0wdFWpff
rfwJecfrrwsRtcXsGcCuBxyriF8l6oGQsTIAXIeOfSn/E+McrYvS1yUMSu8+6inB
LUIm+PJWDdLPFACC1uyulTclspOMgB+u0h30sGcSOVbZAaBRIDURJWW/TIlIlfKJ
4NW30Vs2ztjYnergv3ZxxOJFNHPjEraDIMjg3YuFaQ/pMsLwGy1hCPibaAY3sN0p
eDHgj6eDfhLG8YXVr8B08VpapotW+ORp3lDZ7Bn25IlgJwO+sfgK9O64SaLHrm4F
2WeRVrYzMQ61P0/4y74qWromXVCEd4aLo6kHEqtidREMKhATLH9nsR1000qpFjDP
RtvVJUuke91/GSKZwdhDcIjYt6bXiz5AbXWxJQ3RkJe9ztMFBtf/gGRzSsEr3azy
wnygMsvKxvXwaG9O5d8TUv2F75E9NVHRLpacntWLsJzciUY6JK+/LImH32th+gFw
iDZj4LAWiK1CSE7lBM5M/v6ctPdKsHYt7T91frj1InzncOaLEVAdeTz2ZTDv8+lK
VGBKBpKYlvKqgLcfkhBfIed9knEtHNOB4N3QoAafsL7MiK7Hg90PCfN+I31pAAs9
WjgFgWH6Ios/SzBtbyuYBfeATVk5fTcqi3Iqr146nBACeIEqZY0S2CEQY60Yk/tJ
tiYFV9/Cy06NQuVRq5+uoEVf1RwJKDpaNGgcQMKH2qI/JL7uczc3lgMpjYh7OLu4
5g6wkp6xHUmK69xcLF61KY7qx0vnqWg++Ih+0P5Nbc7chYzyb3ao2t5L4rWFG5LX
rqr9pdiA1DhFW31JUNJFRDSbckzCWji3CqogGjnGTV2CyrRdGlxLgMprPsKyCRjd
Oke1v2oyQKx48rC5cDMLECjRRVjon03RUb1Rej6Po7ZZHIpJpR6gen45dSe7/A9x
ml9QPnSX8WZNRc2CuSEn4KTVidOYcwuIoSodUYksNV6e1lyoq2p3PIcZ0N3o0Nh6
PVdAXwgnR5LB5+mFM33qJm1sEFq7IjHVPVeUS7KGipq5BM5xTWvrixpEtUzXBFfW
XMGAaWoP/NH7wVEJZYPZ++JysuSVJK/KS64uAYDcH0v76NPeYvzHos90K+f1kRj+
DnvMXQrOVRLQ2XJOcbhDWzBJsIowCagc7csij36VrSCUimUkP1KiRd1pAmPuWuZk
pgarlBrDVucTxVwjLvJJ3JJyz6LE+g2D7EdT+28CqiM02WVQkSQlSan/yiHYnsaD
t6XOYAT5XidvRf/Dgy4hi+39z2jYmBWwSL10x97UPOAqDExK/ACLvWAxvhKlgT/R
Us+3TRwqZpSm5fkGgpARWVKwD2sgn9Sx7NfyYnNIYzjifsLnV8Szsj+p76Wv0TFM
AkVA302J4BYpk+Vla6m+d9O3unPvtH+m6dODhD5N6GI/fwXdrpjcaCDUwaNKadMh
AgtTWBa/30cLmRMkTwlDDF5PVKIL0QbXm3yrWG+XS8KDYdNN8awirYga0CY93M8+
BMFTyqQgGDk/u8vXpaqpv0ZjTUfoNva/YJYh0FEybpyfjJR4dyJFHMG6i3egbRV/
7D0brV7XOnJbvFJyazKkXiZWKx0C0hv1B1HIZBC28y06QtoZD+9tJXOG//n/d/Nj
y8+CRZinDc75nX2R5Ce6sHm+AKckvDg3dHqFHDZh9t4qaYN8f17l3c98pZWwiqtK
ut2f407FAEwih1sdn/knvm1yP41sLDINc8hEu8f9qZo8lhh2Ra0yTl5YlY2OtfRK
E0PKD7mwwMnlGlhUQL1tiiTuKW5nH1vorIODZySPVSxZWkR8z4e29odQsSxqZ4pr
HRR/614mRPPPBGNuMq3PlsrfBhJatxrGEG/4yW2Wue3bEg/uRUClLTYyTGw86JL6
XeGkXsAUYPtAXEswkUO/ekW0dCF6eHX13pOkXLep3Cd4SsKzYP+/+Iz8VfhEpsiY
g/JzDAvPdWF6MtZqaKKzjBH5OOht/m3K9QrnTdtCNznxPNFccMGdqNEpoUOsorvV
AJWgmIZNBnDT5RQ4h+SdZnH+Zwh42f1/ybkGLSb63WyD/zlRmYvHHeH0R9JRoDjb
9Y0G7mX/KFkkQUU4NFf4nmCMkqlymqsVlOAsgwH+Kr80BWcZrrXquJQB0m804laV
Rgr+qRppQSaBLZ0yK6CLkBUSMEEbf7qRHgKZ87YuOWaElBDfHqAuq5mczuH+KRtL
/o3qOzJjlmqBo1a/M9KA5t8gREXml7QmAtKmrKsnBUShQcmW183hKBZxEa1ft4lq
AMfsBE70bU6pOLFG5ZDwtUfPt4zVJA+kt+mt286sdpOh5G50U8leLdFGYpwTX6Ky
VSzEHNUeHjS0EaCqHNzjlMXzx/jdljZMwokBJcQxOVZ4uMqLn/fBYTSheVDSczNj
wgf1llvvYsZuxAHSKXc8vN/H1aasg+EBiWDcDjL5XBn2Dmnlb6uxsCyZfiM+OFVJ
44DO0DbyeiSoZeQBbgYKJnc1+EYMva0OEB9joYrTGEysQS5JOM+e18KA8z0UCbPk
28OhHTtO+iaEq10AZTNjV4YucYLAADvm/CQAjOmk2hRJ2BAFr4GnU42KIW1Z1fwJ
O3HT4NgvJi4EWO5jxMsemO5mPK3jZZHQ5STQp4Ly1T/k6A94RNFQq5tzfC9vi6yN
ob3IAZlojn+iVQJckqSFhv4+hLWP+etsAWbR+F6/Egw6rNdan2piwXdauXpmDp1T
blmr44C1kYDmvsr6uW7qpx59kS+7QdqPN5JxPljLe+senh66E+gUE6iTBX6963u4
Pv2MhFwPyOofHazZ5Qv0tyb/ioGPnl4nIiRbcdNOz4XR1sZYTkp4FoKC95ARqlk0
1UuxOC7peBXIzbaFKNH6AIs/w9oPjULJwWRG+vqAoRJle0b5ZrdZ26w1FdMjjTb9
62VVR3qp5oUjZ71jRehYC+szU9ACDjTiJjhINwgfes7WG7V3R9Yg4We5Z8VYic5X
jf9WNITGUFDOpMo1uquh5IMYa3r30op3GrUzyaZvlCSmjTgirK3WStePtr1x3jC1
oKExbLhuZcZna4trdc1XqyClkYKy08tMdCNShEj3Wjf83Nko/N7v61XbLJ++kzlc
nCt8W9ODhyksq7F61OAbR00zsrGYIKtudW+11fZ74C1CwXZsjl2jhS/1UM0pr7e9
GyIagKMQcVSPDtD60SeNNSmRRweX/5MDXI5NIYLBtGUNyzqPg9MWVZ6uE7uHYwME
jgXAAxrinjMZNaEP16irBxaZExa+u0DvUmKz0djo8HuH4lOp01PwTLyYf13qeBsV
HpmDmlOrdcX8CxD4snpORizgfJPdlD/DqbjtskPl+zZQJ5lxjXmAJtRnffaDysK7
URNTfwdjLFe5PCxK9eqDhe+IKdRwH552Ie+4rKWoZ1EoctniVYM3L/TMfzXyQo+k
wHR8tZ4nsxj9asZgseA5gQKJjvkvPRGJsuy1HhVJn+FKJDtkxCsrX+iVdgs2BueG
ruDyAyYBGhslx2zeh4BM1KKmR2UHLhT4UlOUXjjDMm7CuoFe2n+2fr/guDoYpD/K
9h8HKZGQm6v4q4E0G17Y8pY6dagr5y9LwGWaXrIMtuE0pwFTqQnss850LuTIAFAP
3ZC9VI6DJMLUje3GiWS28dXBMldZYk8t6HhR1rFAcMcQd6yeutIRI8BZAgKasxiD
xUxx6/N7S5FRrurrjWoTQNuYNq+eqi9lf7RSW7uN0rSK6gpyAwYCclYu04z353Hj
9Hkax2hdLLVH7KTse0CPxWNQWCGKg5QSiSin78y+jXUK9G26Guf16npa88aRpr73
k9erUeLTm8elDS4Xi9gPYDHHN5feF7SgDyxiE3S3ctzMk9tWbk7IbSzG5tKHnV8A
ofsHp7dLAToT59pIx5rEnRvm6xCg6/Ji+XG6ihD5v62rpxS7pJIrOWHfcrJSyJm+
C3aw7YYNS3OFMwwlVwQka8W/+GWxt7FxaqOUFHcD2T+NB4zKy7HDbc341Z+Cgbh8
Ph2CecL+SzzzO0mJjOO7vGB4JdPO/hqZ/QasShJhgp3+Fr3rz8nWzEuukxR7nz7w
g3YS2GMIWrrViaQ/7qIEDHtuA0hc30OsNjTUTfBY7fDUtQvW1E5mZnyVrWjPaKuP
5IPhMFy6hGrsan80WHmV1AbgKaM8BqpiuHacUGzmPaBgzSbu9HQxxbTEfPgCeqLq
xDytXWfUXAuVp9Kmzc/myWIj+S4Gs8Xe6gQSGp3KxWVBnXQw35irYs8r8qxNli0I
y96UV0GTmmFOB0Y3BwTJ5iZBkczGY8AihC1g+n1QZAK9847BnxEQoMvBIPNcgPf0
fMDhyeVEPMAbC5D2Bm7NiJcCwrbOR5h5vpI4//XsN4RK8osm5cbbRceX2ZEkCF4G
tSsrsNR2H0cTFHrImmiw3MGeD6TFPcDZMhI8O090z516NR7ydL+XykM2SS5585jE
+l7YRuCtbMOz3ZuD6bstHvdRafhHPoQp/94wDeb2RE3HEEe+ADUOjzM3K1Z2mFaV
iMTjdq3REfufgzLAIjSaLPjHVPW5sXiPTwQ2u+uj0gouMjmXcRlXDD6AIc1Pr14b
onGNwLIieDUt4yY0wPg+uB+a92tz9b9qOVfVzRtXCTGcKUpfcAwFEaD2WNV07+OE
5PQE84a4vUPwQxLaq0KhTIZj3Qm/GS5tmOzY/5KpVEGqSsvAqDXxIdw227lX/tk8
JolAwkmIlUG6rcEAmyn8q9nBrs/b9MyZTgjmG23PXM2Emac6ZILMeiJ8pz8vMdzJ
+UvWoEw9lXLWzUfaq8JmqzXR2p4w+PbIbspFUPF8XCTkSIxCuAszwBnjosUpL9fN
6AcPWOw2EQr6mied4uZ+YmI6wKR+MsxHAdRp+kvU5Y5+9KayioDNjKf9AbzKdVIO
uGBV/BOkPmFncVDM79uKECToUN3sJt433IU5BR9+ije4cR9JbUNqMKoGpcxasWc7
deVTyqRFawA+te4syw/e24s3uuehMEVy2w05Do5wghHcQ7dDFoKYOz8LXLzI786o
JN0Y2NcHakzvibhEAD5CuY/Laz3jWRoGcbU+1J0qXwK3RhyFaIwyz5zIq2QZkvT1
r1jPjoIbJr9Y8I2Ns4c2xvUJXF3qd4r6xIyf2p+u9L7CzlKHemelKIqu/6HCz7W+
KZaSL09t4yRJzYxxbcJTahZoUSgxgkebeTJsfQ6X0dSjSRT4dHuXbfaeIVX1rh60
6yVa+H8GQFEEbJpmOYB+Si7F9X4oPUEYngGYzGZKXlHVpaRyCmVVA5HeBTczMA4o
h0jRCHpkj365+PHprR6nqHLY5jcXsYrdcjDCBFTM2zNzyu2yPRZ0fOHHuX14+WQJ
fuSIN5n9iMU32Zb6SHkexJhO0TZiwxLPmfYbrxvlosgXKd+hCJJ4KeKvY33AXtiU
HPIAfRjaHTfpKVBQouZ2UsQGLcKzMk2GJzJmOcsBXnztNq/tVayVHbisWF9WNrWT
r5BLJBC0AuOnYEm4oCvqKyv1jaN2PAIWXPUGKjPtMMhuj3xTcFmHXb9MDD7uPVA2
o04BHrDAriPp1GB1bQTSNsw40xDMi9hO9feasogCDFNA2F2Yv8hYz4PORDHe3xWi
/1i5mQVT/cyVX7LEBfeAyGzQWBgw1y39IuhXWUg1RgXCdkQldDaMU6wO/5YixkYB
8fnVGz8vfp95uoBxsKv051PbeJT8z+Qc9voSuFKWAPpMFSCnqw/MkTv/hDFu3Nte
l3GQIUIkLMk5T/PI52KFIQ3Rtgb/WJCFlSEYWTnX8VsBYrN5Ru+U8HDHN4wdylmY
iseSXV9ajssNxfl4tQTIxKZ6orIdtN6RJXT/VTiZ0J5F7UWjclA6TdhaaMb5MQ/2
VZ1+GjKNu24cL9jgBGagsFtRjXtFzoeF96Uxm3RnsPGFWcM0tQoj8dYbkk6dDN/D
dCkLU3xEHmVAs2PFSfdIC9MMDWtSsJdX46lQjdvIqnal17q3JyWwUFYIr2dwg303
Jf9NF7f5+wUs7sTNgr2aWv0BFAhBOnCu4L1Ex3JU5wMAJEn14sdvycdUwbw7Ygvb
4ghMsRWd2h5nf2RQz7lU2wGkD0CKmoN+RiycfmuZhoypaiOWaNBslAnz+DpYoMdh
myfZF3JPC2vBcx62lX+WRSRqSsx1pXhwadTVuBsPGw1NpBL+cUs56SFCChH199og
ZSL/RN5ADqLyYVTBFU7qjvRZbeax1Nq0/dg/7qZgbA+D8DZ5vYsJIf5hcNG2KiTo
WTXpBSXipI5OtarWtI4E9dcICxh1je8UmRL9TtJ37RGMgqI6bgjkPaw2ULwQtnG6
rWA0H0cwImIP2zkRzvi4VNB6vPrMpnRh9Cpn4GiNmXorEn5J88F2DC7LNiIydi1u
T2dW2aOokotMdE2Yq0S7u59IfkQN1K38Oe1otE/04oarRuPcBl+8Wwvknyvjuere
Y68P0G3hxsfZ4kkM9uGSgwW37tWfhDOi8ZQGLoY1OAM0zw5P56ud8SCHtsFdpPPF
YMjj3u4s0AOLvLImOl9LNgibOdsY7dg3Rzag2kNooT/OIBfhqCJz7dnYH7NCEgrA
4Fm9QYnGEijwKN71QbtbRU2XEZ8gDwaXcQEBjGVvDUFVihvAEhybexBgKP/XA0cz
dTLKSJToEfT5KRRXD2omdgXkRlcjT0Xud4QAu4V0qZXO9MUvo1xj+07Ae9b6NQAK
B2+ukh+TI/OX6DZ5gV9hRRH8QM9vHyybAUNsYsPqHJGShpJZkdqPKNfEL0IOOwX3
DOy7Qm5oOr/6JYpeP7Kl9Nc40viih/NhxNGYpwD/YbXAHzC5XNSW/Kbf9f07GTL5
rwCdFfxiLbwtyNzNrnoAAJ/moSwbY0Neevhbi0I+KkZbiC3PrSw3qbyFYxUnb9IS
9X/wPjw0xJ9To0YVKt+P1SAU98jRyy04Jdzh/58lHjfQckEJOzSPTXh53fqw+2QE
2tDyAz21F+98xLzeApgy0Pm8unJvOBn8v1+Nb3VGmb9zY2sl+cPnoTmJUPIYVLNH
8Kkg2hsIPJ1PeQkAnABwcgeSLdH+JxVMH1TDHJb8ynKUxMjy3psuPjgiCuedGPM3
JEoW40d+eLIeU0HVN0P4Io1TQt5eUro+ueaHrxk+CKJeAGszJxXRqpCKF9sp4i1C
0VdwcCvE01mPY/FCqRLDF9Y4XO2XxmL4Xb16VzWKXY3oogt5b4n3MZ/8qdPB2kY9
nKKrL0d9iRMwBc32Nbae77LJ69Px54DtAQIb2Bxt/rSnSRYoVsr2O0t55O5wO1cm
gpZrVrdrfGIX5zXKwzmJShdrrdvoVf9hqLCLl/5H7kegHTvAeg7c4CFiUyz09BMH
/2Ja4R8vF9HxXrdMYSWTcI64o6xCH5sP9BvoLfP83c1rRUO5sfaAj6GBckIPf91A
h8LB3ZoAxkcRsZHqbNGmCuS0AqZMNjzv/qESL3NuA/XAaXe90sZT4AU67N3oFH6Q
zVa2AZ3wcRKnhQW04EQxYX29gEiEFJz8aWhQS0RlVxZxZoIgc0d0quTkyf1h9ru9
y3tpmcCOoak1aAykjTB2ERphUfkFzqx0i26W42VKjK7OxoUOJkMllI3/xfLsDODn
m0ogDL/AFeQNxcYIsKipOXn+9I0dFehLq6te79SNOM6401I1l4U61u9LpzLDO4Dp
WdjSYwqmShrxOmAjlY5YeB+QxuKhKpwCcYO+Ic7kzA80sUfAjUkPvl91YMVk91DR
erOF/a/Ws+lhkstTLDEJESGkvtXVFrXJmFrpsp/HLCjfIWJNw5n1Lh/y1Hto50yh
ybgpad7r1FOhPd1H5ow3cM7rhTY9QAO1aEuhvNswma+VHActgPoWK+38VdsODA17
Rf1yRwn33GXJvARrrzcBAdE6sHfzln/8cSQ8+LJnFDVjLQneLic+SaROhWm4iF3k
jRjQHcC0DJ1mXIcZlUxbLuc568NS4fsD0BBffa1+ygwfX/kfBdmbzMqD8zXcrA7Y
3jui7bs362wiekBP4xNP1zu58gAIJIfSc75E3WAgPdgORK+G2fTacXfAi0qTd/yP
boKTt8yI3iuYjSZ/hsBufqQLqxhCNzf53U99gWWGZ5v2IYXc+azkmkZ0adY1TiUp
pSFaukz23twJG1mwQWCLKdfRYznMf5nmGOJQY3V2tY0MalNCZTyr+8s5YUkeGccY
O86wr5/dWSqfHScDlvUevxg+rsRzV58QizOTCmzEUaOsMMJduKFQzFup60EQj8Zp
SJ8elPNf51L4nBodf+2/RrpNOU7RfEpdftruzR0P1s+8d3+e6m8yHBUgti8XyQRh
T10i400b++u6fH7RClCoMrZwp3UNmhEneyz2ghysZ6/r9WVx2zCbJbU4KJxzUcIr
gXxtVuaygWx+Uu1lAlV0YrFE3+zABWfrlMQaRHBbkO06mN0tje/H1ZKvCfTN+iHB
LfXHyFf9T6t9MfPQw5P4o2fH/OAlma6YrT66uwyWUaOhFCSZUTs8Zgck0azuc2jU
DNCc9PPxYwVzMVjDbJ5/AQHXBa0kf7b4iyR+nsIDq7P7xCtZphD7PZ51l7Xpdgf0
MldRKuOZfkTS/S5nBWiKh7l45bghfswR5+QG/Jg6jep6A7pZaYHNKTE/Ak2mcPG4
+EnfO0TQmZEwFkTlP585AdwpDAWHz0u7Kp0fbZSYXMYBBQF4IBrz9p2WRrM/9oZs
DEqTPDu7TILuanbXId889bj7pKJQLd4WgpdmbY9tRoZb3hwbkgLcDHTnd5Mb3xtz
7+NQtgKHv8hlBUVIE2V/5NyWqZ9t1wtEq6Gnq/UsCJK+5PbB8ZOHeththXafUeWv
q4wgEKTzS4Qv6W5KpE1ntADe10czwYCAOYN32KkIRxgkc1cAvYKH1f+16JebpWkO
0SU/iiZ9fuLpECTzFfVuB7P9ShCuIMRwOKS2aKWR8EspfXZMMdviN76iSOXwhijj
RHVvGi8BTSEtAQXzekAtH6zzdwXUyBf1NN5IKmU2vUNsg7xPloqCrlSJdGe0Q84J
SHRR8uOFuxL+81v5fs0Ziw6qBzjXrQMYTZHj/XfZtdrLTIGVli2vXof7ywT7g5wQ
ewM6U+c4vOFAWAh29pE1LbGHFRiGAiPUo9ilB5ho00MCH8zByRPC/XWWQOifZNcl
BWb9xAeGNP4pd/WdJQroS59yih56wFiHc7v0gj8PMr4zaBFn+ra/t3h9ST3+7AtZ
+RK6zcMFsY29blzbFn0mlbuTX9jc8YMY20FmBTjIVqy2TveJLEBPnm5Qh2MEjLVU
4Rl03xCX432BWO0VZXl2yZq0yFpOysemYuABTv0/y5Tpcrw6kEoVWlsf/SAA/EjZ
xe/58ONu57OeWAKFANdnNYT6sMY/aD6KGAFqnDmODU0YPDyQ1TJcVG92HGgNVjuS
cMpzf8VmR9Zje8/55M06Ry7WofFl1NC3PWgzkL5URe54i7NYImp8OAALoFNbSapr
M7t8F2+7vI/ymiCoKtDNkux+pG/+mb4ibqbxt57fniLFGXkBcmC0PZyjty6E89v9
MilsoDuYq1hUU4asH1n3jPkaasa7XW9BqQClI08JvevthcnATfuMP4BdrwfSQh0y
9o84etRkMyWUUeEjZ2OrJziIpMcTnkat4+nNFgNNkNAon5R39LnTJWtkVLuxzmuU
PNc3TdtWjQxXzM2J+B88vYjRvwUw0H76Kqc3WAbBn7MApFSz0xSBD8p1oyvs8DhD
HnxfyaqpDD+6FViEJpDZCYW75hrYxKu119AHjYUWNfQXcWYkLsoShjbMExcgruFr
MCZFvy7Uan9GXGE0AN0k+tlRhDiGuZLZ1B9YyO+rZEhiKhZa39WeCa95CH/VAPVP
Rvz8rWH2LNXRJ8vixdHjEaUM9CVqCigZvTG6dkegiKDhgofAoJX1Y/HWlp2Ivt0h
0zAqLr2MHwxiqqkEPzfVqcJtfPuhbsMLgN673fHj/GE3+MydrdlAM4OnReALC040
jsN/KiQtojnmfAhNY0JkhyH+hvHLYO/HQAMm6g3UKbSEIJoKLdQJZrf/ITRBfbZg
KPsN/wB6P0kzfID+4a2dyzAZt5sPTWQ9KAFRMvG7weByqZt3lTYxy2iv47DRIQ+y
0fK4x3BYUs1Qozhm7UqU3jee2Ij8rzOMaWeK115QHljKJHh2lTqBjNxVJVdp8rFg
e1LzffZ5G01qqRTNZPjjNCFVeSXFo8ONlHggRowjXExRBDLUK5Wm27NaKhvFfhjc
/qLoWSUIbKfM6K3LTkcnyW02DtvfKpHFJKMyPwd0Vvz8U3/lEdpZr0RVMANSRzla
C2D3AIQ01gH1KK0Xv1hl+j+PyUvB0LnGpzlLc1ZrrwSv1NIS6gaVyaZEUsKtqH2h
AB13AjOFa9IX2cJejZUSH7sc7Gsdw6j1LbUJxNHEWpBsM+4SrLfZXFtmt5ukjdio
GgDhx2XSHGx5wRXXGikhGxYMu0rPey9DnUXAEBubpNHoAKwUxfVNCYEI4AlVEM2O
KwT2ArUVLgh5Mlt9qCDN3shMy+mbpbSiv/jruAsV9OHYT4q25AvC35gLHEl5gugI
u4JIUFBa3xg7VGl7IKVzGd3qhrB0rsJEl20T7dFc115U4pWDt8YYDqzHrGdAopOB
H84rRrB2YpK8zANsd/CIHCqk86+bMkPMN6gXHhL/J9r8qBrqW57n4/b8sUDs+3Y6
hS4Kffw/US250z8q7N0nJ4uZSZesW5JbEXGcYAHOQ5UJ4zsVzYYrsWE0Gvxs8C7x
Gsr4FBjIw/C1eSe2XfGEYekAumq7/SOT+DAN8QGQZRi0kxxOQ7nHYcChsFAAjT3p
7/heir4FN0T/tMCT4a5lCw3KZhpgJVx0IuYUGh1hYf5385nYKKTXTWMPNnhoMhOZ
cZsxz4gqlYX2cr96L5vDJa5c28Jn61hreZEW9dKJSHDtb4OiI1ZAs9pt4PBPY1cN
aPpfNCHujQ3fNVfB7aRS4Rawt5pBbei9C58KjIWa7XuB9pGd9dtUzaHE0wvVAiqp
EEAxYIVFsj/A6pd6qAokDbv1Ab+Jemv13mRPBheaE0YZ8VBvifd00HXihFxY5ujz
UEPZ9JktzWVIii7/tDXE4zs2s2PMLSsE50LBwNeIvHW5cocW9ZruYBf0L5sqSLba
E8lcQm53sLEbnd4gXOzdR23bWFUsqgD1tmuRRnFPrTRbRaiYHNfVyGATYduECWxn
89+cJVAX+0CGmUV7kuJ0oMSplaj+BQEfehtAbH4OobUmDiIAH6bKTut9ILHuZe2J
1GegYhhiG8QIUPOVJSJnYsvwt6Z9DCAQhIRvjycA1sBireP6nanvihqkWsOwBDFa
orqqIgfVt3K6ty+bsfNZgt4fiEFDrshh+huDdDJVptB859ysJyVAlHPlecwo7ucK
vQ4f07hSgDnRkXf4u3CuFqnmJPEtiwDKYEOkOhmIQvB2k5mlzcqRdNRGN7zd5GC2
Xn3qbCw2E1FnXH2qy8aE9+XDJQkr+eYH5dnUBpEYp+fp4bCo7qZlPZaELCSc/wrr
8vGP6b3huOrUnSCMSgFQRdmNOZeKtAmsbmgHbogLrMPFMw73J+EJNjAdPdd+oKtK
l06W2DDV8Sbdmcd4QCexINoy2JUy9g0g8ZjI/OTq5BfhyFNjwInGPneu5Xc285TY
yywnpBG3t3zpGzYQ9UtAcaehNiQxqjSyEbAhafmu/Ej7lqpQ5LngUCFJum7SR5mM
ghnCT0OAF1X4ioZRr+kSqxlFTmtXVDJAt4fJ7Aji0JytewI44nTlZzWgY9Nur6Wc
iDH6xdBv3b2B4xm1dyZVtB2RaIMNpUrhfjZeipDukTDtGBor2L+VoZG9GitmctCi
6UR/pFpS6E/cI6FQJtn+CUB+BsGj9lKWIGk1QgwR4oczo56uIvtgSrzG+4/g1iJ6
QwOCuQ1vfMFbTDEscmzPL+4e6RNroS4nUVR2HP/KXXoSS2bQy5w/JQzBsPZNLuhr
5wwAET17MiAEareK5quPNyc4NXot5tyYf9dpu+JDDMZdD+M1qfcIRqrude1PYNTF
oadMZvb/LLXuG/NQVzeKUBAi4Drp1zEICnoYl9jnhL8Q0Hkg2UiuoyzxLNIn/X+8
CK8N4KmnxF8EnAaUyygXETc2CxD2t5B/UlWC8uGp2g8BG4euhhqtWTZwrOBuHCI7
4jEoc0UoNY9rbbwf61RL0LR66/rmDuqwmtxooYMwc0OfbF1rk3lfu+HOSlaL3oYv
r9mCyWWkoHmml5YxT3FPSxvKQ/BnlTr+wTuUZ4O/A3u2f+QFsU76zXsKsm0G/uz1
WQ11KedWoJ06+T1CS63i6R/2ervIOF85dxNWW/PpsXwF+uEZBIp5rxIl5QvJHVSE
KLvDcLw7YmV9iwbZw9n88UO4QCG5MUJc4ovQzz7lqATMl86wDcOzVbXH6OaXqbD2
Q1k6DvgOjQRnrDT7Lr2ZboCr7ispZaGyIAi75EMNmz1f9OsO60/IgjYjVvdh3YD1
mmMfS2SU7MZa4Tj1SXREIjML4sJy8r6M7SSfiqZBTW1CcmToRJdzl52MXbvMU0AW
jbJhyrPM0e/Qp/U89bpF9sXm/tGWNXwQ8wqAhlxocaF+dC+5DggLZJxNQM4cg8tr
VK9C+1FwwxaOWs4YZ0rAWz5s3M2NtUokrcrW4AdBHx4YQuhbABkQueBBB/7viMWF
qmK2zZpZM4KfT8fFbHCVm43ZVsCIYDS8o1+nwoY6syg929O4nX8z41RJ4aymbob9
6JQ4wUSh+v0X2VOsTuGlvK5+I0HnnblETMSOY5FE5RZwEh8LTpqohuNw3st2dQ4i
EOo+8VWLuxIJ5UxwAepDhXPfCfkK8EuaAojrV9n2FADB8VFG7xcYxiaJL/c0kR9b
RKj5/vGyIhafWPNFuWPDmqEzNgdNPD9aEUYtKP0ATXX2qSwGcTtlzGriPwcTZ7ZN
uh28bGcwtlUA3y7HaHS3t+w2LaQSzYAaJ7io/wGuPEidHxJfkhuXRIpXLqCYse/N
DnEu0l7Prudru1nu9YhRwGK0fGpSYS0j2yBBlnhZqKor3nQeFuahSRoQlFqwa2qT
PYbAsueVSoacHjDXJhR41nKelo3wqtzDq6ajdcsBL4cHWgAQ10zMY84EORe0jSSK
GsN7KQsNf9Iu1Wx4KYg3GwN1hofShnaGg/ULuKvDv8ddOGqlvPW6Zxpnp+6ttFtR
icGF2Q1hcpSvD6RKZBv0fo2804+m5FyaNYMwPb9woDPWj26PEtdrFF5R/JGlO4h8
f/XoA82UWN2O1SLMW61Q1Gr0eOKmo5AfpTNBjP+ObgaeoR0Xe2h6ftn6OBM/GR2+
ZUHabBlgvkguEG21wOLqdJVLbDGMKfU7oSNL/oY+LCmevxjA3QPvdHc92V2XwoWQ
7pzqkm4cRlg6VZ8WRvprcAKEZgVvoHYrnwK0jcz5SpidIHwEazuKIpeUVc+6j/C/
gMRjOZqp3lBhGUFUnVk0pyFsA+G/FNv09/PzB0mjosMKeT3kCL+9XITIaCryyVko
8R3qL5OBJEo3POLY9wOU5oZmelztjvbHenlXkPgpHA0TTjQse4VyZeQA8TyF284u
mCe7gEOaGvnq5m0tcorCtAf1zwpMVKL1KrsUn8ETH98IetP0REBZKZdcH1BS15T5
3zLB9dn2fu6Sg6rAMf9m69dMQAtUWQZ24zp2yFquZRFWtlRgVJW6RBvNqU/uWxSn
SxZiVu9NwT8q5W7I9FywfV7fdj8bGf8U9Wzq0kImP/thQXOjzgMtXk9htALOl0vP
ESJq9r95iRRYDBSol4BMkQEDJlfvvjTLClAjjVQT+i52JaQs7j4bN4kcNIuQ6btX
hWA9KKX+KJ8nS6+QnXVXeTQdffD9kXdCL5BrPCAXLBKDpgWFwUkOjiwHzJBNbayz
r8JAMK980Rs5sb13YV+xAJFlVrgFUIkv40t0Mdw0cBW+fnESTXYnjiCrd5TJpgDf
SiZFlB7Rq1K7NDw2N83DXn9BTN5STgW9bs8vMgdEZtrR6Pc973Ty7Qq34MGTXV/5
Hc41dybAj8DdW3RdhFkPpArnae2LpjVo8VkxJr5a7LkZddFEwm8fXLQoDlG7OiMi
ZRHFhbSJesrGNrzzCMXw0r0rYBRaXUSzaM03gwX7zyR8QoWkG8TDmBgqQPKGMixI
onVFglGaHUINdQGV6kmSMsx4wXVGNyVn1kOjA2P2IsEBWN491pf4yitXsfR6CHtE
HUuIi6RWoxPFOHhHlWMzARR9b/6AfS3CAgq2kU6Sxrtyh0BGdmMfYMF8ux9p3bC9
eI0W5+se6fHD/lXfcogP8q+1iLWjs7T1futJ4+RmQZI7Sgvs8v+GSX7s7Ex7BAPx
j0OwIjHyYHgQY/FEvrPtLwltwSbTHmSfrGPw1bbhSWF5kOsMzehaKHJLT+YBKZLd
gSUDNIMM+RfskgKS+N8azwiDhR17oYAA3opqVgoeDWGNbCDE2aqyLlAf/9OGSfiy
/vZFAq3FG/xhnRSHpQuvVFWcuo2VP7vH8dTKLaKRuFwJX3unE4YMW6lMimzYepHw
dKiPudpNCvIK2PFKDH3XMxtOMSFcivXxq6aFchs0kIm0OWGog9yCICBRdaJzj9tT
WVtWKjwLquETO7Z55ujfg9W7pDvgbzJpneQMyjxsaupz4oXbcWb4WQefMS8AreQS
c18WlWXc8w/wmPwGxF96mUv+YrNYMd4IC0srMVjegELPPoVO7csgEjumPXWQgj6x
FwPez4u9nMI1LL6Tv+nQd/zA1UMDvyjN0vcSiyBJT4EV4smQEgBvfJ1QVJHVwaw/
wcbWhKcP7r8UeEAO7Ke3eqBuogz7j7ZMBr9JKiTvYcC4RrkfhZvm/iRpdzFXI9hA
tXPU///36aAPUXfMnyaroDTMCc9ZredjiP+xEWQ7s1BC15iAJa1CeYgvAQG6w+PW
UVaCxyrL+WroWuOF3YRpjCDhFx5v2IWQoCSSDiV69wWPJi1JU/yIHL1xPsemHpTu
28IbYaLIiKjK2gDb6S5Q50W0c//3DfXEH6/4X8FxVysxunFhGvMpDaxNLeKxCrI0
Bw6f/hXyYEgXjHngKKqKmw5q6dBPb/d2tgzs3rLRxzGzysYURLizBeW3zwmaOZLt
6edy4DBEcwaXxdI1B99Rnbx8Yjpwlr2K21Fngki8xbDgbsWNlYzMhYWxzplgUCVo
/SZNN+acopqwle5NPhIZ4DthB9yfa+eGYu3fcAH4J/92LbrEowXWpB79GL7uOVPT
7M193GTXoViBTgMGjNOV4KigF+q642t8XQODi57Uoyu4P8fZS5De7M2AEBXT9hRp
bUnSk1OzjIYYwf3jqrQj+uCIhpys83bOvI9CGpHmlctmiN/Sv8wQG0uKgwd6gu+f
qTpJr6lHTdv5wntHEbvHZGhb6/rfYatIOw3anXU6RrSoaPi/jSL+3YWeIsDdfzZG
rylVEzaysCyBXlOxmiKOdmsEbMwyOrrRaPcKwnVIRmZUOJei/O1UpgqOuU/MrqiP
p/d0p8mEsqf2TDVCvzpysGR6Jd2pNbwh8e2zGu3qIf9knln6WOM9T06j0EzvZYA8
0htOzg+yzUzpccOepxLE9Mo363rXVIS3KR5U9fvIbyR8d+GDd5/bvEHvWsgYAjHE
919QQqN0l+r64E+xFQLUGbWbrnKVswyoPrtfduAtjHGnS59ZfbOGCf288qdBVuD4
HTI0qzumfCZFJ/kRsK79byzIoIsG5TxnNKqHCcBqXmrftPXQQWMyoGMQBo1u3pFd
STRFnti7ff8caglmcqQrxrCNKEjGF0LdRBERFQ3JGwyKrhR5QnxGbfC8WTDzSAyt
Sq6qLhqilVUFvbfgMkcxFLveDw9QYxS8NzZTa85RWrbBjUsGVsVCHyY4XzsoQeNQ
3+jeTAVMJwAmchQB7PrXoPbwbx55zX7jPAmEuEqFthIoZqXP8LGZqtqfFc4rbe+5
ezm2+QNCzXAYPSswEH5/c9qTuqM2CvLipnXRCtO/Un/KQASWlThsIHC46VWP2I/z
SbArT9JfvOpJcToR//ul7L0isrkrrc5FU1x999AL1k4lRUGuRWsO8VPACzT5AQS4
5jQ0o336qDOsUGnWr3YdLXajCkEbPRVF0tAJL37D3ySrbSvMSdGa5Bqyb9nxQ3vR
bfuUkl6KsLwPveCftw3tRDwGdUNswJxCEijmg2TA6T16ELsCwykhiT17+lz58L3O
Vs0bh0r1b/UhrGO2TJMvFdDWtH2uGUH+2oeGWsoj4qoCCx80oZfus5UzZDumfWWB
4TOZqSIAEVrYf4QjmAkoRi//x410lMAeIVxyR+a6e4KryVXgzpWAHRjI0ureDswP
tQ71j+6Q5bJVjqbp6Sm+NNelO5akkx1jLfLll8ZQM5UKu2dginIpovJyynaw1f1s
cUf8f5Zg6uxFq6bxyLWHDjapXH6+esSMWMGxN+xF+hmUg49wIBbf6EKW6pdDEVrC
5bZJ0+ZRgtovMejK60+uQvXU7F+KsvgLgweVVUO42EMVijG6W14N0zGqCkt5Cu78
UOJhpU9V1ZSx/9F6Kz0ASWhw//MLajTqw042ycDhOTLyox+SzMaWhf+8dbevaGlN
y45V+cf+Ls/ThZd1NSVYaFibLKTYIRoEth62N/Q+NXZUeCsFPfIBu5qLD76ODzxQ
sD0Bu/mHyCBovNAfnvne+2skRp78GCtbha4aZeQv0jxdjjDQLdbI3cSuAMliJCah
b2ICBuBQL37XyODpMSESfrxOk6mosb/S/OreMzFmPp5UkGqwYgq/xYSOjnARk5k2
zM0Hap8R7Tzvk1MJZBaaU0B8hCfzZk/jCUpZ1ZZGEKe/iI4qEgmYb99NR0caopvS
rQ7zs9N7jOPQ2PAi0vzo+hhobqVBTevrvLofcwBf3bMkBbvJbOGPV6LHpBVCt4jF
T98UQsnAFD2RIOvNT2BFN3c3DiWIWL80hsUAqpGmYrpbhsFVCieImj3w8k93amiB
iVj7K6BhnQQgJgxp+j58yCt2gQME3tl174/dMEVg3yjKwrrs3SRgTZ1dzQGu8lsL
m1DdkPS0CXUgXAa6SwAJHRORh88rfECrdsxdnebbUGUy0PrdZonamkg9ybQ9SoCE
qeixT2oYL9wBDV8GLhdpRAyRhoPTV0wbZPWQNlPAl+S+/RACwqVdB22isHOvrpcs
xY7G9M2rkUhpbjigGE7ynIQzFDkBPmqwkq4mknAn0t6RmPyYZqQ/nQ/HCAmZK3N+
NJeOhaeb3CKsguk7chWqaA09mVeoqWSEzTEfdpZXqxXFGfueYE7SDdmmSElKEpG0
X4XonHz9llgJzOo9Z8RgKyHw/nuH/fB0dMvPNTibUeRZ5Tdjwybzv38xcveQ6HJU
Y4eM7i257RsQTKi+rvMHJx/cPJ8Uvd/KQW1QZYu2vKpDSmusd1VvJxxM35rhWCt8
pZRsrnt1Urdh8cEtTdVKBHAJ/z17hmITvQqWpDp4dl67i9P6pehJ9jUxPL3FUxSP
BCyjITrYlinuhoLJmmwFuw1hADiP3zZXDpPYGgbP2yYSHf9+mF2TPwdHT4+cjj7P
pS+GNM6hyY2iyxfl2l3XW0XzwY8cj9gNbSsHZAw8Avl8kCvKCKNl09MF9JjkNv1S
/qzilU0RFylXeou3Lqgv4WqmlTVV/fTSJz8gUAlVdBMzn4OsLcA/Aybfrs1WrzJg
35S1xuWDAzmFWuYGhpTYDu0gs5C4JF4je341M2EwtY+heGvfOmEsM2SOaby7MKNx
0J5ZLDyjvmNBUeOfwLoXStCVm/9rdBvJqQ0rFYUrvTjxV1UHP+tKBeW/Il9xY4mH
foQIqUFbeB32IUQCWl9aFfecK+ZrFhLWMIlul7RkzIdOwZ/0/F3VgNC/FBshYlYF
Y7v8fH0UqqxCf2wOnLnkbmp1t9jyT8w0XZmT4QJWBUxqianjb7intYSA4wbhtoqu
Ctkr8JZ7pfMOb+MIOeNWl0LWmPOVVDxsFUooCKmkBbPXinzTyqwixUhNedgQ2RNp
IVjvtAtgnzatKbljETq3kltSzfwia9sH8LKTfUdGNMQfmSEbaHZHOko41lnAo90g
GKWkv8dOjLIcqwriF/yYzx0S5LZ/OBf0sSw9vkMBaaQIUiwsyNUD4GofLzHHsx5v
q0i+I8mKFAxbh9jvmnGUbSkU5m5XoX3MBAUaoyK+G8sV5fu0UBmH0LQYJeeNLjYY
6yLuv2WyCU3DRaccT/BNtsLnjVj+vbb7sUjDAUWrDEOEGSsXoaJmgLJk4r9+sXjX
vIqeGCo58OVLD3PS0HX8uFgYAkOjOJQ/OoJ3iygTL9A/8/UAiFz5enUh8dCUXBXq
9myHWJ7zVCEsgQjyJVGczME3k17kLfYRq+dWi+AmSoKPPPkeQF8OQXO3G0kwbiQT
g7G4jHOvtWo1/YnfWdcgBxk0zPfiFJDxaiU2uF7a/ZmjhEeFD0XtpYrFz94h2QZM
xEGhmoiSJjItgK3DhpQx0A6uLzidSqn7AQmRUfOKgfJ+EtZqEUSUkHc3ljl5Y/AZ
XNP74Tt96gNpUNu1sSTahF8qHhBHxcsDverYmHgOn9DFFef3Y948RDCTOwCFVSUF
NuqPe1NPHe6PGqpXU9VU7sl6zh3dOJQ3Js4Cj71Fzmk2fnMyZm37RUGC/yBDKvyu
NwPKkb0sWA2p7ZA98RJ8IdMgsPR4NtTkOWOl/6X3lcGGEGtrkgwyH1hb67RowLEe
2+Pb3MOr7oyW/jLCd8G+0ymL1rWx2tpf584IjkyVogKE0MTmeScO6ndSuEcbw0Vf
IAp10cXT/frkFPeNGBgoTUqff4qHx4c6l0ZKNr6eie3QJhqsKng0g27+DLovOHAr
mxRE3L+BTYdejXDrPZbrJBFEz5jZnwj6zrw8KrZkFD/ckRqHSGzWGuY7V/LGlS5R
orMNO/U+q1I2Ttt5FJMYj4F1Z1kvTdkPwaaqm8gqq3MifP6iPsTbUZTz7gUMpMTZ
xL5f+opA0j5/ApSPBoaWyCwB2BSYNp3UFgjpeW1jDHZqt0X22QHl3TsKKXR0Lo3W
ZhyQWmJfqW6UYj+yhPY6jaSFDuJUGHhj3m73gSPT8Prb9lD3HD3qolF6xvZNYoxH
cwwiH966zKp74er001dCLdAJOc/Q7NdYs5hfykmcv8o0hUOxxyhLdvzg+U4msdQb
yVvhSvK7UsNljocquRYwGjAcJJEvJBFDq+IXcKHmtNTam32Q70v0XpitjHXdyyX6
EtOqnkL/l3oDftOX/k71mJBL96eRPnYAFJ5kOdZE19p176egw2D+TulTv9qxPAZe
rYA7aF2w5WpbJ1XELfQ7gkf2OZxCfvkubeqEjlvt6hFG1u0ngbqY0uLKOASCGb6t
CR5XU0rVM9xgOawXNDXCpnvEKb+WK9QFfXWiU5TLZSjElwMXxEayZBVjwyEf0jBx
odS9Ot2RQRZVeWwBtd23ll1Z5RlD5G5XIaaxMbrMjLHk7hMBDi/FBsA76MUouIF8
QOd6yILoZoEpEJdENHikyp8+jx5VkhyeqIJCu9S4SIJ7ld5kjgBDsAm52w12DNiI
MWhJe0fphNVVmOgXVSoQECd4CQZFb2zLJD4I8CXU0Kxa7frhrcLUMj9XwLMenpD+
A3+jejmjXV22mjqw8AYT9ADSlC5vYIWucHSZIYgOhXJHppvWar8/jSx4+h66GHNq
xuwCfainJv5jel/sAYaL5qh77RyhY2z8wP2sLw56Ic48dhvwW+kQqjMRQBKcOisu
V7J0Lh+XuWI1TuDP18Q7ia8IPyba8PLlj4oP8cd0UHb9/7DGKTv1SL/3Xk+yAzcn
v1YfSJkJmpDpX0vwTZhQovdyOFG92my0+Z9iJx6LlhiXTudRv1/qDGRqGXy0tbUb
iEKn0W76zbPKQYot5N8DLkPCRYDAk0ypR/HI9hSKl8bu6dIvYCsltuQkzIW4pLJL
ypoO+LttlsySYDMOt/osupyqS8qXdGDhzVqSYApiiSqXWz+M3MrThjr8Kymap3sz
voKgb7TGcuVA3ytVgxouZU1BtwY7Pw7ejJZtgMTXHWjJafogTQthuBju2rl1HreO
0wSsI+/97zGzq0XUt3vaJPoNi8omUPbOE8CVDi6RYD1DN4dree0nj5OExdqHD1MM
WunD18GwopVeU96CKwXwqBGbz8ggdVtjRADvWfWmRuSosR06ZPlQj2xDnXx8YIrq
dyR1yx52wa98vmjKKE5rSuIniQ25/NckvT3sMEuBnlR4cGn/QcsTtdW5fprHwFfa
q6gEGkKjkrYxh5W4tO2y5taSjzd4jWT+1K6Q5JJeGG92ZpTTKVF1FyCylertL8uw
zZsApQ1x5i8lT7njDRgEwlDTDG/O0eHANDgSFAym9ysMUBOgJ1k5zxTgEqnHjn0V
tG24c4YMaLiy+J1/msqBZWPSOidmnMxtn/B5TPA8rZCAM2Xt4+vYsxYwK9CbSZcE
9u3HzghEz/BhxqcvOTRIQ2dPVVG13Zo30qB4R6PuLAApBV01DZ2JD51v331QYMJc
ek2nU2RhqmsF/kFh5NkwpjWyaEPXfMPGLThiVV6B0NKLTZ9UKWWDYdmzVRVFjUxG
5xfpLhX7NxDvVrp5mCuNslgOFpDZKvxuAlJzmOiScPy3joFme29Y0AkuiMrmdycR
6FLk6wmJ8Cj6QSOtriFl+0Hh9mdDLh9EiZNnEbSiNhGWqnb+l0kED0xdNRCESrBO
pGnFv0JzyEU0RFa8pILHJriDpcPm8KO/jq7T5H94Hb23AfohV3l9najgTchOn3wA
27JwTMT70KWgBZrEFrrmjxWSVobT56PoJunc2RBZhVEsSpyylTejU5JrSM4KXRu9
op/D/tlGm+T/yxgCP+jB2ZmGWViNmRnIuesGWtDd+RswRaT9beH3rZ9XBvABX1ki
0xS/jIR8VzsB2ChMzhwhrQVlb9yN/3vEiZFcRzp6yTSeJGNuh004JFc9tZCtvJcT
zCuwu66WUreb72CZ3wBV4wKSz9gSu8u6w2b6YsGmVIrYSbg2HIMtPrChe1nqNx7/
xK1nqq1REbvtFe1RB1M6FN/ygKn9Xg0/U4VU1A0UfY+cundSwiMf6lpQQYY9vLPE
JwlS8B4/WyL0IDJCIwx54COxNv4r1CnApRV9tlLkKCmObOMWpHssmVVLifrpcDGf
CIHruNe12j3WoVWPbju5km+pKU7m5xme/gyM0GE77LuQHRwzyux8iseOedGE6Mf1
ihtSvUi+QaEla95vMDAL2GQDOV7LzUId88/6D129v4tzzSS8HJgpfwI0doTuPB3u
DETB2ijXxRjNW+shBVOdInBFxidH6HWyfYRqmGujRkWNinsbXXvkyE96qNN9KCRO
I6MKFIFKthykObuNa4ohRwlSY5P9rjExwKmQCJ+oFU5WgFiFptA2T1dxzwHUDcix
HD1Z7d/eeeHsU7RtfDRUFeYciKv6ryKBqFPz/h2xaSzBXL6EZNAlP6ea08HDF5NT
k7zHbVKEzA7U4aYu0fC4YLRjaPQylPjauTe/yLieEDkYnjXjv+Zf+5qPvK55mj/6
YuD0P7R1P1po/lRqPC9aLH2d9KDrSH9N0Z2w4W5srZ9pVFOiAZ0IWKgSwJZu1IKS
+XvMtEM31ADZcIS7subfFs8HulEVeONE9m1j0atGtMAfH0shAf6cTE3hNHskUqoB
B3cBPmHyoeLzVLIv/+RuTQvAXHOKvTA3Bf8sGnzBIHHofnI6q+ZBF+yiX/4iDRRj
uUcDGAOoPMEGzWIKdx5yH7WqG8SCZZfDAogc7jiAMgtf0oIO+xmUWIUfmGfCjjsA
HNHQrQ/cAGhFYAY1WmGMAbMLn9hrHy/qZNVIqYaxR7ttLdiBeRkyyi1XN7DZWD+x
78GYJBjtZiO62SoYfnh4H7v8TvnqhiwFzf3ljtRCZIIjoTdEHECiIadPJFmXgJcz
Jl6cdDdtZy9vxmcdQKC4miKKffdmfq6cdIAnHCdrc/WS2OHqIbGvd7qEMlSPOHQ8
FhcrLbc6vE+7Djfik5k1i/kcn7/5rUa/vLfeDq2EdrWAZ1FVLm7Vv1gGWAKvJwNr
fOkBDgY17AzXjPUVSJGNuP45aefvUSqqgk4iDd3kcIDhpnsjJsSx+kdLK5/tkcU0
Gfuj+myohyGcbTkOY7Ni2CG9L3PR2Qvkbhaz99cSoGxANsadcwGIpfqp9PWj1SsV
/EzzvH1FMZ4CnkSVOQFDOrQRRNLhVUkztMCZ6yW2Ldpkan7z7RK9SzNskhJQsd3e
WMGYZlziqb4Vt7uPNS/doUBDEctxJgxdOwYn2A7QT/nDM6KQwzoxrGwLozslPSEB
p8EJdl3v4hABK9BQ0txcTG8dHbhAIG0jhOZkFmBunJGATCsTr/vYqSbxvNDKw8Pv
70fNZq1vr/eDp4VcVQvwzOcANo+ovkTlw5rEkK+c2cDqi2zd2UWScqiP16HNdpLy
iUDpd9gSTjNv+zLQAa/IgDcScSlLTYpgh3ydIy08EjVZocAeb7GZf8L1Z1U7LMb5
IxPmV2xkck7Z6fhjXRxKhJSOWdQ3km/FKL7Yxin0PWsa/efjsMbBoiS/00Wxhbh7
RMnBrVCs6j8sUokI4X3sE3qf7+zW5UGp07eOQp9vsSenU/jxqKakWTXHVsn2df7Q
WWwAln9IRruj+nl/cMNT8EivzrHyJElAhGpPAJQLBn6EayMOtMNLaN49c1+j/1Jo
FvmmSyZY0bQn/DAkMvgED6cNz4nTNAIsFoQAVpgVZf8sKZ/ssr4OdgY6i7gS6xRP
36S76n8eCLjj1D8tZEqgQFYV4XodLxAugscR9RCrwMt9vN8c4JGj0L+dE2epSPi+
BZfDolNnyIZ5HH3N9lHVNh9xnfZL/O6DDEYxb6xXjDk0BTar4p6hNyTbEGn3/64L
CceRR99U/nDr8TnPSMeQB05iguw4lthLFdU4Q4FXj/rFw4zZljkEDTje/xkDYVob
iS0goeNpCHhrZNJbFffWVi5ERnwSDHVHC4uF6vGyDhm9fvx1pjrgv6CwBxz9N0lu
a0ottWf8DwJhS4qZR4U/WD4+pzv3Ew3cyPnMBIfG6+dBr0x9AP82I9eJUgVyXAGb
kMVe+4ubji7o/pdJY3aJlkn6uliWI5bHTC7eHZaPr6i2tCVKGZYiwRxFks34rZkK
WlR58dcJ1YJ8sq1pyEBGTalYaLOPZ82Gia0StiuXKjRYVATCOrPbOLJtzhzrI/eS
dMezEuzpsc6Jsagugq4ZJILrdtVK30mfS4FtUyUXMBXHBUGf++HGb7i7NOgnyt/D
ZhpLJOJiYu+LnRb8vMJOcMabcgVo0G8Xk21Iht394zlrzDNZOvpOpNIUDwxpSbSg
ZSUKUkI7npsz6ojkZ+7AS4EnCwdbW0xo0lYPr5ND/eg1W0iTh9WfnrkRMwHi7z3e
5ysDGmtY7JSXRrfGHVbc+GXxmQ5829a5jiuD0pvEmG0ZWANNrxN4sIFa/ApZTajY
cJ7YqbxcoOkyUk3ApuATgzkY5VQtRVj5rOjSCt0V/f76ehFKbWjk0aqxvXqNBfTm
IDrq7TtZ+WZbGOQGBdJE3mShbyt0sj4JfiIddaVGyC9tcy8CYJ8bD/8MsMy9GhEZ
L11+J8/VubbDe3qeR+i0gnebkk5xJp9vkFMfXYPYntxxhgnTFXHNdac23Sl8ezvL
t4Fc36TpBm/06i1ZszFmlfTL1FKSQXfUKVH6W1euzewcsqpM8P0mIu744ew13oEg
yVGB1kQiMuxLGevrUsplWhnVw+LHN1NKVsQ73MdTiS2rFN2R9GQWM2UxC2WiURCJ
kF6EE1bwaHYrODohcQShlCXZ3uEpUPXWhi4SUbVZC7q/EoBcuu9jHC1t/COSoZ9j
NrcqU6osVqNKmqwZ4Lbr1yT2L6DZLr+Eo+2tF6czcXx+xdEIc7yeRw78rCDu7nen
l2IB9ZrDfdNBQG+oHO5nC+qF6TxSPfwkgN6y5tXjEIc5ZtirbtfRS0PykEe3eaQx
JoLYvbKxdfAQbFjnMeXY4gGJgCeR2brMfnhfAiijAkSdgibfEZrc+uMBAZoCqjI5
JqRfUKq3GJ9cmMXDN8d3d5NTE9oLFoHLrZR/VvnSo2PL56tmCHKiLfvIDFyY8u9S
Hjrp0piJTQVogAOhoKprnhvSqZq4I4JWGHPQB4vauAO838wnjJadvblchEB/zakO
xKhcXvIgbxvNLriCd1BZ4EycqUFjU0Tggo7cidmwtuxKretkyRFerqYR98pXEL/c
SiIJS/09HDCGWakKldcytNXc3SknqZHQNVfW2mC20UvrVGxn8R6xovu2mGw0vjFn
0/RVp07J2G5B7mXqFusJ/S2E/YEViCUCEY0Yb2ZFySHDG+1b/ytTyou3F71oOo0j
9NOwNlnk65gcnFddd4/npUAPAIZNUDFpB2y3t/HIatCgY93U6bHEw5kBh3W/Da8x
5A+N17xlxzMlk25Np8J4uCWG9Xdeo/thq2+Gz78sgYEbq06rxByApUFp4caHaGiO
RJd0VfEaPk/ci31TWZuFJgFHihMa6vPy2A/xyPJF+ISNiYuIm5++Mk/AhUzSjGNy
xnPi5+43/Y/lgfZmBvmnNt19Fm9ZCoqys3f35Xw3McwtQXQZn68lMZkahhKQzMQ8
40fr3wPMrYl18zVTS0EvQ8uKDH8cQhHqFHj/t+sTZcwgSOhgQ+zrFBO9HFObvyiL
JY8sbwYdmD/2Wd8/8pOSxx2gfy6rFElsRAsOcen0zajLjRLLcbneLLYzsS2vwpvK
gvE268RFicZPgTIfN9XOO6NwXMm0IsVvVhEJ+ITjj8amGkbtOpB19S/OGWomMpUb
XmHpf2baw1I8+nVQp2bPTtBUm0PRXOtb9bz8jL84ovGMFQYQflcsCgSNSXx2zfIS
zdEHeeS+nI2BaUysx1BvJJmTG6WwjppfDMPsQuzJMIx4wmEu2eVLK+m/iLQlnPOA
MMgy/cgrceYIQAyFub3W/rWZ02Bn0n7+589ev7+YAUTRjEMy/WXLT4/cr9E/6de8
LSIWJT46BBe5ibO5RrZK7/mPFEIMrTe5HOEYWOGxcm29VOVQMw8fkp6BgnwxISz2
erKsvvfJsNmot4ghcs0BOIxdYZZBNz1uAUvMLfeQ1yuZ9CXAVawdI4R23L39dhP3
gBfBGNoYk/qX31BkO1W4liaP+Mh4hgTZ04dhgJnDaEZECNaOs+14+v0eNoNGXNJL
Mqn24cEGvh79T3MAdC99U+V3Fw5IucYBp+PdKdvr/6UJ1QsbrfJUDuGXU5qRjZZR
G879F1ASBVLkD499iP2DygRBEaxcl3AmbVFUX6/EUzIyGU3SWQUV/p+uTJIEVqOQ
NLlPg/iwe2aGTtYEPnCrsUSdiwBl0tZ0jUjnDSrF2YtUXFPHq8vWmQvnSR18ATay
/D9mzEglTUpgUO9nArH/RMjGeOxw8gQXJKqhFlaNRtcSUE91EHcTeJdaPosMgvC+
N0cjDgg5Q6aIEGWLGPap13v5j+wkVjoZC0PQmmo4AAT1pz6Qicx66MCHgnBgTh0o
o4qbNOzBripPB3/d6br/NWjrFO1KVjOjMytirRvSv2WfG+tjEthcODEYpsmwot0W
HZH0tBx1G5id0N2XdKsmSgQ/TxJdov8sb08nJ/hVTQPE85My4QPKfQgRh0OPq04A
J9/95/2TTTso5vh0JaIVYa9kybygZTlVUXwbPrI342dVF76TZFm1eL3Y0BJGXawH
3P4FsfX07fRutLcOFN/OQZTQqDkIF6l/LyMR1ZE5ekFpevnCKljfCbHtMAS+5OzN
sZ+XuId/8t0W7kHHLpwCLlD7PO2AvCThoSoKLdyuKaTGRNtiEqf9rvfUYilWEt9S
41U93sgMKhI4PJLvG9aXBv6jekQXQBsj+WRunyJ/SxoBbzhfGPOzHDpVmzxGAcl+
mm69wFgvtljymhVrX3AfdNVXmI7XFuUuzK8OozgesxWJfurno+DWY8UFMnj+VStA
5izOrKGhineM0bPbYYjWr7fUQUm42MoC0NTeXgztYyNVjMPcwq9Rfr287oP1iury
VxAWz3D0CLd+UnzLr4do8oSJOzt2AvtNwb35lrY0BwK8KG+ZnuGC0cdox7rE+euS
Y9lNnYQDFyzG+kmGMtAENVOj3nmIEk61U2vv06TyzQqvVdlXbxUZQubKE/GZ++4W
SLKMylj+q54uLFlhV2BisvOnZzSdNmulmndxkkEo4wnha9nOtcr88EGf4SXGOej+
V77EhdRKpyxKGvpzFopub+PFf22PbjIAsyDTZtqvn7Q9oIYOhqLZo0ZadYWnkJcB
6tDnvKkxNpXHhFu9scBskeZWRWofqsDyHrzrnKp0BHeT+BSE4w4LTOYOpA6Y3en3
qae02SUpeUZKNyqyTmjY7Kv2IkihvIrG5fJrkoe9Fl8Y+IRXCWt803u+mQK8iBb0
kGlLYkv2VVdn+3tcdox+mNn6i/8WAXYkRuak2nisOBCmkSCpjfTQOJpiVMHJtxJr
dG7Rh4L9VGvCah6NIM4NkASbMb0QUfiET4wzLUGDpZVJll5oLcr85xcQqswD7lh1
nhoUbSAPGV19eo51QhB1/pUgJmX2dbSUEJdlrO5peqbkRVZAsA7MZfQnjN6wTaqt
wSF/F3qOiFp8aJdh61w2bdhAHBZ3KltS+xlHDPxg8JH8FqeH9fTGmpq79Pv+LHRo
vyqbX1IYXT7F4aw4vLyJhHpyWGc1mnjUayvCRGlHm6db54UrkD6dL90F+Oy7BQyW
rgfLbei7Lt1NDrxQuJE2JKmonT2AjwRGbxuVhru5f7GdUc7kO5x74JAL+T5LCkZy
7cZSQRM8aIUTCbALr55AvKmeFP+bYzDeyV+nsYJTwV9vVekxP7KDpYOWiVrLAWA/
zrZniMIHIhOiQtLcnNtt48wS8Ls4eekSCUMFh76cugwzp2W5P1CXc8tyWW4t7kKb
k+aij2Jj5YY/BauleoFBBBO3vEUmppJy8OkqczxJod7F2HiNNxcRZ/V/vXhiJXQW
ZqOYRNdbzgdW5QWRgPYDuhR1qLJO4tFg5DFPjOYdZ2qp8KlqDECpfnRoO2x4xzGb
2O6/rh5o1kox/inqBLKbueKVFUHtaimPU24MOiqO6yDOZKsR8oyYblKDX4/So/+b
vfNTP+Mx23zFnCYktKN/Q0tl3yZqg6XWHIKQNO/DhRpsZETIfEHvQH+CDcXBvZ+I
1wxVwtZqSKkwabR904DADXICPmnVssORmvOca9S5bE8S8G0RMFBINurt1igaZtWp
Edcyw2dC7LTUiovlSFDnx5obV8noAP9HmEgef+U2SerljzkqUFTIcii4LzHGpkUr
45TG/0lF0zuccO3OWLEuzP1dHNPZ6aGMPm0HJwm7bx7CtZj27MmBW46TIfrPbVlU
P4QO9whOyoARXweGg2TdAX6fCibDQeReKg+K4KyuxozqypugxF2Mqfq83CZ/uI+0
2WrtG5OpqZxTfMW/aNGO3HqYe/C1F6+XutiRkJGYXvsm6IdGXrQRaOI8mDVu25xj
95ySEy1fNbwRkDnfOdpxLSeKAw0ShUO4gH6t4XrUgfX/R2kYoUzjR4VZdqQugpfM
E6qWaoVt1rEthQ3IJdQhXd9SY3RlJfGRJ6O3LZCxPn7WzouFzoafo10BDRCryzeh
f7OTztLHsJyQqu5xzyGgyTTBwzUY1GOhQGVwx7e2ugMnKUJmCPM5lIUmLYNjzF+7
/N4tZc4kPc9lXPqcoL0eJJ0+Ur8xBt0cgTvtDjraxXETL8Ycljd2nMeWUxjcITw1
n3n81yqqJX9ksK/rpSgzGMb5AgRfVfaWan0iA4li3WbYG7SMoNReml6tNC0nYeP8
QA/fOJ6oB/ji1jWY9xAp8WOnrE8FRw9nO1EFZAkGj9/njr7z57KDV9nqDiVZCg4B
2sZ4OmeIDFxkctCG9P7BJqEdHoNqfC8S1TuWQ1oFgAlpJOKUpbYERARPDApwOPCJ
hmETuEpSiLDHPtmeFxkCBPaByZ1zTV1pIi+c6y6z0al7FKbUZtRKITGXziTCC3xk
qBD0luwHKJbOYQ9Ych/rAojvUDhMZFoF3So+Xx4GOH3xHid9Hj2vKJqk+YwmFz7Z
arvEZnnktgse9r1e5sT/cIhObNMCeqgUd2RIAjyIgF5Ldl4pOV83slF+z6LmUSRY
0OJOHnJON/WG9E3tDE1w3SqtFXR30/oMltN72b7wk+PoeO52NkMltZclS2AeDqOA
FBEBGDs/sXFOEMzjYFM46Y6kia+6qPxEUhPXqKFxrTHmy7W4Ke2KRGEoRkrGE4YK
hvq5i2ab2pr90e6upWDpQWeIkO/gfGMFfEM6Thtawok89WadkCvDgEb8FevfSQrc
KBeoC1qrkqty0YhDKxj4tnCjht+C8XkQM8WFCAkZzxpQoEOz3hFLbwsn6C457ZVg
uHIrWGPI9k9jL1eVL3M5Mzrg2ygG16/bJoSImRKq2e91JZNsXFPTOFwJ2cHlZyQ+
IM0tCntIUd7edT6vJUiMQF1RMOSHHwKJhQuqKMmzYbdxwwZ2S9PaU4lxV0+tE9jH
+5N5/BzeuYgJ3T69X/z6jp/16jEwMDrC9pDGS/5s3U8DCvlYDyJYMCnIyuXIVHKy
+7tr/4K57jjHo0BF28YnC3D8j/tEvB4+0OOAqUuqdm5QwywJtkaH2sRYqI2r/+7z
tD0cMi1Dny8izK9d4+9VqP9Dvbwkxi6nt5rSZcDDlVvf7OTBEHsJ0HOprWOxhf22
kCtySxbulpHcfn/2ZNBmU3EO2bLFI7Lf+4DbbMmhw8aVaBDCOyLVNyNtgCXcYS1C
B94mkR5Nh4F37xFaYrMYPxLEZlDk6tlJGTwDfPDBz5UFhMUh95ocdDQ14afM1gaE
szB3lsjbzZvUhXFp06APG/9mOOy/cyJw7X3CmoDNp1vHUiURPJUcT6vQjVb7LFdK
3iFNOCfT+xyt+2UoBpeefqIAp1R7EuDwFUyG8VHCajP8yhzr2k8okOTQ4xW4ervg
wM9CMhLSZceHiZ79/4c+DLa9TKZB+oSB6zV+nqDgjo3QfWuVqTj32VVIrbqEttxD
69luGjMhm2BpOUbCRZjWxGrFASfzq/ViMD9sp+8nijvukFyMYLJcDGebYUGqdygb
Q3foARwaS0IFfp555CHzRcybrDEVhlITw+CkZZIcboQtD8ev6g1/5Z4LBBmLCmyr
2a6e/3F91NUqL1+pUpEBwSgHj405aOsc1KxOMzU/BXz/oGmCJ7e1fcQu7LX0uPI5
sP0CxuYacepDtLuEYuo3NI9buRaCUlRk4yMN8jtFmjbH9qcwHwdXrTxH7WsyAbPc
OZtOlfP9iDnSJdIysq2yS7mZTuvgeDq5csTDW7SGPcKo3sOFH8wv0BQIwC4Svy+L
A3qdWYlLnnke72JyzmKSdaUNAbQA1iA96E5Fa6DXwCjwZ6tdFB2U/IyCnpLP6q8Z
nt3LU4ZH55j1fifCV1NNyowjnGUhd7hR+F/r1v68KmGgQV1wxnc01Fjg+dNkuEYm
rDmnKCCoAbJzkUAT74zJWOlhldwhx1rFXvZ8ZvgypjVfEPhU9jPVXxcdFIDCLmhL
yEuXkXSXn9MoA2eaVei8APKi/a4d3sZo7Le/XrzTrurbm625kFqjN7Vq/A9Css6D
QCOfHxncUw86MgApup01H8uB0bQYAAl7/Gf+mkrWMnQSxs9FahTe15GR1qf6KIsy
k/MuU1fCLLEDXy4vApiJA8vOse2zZ5hJyypYbNSSg/4YS63X2NBNhFijFLDaAEJ1
CxldMyQ9kuje3nLbFD9UjzNCXNQc2FySiJnAj1/vWZMnNi0cKKFA/FG8vQliq7wk
uRn/+MWob+yDga02RYIB6N5YzxSX84ckaAxw1Bkt/yGw4l6IAUUtvHPon3w4pq/7
/9mS9P6S4/ZmXjn7zvIkqN2lPz0GSxO9t2tzBI7xIx26hX6jk/DxDxRtpZImci2p
wcNyIIKDmeHKDtZakV8bu7ELh1NlYydZfHHupjw12EkmFalKk9QXQhN405cdgX2w
JvsswZT1Rf1qRCou2YmVUD/kGf+tp08D2AxgChaDxa/aoZH3oINLxfbGvF4FZo1k
+dRBZGKdhxUm0zq7sZhSQRsiknFhEIbdOch25VoNm/IkBYzJopLud9J+BgRm+NTT
s9CFpb4XceRJvLWgvXEA5hDRYs+EYIi5jTlurlOhUi5q6X9PiTTk53pFpK7lJsQl
LhuGIcbugsAYpRtHIWUkVHR95gaqHrNedrTkNwD7f0wxiBYCMrfwkXIW7xZ9hPhW
2P4HUPqxDdN/qkMtuOnsHYwp8NFIsT6oyZTQiSK5CnWc0b5NtnuifaanSAvU6G7A
3W/6EsItAlA7T5/8PlX6vPbeul7yqmwuhn1HclOfvnXcJbsUXq3btAR+HLeNc9x1
CA8DRlz5l1aW+i8NhIK0V0iXrXAKUuC/jffcPNKwqVxSDYDGHB3z++nWWuuz43xK
7+J4vBNxiJ+Yy1khOBg4ZxasuOx79RARHDYVq8q/2SyNcIrgTbCFJAsiQ7rDHZiM
BP4mGRh2yQ43qsMpGhL/mWHywZE6GVuugKeJkwgQ0RGkuLGpr/ZOOCrYooMSvyXd
5DkEBkHv+u6k2FepQJfTU2N6eeLByB0Gn/6h1pHWV9mpGZqRezGgyr1rEevDRcxk
cX73zRlBICVJMj2fD1kFLm2hq3ETfHOJ8T45Cfz4+8CvaqaQqLChgudPmlKKlvuw
Fs16zBELPEAH/pg8O+Q3cYZ/TspZllJgvcqYf0fu2wxqD41yIsd0sdPot3oBg/i6
i+f+HxscsaT7ydABBIjfy7ZeJgKrieYgl4UXV2hYqXM7NdTMCkWTqA911erKGCjf
fn1TzsOPcftbByV69sGLwAMrkqCsuFh7X2bp+APaOHVJ+8g9QWk0yjm6KD0BW2PY
+vYMdFPmhypb7RAH/EVvVO85Zx4V4fAh71CbXmgiuHHpPJ13EOKh6nkrZL4zpi8W
1KRzDBB6zVBEnQGkxOspn4xtW7m15RjBqEFDEhMhC54PSFdgzwJTMAFcKqYOv9d0
6QhnXbqTufgqRmzEo2ujbmSKS40WFTvsNH9YrAjH3zugLdrJBhwkeZiu7y895lfV
X/RKii21sRtR/uhoseRwrH/UJNfNDBWIuEXgSACDv+g/c7MaSmeYJtStHdLm7zOg
pOm1VQ1O9DAlMV0eSbQy1O0bIqIdPqjZv6c++LDnt0CpWgB8v7PsAgVxgO5Ngisw
h7A2I5m+82StWIqnPi+fiosZ7jSIOtuZq6rDZqEdKRnrY8oIGVYelQoYGvwrXy3M
opNT9k4q1zyVHF0O8zyEtgT5OHKUyFKUlJamJvC6B3HCoeQtygHgsGfSduKmDzVM
sEKVZnbs9SMfFHxPKI0EVZ4RNcoO2GZ0mmlNLHZa0o8JcuY4Hhh4FY5xGsOygOrG
plGyVoI3GjgD/5i/FoIOT6bFiive3SIjDWFlCUrR+3fMr46w+a3IsEuVTtYcfohy
mpSMnEHz5Yb22YKkM+OZkjbGihqZ48Zq7hmNpV7dCHSMYlUwWLWK3xIL8afe9YT8
pt3sw4Lnq9A22JW0LjV13gto/h4fpndrITAZCtFB95tpkGHgmgYBBxJK7X7YFsak
yKBPomjiUHK/OFUry7MDP6rJKPiUJvkFwtbUWLI6NgkiVPXTpdT58coo3P0HgmG5
w48B84SsBEM/Ynd631Qz/FLQ11iNALEn8Ucsmvzegu0n94yahBqnB1cs1eF56OEY
C367TQtta27cgOir7Bm4ECm4huNs5jha3AuwQ+SD6f2DBKclIv3KQflcyf5Q68hS
X+CpnZSLc8rSQ0NZAyxH9h2UEsPwuLlZ2xgo6qQTreVO4/PUF+mZetdZCvJ7gY4O
fbiHtHu8HwZanv7ksiioB2IAmFp8bupKuiZ547PT/yvghwfz06MNyshY2WdqN6Oo
iKGx9iIRr/sK1Ze3uHswzPxipzzOycK5uh1GjWks6t0K+AiywylVAstg+k4gw5tT
OCsrQe1DIRvmeXJEpyeaWyfy6L2vN5OfOdv7Yoy1S/jSJzg09dOFXHR/IohTpTdD
XM6w6JDU1EerT0hL3mMAGimY5+U5h2y1z+SjnpMTc+fDytWXfzxukEjaomqrZy1L
E0oY3gnozhiQLjZbV8S9FpnM2ETJmD+wgiR0z/vVDFRc1p5qTK+v9KFZNbwAI8YL
vuFISktpUYbrhkIY70rZRgYsYcV6LyGxKqKRWyROd43sRnnXoIqPKx9wHkljdmhL
gGnBtEB7AJ4cy4wPHaknBjMsTV3xyScu5Vaad5dVcj2kADzX6r/3VttzXxR5fLT/
Su2KHiU1MyVMoFlvRsbSW+lN9bV2JrrNBnbkrNT+V8N9TWtHlt9OrKshq+K+8Eju
hd70985wuIJ7qJWxHrTlelkcJkUVP4j+y8lLC+qJdORMSHMO8MfHbRlBDQF2YH0x
ioRPFpKwe16Tf9F6W7SnoYiLbEclfWMX0cbz5RMn9/XQAS1HCEWN7S1ztNdpoXX1
UAtcJYPHSHsK3Bvc0LRGqWv+r2RvddzlXuXtzho/pTl7ZRcFswR+T2irQ5b481C/
rlUKetTAqTRuKWKVT26Dil5sjuaSbNH6uvt6OzD6pCUpJ1e57mW3dxCeOe9oEqgU
6EpUuFuI7xdkQcuolWQ/FgjPD4evmrDUxL7RWQvSxO+o3r/jF2KY7p5osYbAjsEL
3oTptNP7s9B/kza1JOgupkpQKu4qFECPlsCzZv33B1ESAmE6lvUscynK80Ynbe5V
/GGcPJ5zv5dkBmv86NdhnakJ+xZrPnzB+Ws320GynU6w1h4HP0sneE1VPccK3P1x
9BhLPj/oai5LKcNXgd3GNKke8WQROEgpopaP6zKIEf/Xj1a66otzVplKLjH4CXlY
jbnMkTrjJTI8boyMT4OOVeatLfZJX9lCBnrRdTssXBaFFMNkcBp4FziZ1uy+ueo+
P8TQAa4DkevCK+4Fgn4U4g5249RnTaudoE8Bj1G1p90He9OHesDjgN9CySpxgR/7
GKuslOWGOtF4/ar7p5A7MVRhByZ1mJ0nE/Yhi3eh2uoKJGXBsNVC/yywUHKVJopo
KacC0JCqPcaGOeP+he1k1qxgMOEdrBvQbcgmEqdFcGJeDXl/Sy9EkGD2iCUXDCLR
2JqgnTx5ZRvK4ZhzA0tcfRy30+Kq2/NUGK2FoG1b6KIu6DbSNjIXCtpHkm3VofmZ
V4BIXqEr9c+laItaELlZuYDEe+H32JgZZZqPCn3IYML9xCN3CtWUS58o0qjmUK6g
We5UvXePBgXeCGz9Uv5Ge9NPF7wmB62H7N5CwVe6llbbFNqi1btDUrHXNWjj6ahk
AfJM1ReBvw7fLv0kM9Xzumki+qFeiYriusjvIIfDCDYJgdCJ03VqgIExrni37tdJ
WaX4KoDp2qookr10WiEOtqoQ97yahDWr4oqElXxTgK5hST30ULrL/aDs9Xz82h/M
Z709M79pbq8iupBhBx5isvw/HMfiOYixuFT6xNF25ViUWxcJ6BOuxO1QlE1JS0UL
uxcvVczvIT9XBGkq0U5b51VEzgQOy1UCjRCGE6H0OW5wvRSD7+BNfcDFUL4yhRJc
xcGyTBNJa54dyXUeOU9KaND438BuuhnCMY2f/TJgAJtjAVJWh9uN7b6CF3Mb+Z/I
6wPEJjDiHZI065oeL4Iae8jc1mc66bkVI8fSlGPYmRTcD1pqMNvi9KlzqxJrzvx/
R2VU8miDQAxFqvI9oYk9mK8mGImFrkC0hda14lhRzxvpATwKHw22r6QdqTDQo1nN
QnTBdWjaTTsLwdPxwK44Z36nbMlaRp/w/N723dZi7TKh1tlWPa7bww6wsWIDpLg2
oqkP79OutlpXY9zvN/RtJCAFuemFcEOMWBIvk73fAN0X6hr899CwYevvMZFB3QgV
2mvCelugL1jJD+RU92tSYJTZ1hg+n3qe3J25Yg+UPjZb+31f0GOCQ5GHI0r7cPO7
+oMndkveXy2s95FhlE8CJjgvyppEw7756FxW23abkVtkr4yyPYUBBOXldy9p5j6L
zDWfMl+DlKHQwcIc3fn+29meV5J5FKhI4IYvg9539STNQZcdyWKXgt4VJgzisDIT
38siXKYs8WV+O2gvx+rxFPTsGH9U9d2NGh+X6RVnltTDRn0leSE/EhPIUCI7Lrxc
s3aa80aLePTgft9F8G7Bc6leF7CmttpKsYY+4o9yO2H9F05915/DBd9uVzVxSTSz
9sk+brTISBH0juNKEaICvDnfZlvuZjP6dSD88w4W/y7rv5Pb0ZDiUHsNwY8MjwP5
Txt/0TGHKYkIRmFRdnox6baFRErnGpe1htDUPg7CExeoe+IjIUO1pEsmHtA4g+YZ
Zi7XpF9ayvitztRJSXw1mu0VZ3kc9nxb1ivDAXTP9TINFSKH8hOueQXLsxZ44WNt
gjlFtyC/E3MSHEVcQvSKhvKNNonOOObTpgPJWLZh1rLu615AU4+uC0YADN8nX80d
yGhQKJGgbyCkssjJAWge4rxRKgpXn6yHNwhmzeFWGSfnpbV6cC6hqM6xVtPZI4NU
hdnvSFE30e+CwAlsu1iI+oXGTblFLW1IcwwKHEbKFQTDBT8WqpAOOhEKJstfvS8I
xoamAcBbyrCUhrUXJQHCucK+2yS0zsTa0k7W7bpU6ACWJNqPAeIjoeIfTKPBGf6m
rSmKc7dJ1mdhs2v/MTV/Kr58VdQ1MkuG/egWl+VLiX6Ds7UMvXxSJPDqdJS3BbNm
XTTeyZdwtFmcBz8Xmc745fEKK0X0zfozYW90Vzg81LbB5WvUuNL4POXOMD0LHUEa
jutIimvBkm5jaQSBFI3daE629VB2thdw2cTo59wG5GBObwvlOslMxrGOXelTp5rI
Wv2A3Vr9CdtZ93vm+jjwjd3zUfCno2Q3CS8V5TO0tPEIZ1R9yrYn9/JbAGaXH0u6
EHAzQ7FVgGjX6bj5rYP7mNwhc9laROsE+lhw/GAnSa7Uo7mY2PBoin2sEZo/jwF/
HqVf/0xjK1P/wovDCKnTB9YL1m1wFujpGQyK8baYEaYOWZf1fuB9rcZAAct9yHEB
XZmn7swIhUtgwJF45/v7HHiM0kxNt5IYQApIJs8T4Y3W96pA14hggcGJKHmSfKbl
PuYSl7FqKujapm/Za30/X1Hd7Z+Aw12QNbj3adih7VyAD5PKIc/WiGVLMJ93zUfQ
yV7Nz5HV4s98ULPREPKasNwevtw52lIXDl2ONkmQ60mOM8GxNHp6YgHpArI6CPa4
gSbZRlDU9/90LD8Avno6gZYKLk+psZ33iGKLb3JfueSqDMp0UW1G8INynOMiz7HC
5jSpgXelUlkBtAlvKdnrwZjcgivVCZgyi2QVKiDPRHYb1rz3oZ6ffMqu9yHDkED7
z2BJg0UwFdnPxRKv8B4GOy86jMolcuUWnYHciD6uM+/0Hrw+J/RfaZVgW2Bo8+Up
4+taYzsKZHaJSttoDzPtQhHtHSQKOCXqU1j5VJcEx5O9UEH8eNWqfvLihdzW1+dq
R4yVd5VWTR6bWufc/SBBNUhD3wmlouyGU4E+M+kJgJ/trZdiSxo/jAg82ELuU77d
WdScWzLRIuol/UPe5li8LC6ISLNfkNewTFpqvVkp/f9aWMtrkL49KRSXtaMMkAfh
EQXZfjMisNJBeG0QnBkksrNhaGr76z0ALS5sreVicAZhgBcK3g3K9sNrusMA0dvA
1f2oadcXox1Q7fSglMAa5fem+kPtyBldsm5L7otE2XP8NdKUVetdbwGTyNFUWeKf
IyT4CBngvfYXf3BfKLsK+e7U8T1q2Z3FxofY1WeZXHKhrwfyS2spDRiVrmvqnltK
Z/UkxQHWmubHZ0d5n6CvfFgMDlEFz5qX1zcHrzJPSTKjN1nvQmHxPJ5FypT9uGG/
+eiYOD1/NTYUL2Pah3lj4DOzEV/OBoWWSCPkd3ZG7mc4nOG5qvb4QeD5/C2leR8v
XWGXwCOzrzQ0b9CxEGHLAVkf6YBN27JIx/r+vy0MlS50ZRMFbrgBLblIAVeMCWWz
5QR+y+moL7CuICHVFDGKgRrqD4R3vKvXabejScyATfZ/X8Bj2RFbkCod7CTrSyHI
ah5pQ79AH88auW96c3+Gx+Gnh9pfI/DQIRhGXcZMQSD8FYh2L0VZ1WM544oTlLrd
m6eTvcF429aSJkVqDUAOh5TJ/7gb99f1OLOYQT5r5tz8E/jvo5rCGvPeyW7Pk0G1
maUl6aghjA2iF5YhSc+9EiawieSU55vBSjjCo766imxbh32vvl4GPBpA8EBkoqHM
SmJPVXkUSyDTI9v+pSdX4qVgqi0C0uu/4N01OBbN2bsEiHOabbLdfEctj7Zdx8S0
xHgA6scGYH/ChtX54gV74V1WWhwJ1BrQvEm2aOWrhjI8UXkzQszYb2+PgvwPYJcI
KL9MDEDHn13llkTxXWKuA/N2Be6MgGtVj2PALKivucmtlDyeFiqLCifNmzUlBREI
dkomS8li09J7r9sk27nF5WlZxJaUXpNaOhI8DzNcPc0P3AthkbFWYWC1FtSqC8HU
dNxsYK+kDyOpFkCLQaCtDlBfPgmDqycwFGQEoRTG6sAhQV25aSl8IhSlsierum7w
c9sE3OBv5fde6YmZnoLi1kw+veH/BCdWQv099UIPs9AwFqvln/9NQ4KlJlMXIy6f
ey4RZIJSYBQH+LbRSJvYpIQ2qSEm5R6/32VCKMP337WZhE49tpLO6LyKDR4BUyII
EM47XozXDurLOskPoov0O+tJgm1kZGOgNamgVHdwk78m34hsgYWhHwn4nXT1HiG5
TdVjhUurYsOTuaUGbMYxQhAxdaj4z6S80cDZ71Gw90fVoR02YdtNh8YDni8aQbPX
iibdkzT+Ut7KKEUy1n/jWytLqxk6UQeDV4c4KZtLil2i9aOB51yKjOzWo47dVsB3
MurkY1I/AR+wISbcgyQ1yA+nkSIGY+1seCjNfqL1+w7vBgicsXMvUg3UBN52xAaG
EEYiXT6CKk83DjCX5Rd0aPQ6nWYxBkefn76Ri6zZpTlmpGwhWUG006wwHJq02FKZ
KOutw/btcQAGZTMFJKjcy+aIDi41spAa9uP4Ow51k8hqyN5yKFrTgTa3yVieQdwv
Q/YP41PNXxEhjZZABqTCR+ottZKqb5HySsgci1RWKixVfgciL2t3qv8731Oct/hY
57cJGa48l4lwyqzL0k5fjEVQOIWso+5Qm8GH5FEGzjEqeHvRooYcZlutJbYwAqBm
P4Avv44wX9Ud5J1akn6FNnnWCbEeZmzHQmgwBUFlfJI9X+wi51eUjp+1EtHv82BT
NIqSc7StQplTu6xRkWNsPyfvS8311ct8LnA/1TNv9ofbb/e1/ISmVFhXcdwnoTSZ
I7fuD3p3HPHU5KmB1MpZpig0Bco6G6QJh8Yl6DFSuHIhxc9eDn1i31FCz72/75KJ
U8m2cQArQARZuM4lBvVKiRgCZhcTU4f9xQP/Hyc6sWDBxhPMip2hPl3dq3RmbdVk
JzBJYXtkE8c/3hM4IV1SfulHaqrUYlK1ek+iCkRwQXkB0lvnDFa3bKCtQMzSeDDd
ExTmyL6o8LzSla/+my3defN7yH4BpPLmxjCmb9mLDugK+QqJYFfBBb2pbuOaKwEg
atB12cL7zIO4SIVzRG/GaU+1gk0SRGIHK3gt/anXjVdOPdy7jx5gKv8FSL2wCCDj
Wm1L5UkWH5zrscgYpmLzLc4rx+enszPeThO9oxzK15daBP6oT+mX5M0sfVdqf78a
8kqpxoxSi8F/nIPWVziHSdtCN6pTJ7Ttj1XXHsMIf4LFiQRvZ6yUgE0e2+0c7PuV
xze+O4TojVIIXjzLBBNCsmRjVK6/uZuGKGTei4hzYIcDz/h7QSKGu3dM4u3qAAjN
jVjhvpgeKOGJxqy0F72DtCZO1uHjumla0S4wTS9VYEZ/0OzKNEqe0QOW9LUbXRSW
T28RIGOQIL46HigMrsUxE53oVRXSs229xdwvDYfyLvgHQsMdmvmV6+d+VrYWh/ge
bxUXdPWAIwEgK035djppo/CsyFZVx3EJpjNwb2CoqsYgKYkyimEsW6Ez/AHOstEU
WQ5k8iH/Z6GLuKA6zq2zb5vlHUlasah8vteUROXzU+eJfWkaiY27pDk6Zq16xqS+
WTOjtXninpKZemsu8TW//EIrfCAPJJdsuW39WiL91TZwCV+4455+Fu1/71U+j4IT
kmkamrFmaIhnMMhfDLQ+I7jSuRqEjpPjnXoJpMS5tI/6nh/nBbovim/De/eexzdL
hb9aOV/sbaD3OQR/+IG4J8ahY2yqyqhd07mZD4aRxw4M72mj71O/Y4g6mUIpcFDD
FWNHx1/X9TEocISCgXleBY8PAF4Y98HRZO3PrRxWxfut9C9bydCk0fsP7OLx/LbY
p51AE1kDHbcephU+NuPVfBQ45JEluFmVmndDt5mo4FIM6UmOcaJ8F65cD6TeEffd
4k34nnQOqRJ01nElGeONIiy5+jLsUZsFbFDGeuig2s+OkQh7IwetR4qZy0DvDb56
avBUi5iO4NX6ycNLHigNGNaVp0KlPPNpdtl39tfQYs/2OXsJqYFMx9Nusxt1+XgE
HC8BcV2Smo/ftGVaMkW/71MyWPvHLHdETdjW+f+v6iysWXfk9gxClqZGMEXQdIwu
MrsOM3XoYKWjVGjwEWI3abnyCZ85LNPBB0x2iggqHLQD15MgUfm0BP6M0pywLIjH
DvcZHNgsaJV8AfNgm2gX8ZJjC9gSCSM2gpO1U6xXxGNt/NbjLTqZ2V/58aTnZGC3
7C0JBCLlUDAm8B95xUT6HqEeqYOOLT5U0SMrUK+w63X4anuqT9jns0hFSyLIAiRO
I9dOWLCfApOgh+1NGJDf31ToTHVNeel2sLv41YlX9YOMk9UUr+3FDbPHDz5ypjAZ
zacmijWTEHOUTQOj4NnnVOuCx1R+1kCjA/eZkPnQd3WOsZMQfnvLZJDX5eNYFG6/
qhoyFZhDXo0KQsFLUWiiV5cto7xs4k8nPM94b6z1kY44ARuMALS7miLzQDFHQPc9
oERWkox6K/Dakfs6gJmZbaQ1LsAEcsQRRn/iUjehKWrCNkrFhPS7QPRuJxC/1tgA
SagtakBY4HB61FX9qKboA8gZCcQkiId+x+29UciLNUo3ABCKTcQYBSJJ29eGQjkw
2bsqQL7gFqAv3BUaWIrScDyjn9W9TpFMVsRQktmwf4wn3GLSMidyookSculsfuIH
5ET9lB/KAraILjSD7ABnJmj/E9nZBVUr+fPRom8MHAbEm/JWU/HDrb69Zo/E/GGq
JBYnd4i6dV9XTOy271UQb/3xzrCP9/1YHb5eEaTj3AXTwqPhwR97Faqv/TMJRcu9
GTeoBDlDOZBFEfaHIO3EWXgyZ6xW8qjVmMvWfaLcqOYNw6s6byfxoioX1bBCruHd
8IumcXweLIK4o4Z8H0v09ao5QSB0AbAehxb9hGfOMBkq+eJHnrt3UlP6e0TJ/CPg
kS4G1m1uaANZ9Btj8jppeSDSG3L/8Vf1XE2B/GB2m6sADLULqI1+Gi5Ke3p9eBWW
2FUxT4BuRow0VupeDe6/bw4Z85E/RjlvVA2LhrUuR1wOx2PViwDvCRAgq/rZHbR/
FPLAmcEDytgXya4ibvdeE3hdCL/jen0sEEj+lQVQR1i1fIIHRokkriGjGtN70t/h
ZtRN285uiwpJA4aa+zAKI/1GDOEHN8aajG77ZNVknKyBQMBMLWoJCD4BFqnWO4XP
l6dp7gqMOFYZYDyzXgU/tPjQ1CBtVCfDmi/Oa78tNA4+DGNvTTs6k9FuhkXO7tn6
q2RTP5odDcj5Q6XMX4OY5RtYgf/B3fDO8Ycff3WKY09yP8PDqp9xfrD3B1cRJGHk
/IcRyCnHpm2/e8710xESCqQNz5aFCfoLd7QleEHQBhb8flpva92N8C9slKO7+hqj
ikk3zhEeywKHc/awLyOzovTMDk8wApFa6n4s7kMILsW1VBZwNZWPYsa2AyMVe332
pwDeiotrlI95gOVD6wiNEA232G00T8YtPXEjh77NuJ1O3lnXnjav3Rx4A+yMiKrL
R8uWXWyWYFrFp/XmpXUQGH/Vk5Jw+HFP9iFHanIPdKcJ3olL8Q3EwzpDAx+c3Grc
Bi3lqjHrIAUA41p3YbTD/Xudx5obdD0KGGTdxWJ3COh5CuNqnLQbeM6SP5+1XI/S
d4il3T3a+8KkRoQtoLzdLPeMt0jUoX2qQuyUuCKAneU+Yz0qXClromCS/o+QIv+2
z3IzvfYZ1wc4ueAITUhXo+ylMY3/6NwMDTtKidJ1XWCk/2FKgcFuhT477/pW+qMb
+fOWBs3p6+bqifO73tfOWFsGQkvKuh6UJ6cRK3Ila5Djfg/kh5WRut4WhC/qecxz
bcnhlm2C19IcYYkQpHWSCaEqJ+RtqSEw/Blr5RH6mjCVEumVwhvHkOuf1bnslPsX
qei3Wlsx4OJG+p+uW6vjSEdqWWeUw0lu7MPZi/PxAn8zPiaI3Uukv+FRF1c6YvlC
F4w//Zsuif8Vg9wY7Ca42Bm0d+t/Zmjn1V/L7/tQD4fUAvAy063DEoGuo7FyI2/N
wAUnl2BmNQNgifR6UhVIriAqrHDoqAYmI2ywrHXBtKUQCXwxLallEKSpuixgeacB
qcFP2MW+VgBSbr8uI1zHL/GnE0TKARk3PFJohLoOVLSNkZINNdAIZq3fGl04QHZx
4cthiLjWwu7c9NK4o7bUF0xQxvVJBLzLNIkCsfMvTv3l94/XSTE/C1HbAzKuMfzQ
Z/vxE5K2fEJvQTjdzeUNaGvrr8wJQmVIgs9XEV6iEZFI14J98++aQmezZvTCFQGU
EO5sX85lcUtbJkXS3gVu+s0gJHnw2XoVyMbP2qwhfFOSB3fxnu/FXG7/MxeCvrr+
HtfdzKidTg44bBKcQgvPVNZe1ur8lYfeXYs1LpfobIW4MGnO/gNQBYanPez5tJa9
AWDWSCm6uKqMnVk75qGFxTSJTjMJYTewYdsF7J8s8O4kssziG51D9NQb2V7uF7QP
nwJhQwK9aJguxZWoxoPQ/J6Zh0n8+Wc5f2PscUJCoGy+eOYb/tPcM1J7Hhg1BLY5
GGgMqz2BXHmxgaAUk6oB6ajfG+3aMq9x5LnJqIyKc/3FPAW7+Ln2Vfhcx9TcpqaV
Ir4TkbNLQFypyhfahxpbOe3BMNkqQnwIXMeeEvam6kpg5QB2/NcfadNZwiE8c8pe
W+6xFaAh5Cj2JfnDaMgk9t1W5vQzedgATmRjf0/6TEbXX1G4OCVtiltLJev/R3Y+
4Evs7zXJHZYWVPgVsd4IYIbIiz3af3G7rUbNDFJEJ9sM/cscKLq9WhIvGPeV79gQ
9bBKCxpVxAMOiImlGJpV9YkNJbs4r1qSC5jX4BQDoAUBzPWKuoRRXqw3YWW0bFum
TXe2q13O7AKs+JQkgPFNlLaq511Q4G1gWFLWHJ79xGIaLIoz2L3sojsHU+sT/Mqr
FoCKiLdZvr6GcWVDVQ7wq2IOUhe+arj0TNeL9rSznhsBG0nZMQQhvTOy1YFMwS+c
F2Ew82EVZTVRiLHMQTsPlsrpyB2sTKH8cS0PoD8P7WHT0HyiwpKpI8ihgOjh9Phb
fdjY56ycfqxED8BaoUySKuuSNt0GgLCfkBUYEkAqKG607VVcVMjNCsE9T1OUhO2Z
fTFx6ITKUVtpKPh0fueXF/bT39o+p6jYD6VSli+JzDwu0f59ltXUVMUHLvz7NUGN
P1qfrUT5akfI7DTMnoYQNqZl2z0wblxVLqAUeQTzzs2JUKYOvsM0rqw5TyLfgjZc
IQTbCxC+DxS3GU73TseQJTwFak/XvHEzYsrhgkX4KsCmowXcUAf0trGpdkGExu69
7mRO48bwmAcxjgrxSZZp76++45Rm0tyyiEhuL8m89QtZOQNT4Eyp5wkc7JMpLfxu
lywHZhBUYFFFZ5dDEVTZUHAixeVjVCr4GJHGf9arAMuUAzKGYACmnHrsl+EIoJrf
NxF31oQs3FBUdxctqopj4yeocgR2EAvixXY5OJXywSEtBGP8sQXa83cCix7dfNvD
LKOMHKHi5vTgYafJmCP0BU70LXOV24XcAYKw4Nane0komr3DjNeOJtU0+TXCBKSe
te4MkaSdLGryYXZyYUAP1/wnN6lBz0mLJKCY22QNc2nlrks+r69BhTco5m+FPIMR
j3vmD6BnR8U1RZAa6HY5AMGP7E8AHspi1Y6qc+L0F4w2TM+ZsYmgoNsu2/N8119h
2W9hgzv1RlLCK7iBJ6huCR/h1oJBsR6oBQETMOrtTHD2i2MaqrRVJfA8LkHQ6J65
ZTrNzn3dRViMo5UIrcN8joXk03slBWjxnHaN1HZIh5HOdHeD6Ozohd8hLV8o43k2
Rx+mI2Qw5RvUkTY56OTYlfEph6zBLKf0++kkyOWbenD+j2gafffuhn9jCKwpbsGO
kdgNAzc0WsQUgqh5lZ5aakXFfO7tRgTS0LZ3e8U5APDvilH/HBQumv9tFOL6ZfIR
wOU2JL74uEwnWTaRih7oUNpWDEQpwBIJvdRfyBhk2R/856PyMYm3NL36Yn98y2Fl
RD3NOYB1EpN5GRgbRuzGmFwR1VEIu68mhozi/CTIOIQ1BFBl9cZDyB7V6W+pdVMa
ePJY89mZrLyY9IF3kUSSQb7QMplzNBA1ddTWXsDUD84N6Diu8XmucyfluAzeHSyq
qB+LUA4QHieGCUl+8QbfjKZnTAYNX1MA6lhDXRLyxMsR7xaLCM/j/9bD3nmn2AcD
Wt3/n9NWETnK0nXIWZwMBHEODUowCh97aBc5ksO6vwkwqlrHsxObTq6KSLyjCOAU
yGThRQZt4Gk+zOKmh9Ea1qlfFXdCFwwnVBJ57jTp4xHrgqiQQSYdSm7NqGkh2Wh9
8U7A/XGqla/0rcempMls1CJGkGda9nRgFM3RFKSS+Dp2AXRfdKKZJH8wpYN2pJXp
JPTgf7AY5Q4DKNmKNPsZzukicnxyem/AIUOf/dfPfIfQqp3vrj8M59bvL447+5Ni
imSAjJzGXYUCu354Z/92lFKmKn7H/OQbFD1dztA665KjpaotFFuc28q3FDUJuE/r
qyZcvtnMMhShrtmxNxZfvCGplA3I0y8irGbhuUIEZl3Hs0vb3dDghKkgEngAmhws
v/F3NwYiBf4V0ZfU3ebxfl+8DriwbCgPSdZ88LFKqUUiITL0OsiR0oz3kdrXzMdt
e9YaJXhu2oEOQhLfQdtMz6pu3rMRrBE2WUSPYq3/IaqQNFERwMvlS9lMWNgTnuak
hA47irFfsybOkm1a4hDNjI/YerhGlauR2RMhx2UMiLDhthtOoF7Id567uoCYNDZ+
u1RdI4a4gCQVodqgDVQJ6qKYrKNURQHsYcr384mGxukTvtSa8YPaQLm7F10AWJMh
WxAiVN+R2M/iDSRKPyYUelXsuTsBRSds3Ra4nnnk3yY8tWvsfzjGm+qrXUhLR1Q7
l3H/7hWccmXF3JRKioJbHKF+GmxQCdEp5bmbtuAAU1gTm3+SFUCOpWbLHvbx0l1n
mRA6RAH+B70+sv8fA64oZmP0p44Iv4tfwVC9G1qkttpzNyN32/jUOHpbppQTvymS
MwbV+hn04ktfjrbojbgGiQIyj+PinJGxlphtAmEfYe9tJXLcwBCDlTSRP34uSXy7
i17cw3vqk+zJmG08AlETBM+YH8g/jxUwqRHMAwfrVdjQFcCahr+kYAr6ZmGwZxQr
+fR1xqekNp3VijbN8x3u5DbtLUA80unsMTzQhRRdw/huRK7Go1yvUeKqknbHC0mz
8z5JA84nWgrIgrGEsMAodr4sMI2RETRX+jKgFtfhs5697k0NhFPsIlU+qq6rePrm
sZhHnHDhu3AwBjM5AfQja4dZkTbqfoJaEfT93iHejjbRgvSUj4AjV9dbgQ1B+lii
o9+Q6S7zMkxOsUBPWA2Rnfj4svyQzbR2kVK/ZHQ+B772vuVkfI+iqqayUctQahHe
Yw+u+8GnlKxn6KXOjMb17CHHwjZZN2kOaKQs3DUiM0NT+Yw9XHGeGvTmRVxI8LN2
FJbG++otQuzyxb3+t4SSZuf+TViEqPRcUtDiZZR5k/rfFGgl9/lGiQ9f/rt6fZDG
7EPFTIJVPCcnbzNdEpPCrq4w/epvu06LuSzAutDaP86CjAFy2c5KiQUWNUgAqWzY
UVf3RKuQY/9ftLhoIZir9L2Z6cUzjKKEoVAIeZkIfjTdc59ikHNwocx0J0KaRqom
+7p+LccgYq+w337x93dAuEzJwD0EnKRrU7solcjKM3/wXzoa/S7q75wAUeauxfQA
rAShSnZor06skKhVv/oKamg6KAeWVDGBSNyU70/VJTrRbE3nBtCC74AzYXMehr23
CT65Qvud+u8Vgc3X/Ae+dLLwGgvMwoL1gm9g+tbO4WLd7c5Dx5+QftZdjBKoq4ZA
NMENcMbtE/PuUfqV3P8HoJT+U8/FwS9q9x+v1EKaVo1+OYqIYTMSnBGbud1wwqWe
Rpbyoc2OLXJkxLRrCWRKvBSNfrinM7arbI5Fp4+RhMYmUw2g046k+sybzUtwEBj9
8DpHUgreNv5hbd12EJogz48VaVNs4I33V0pcKPg0jthK8a/mR/nGI3tt+4ievF8c
cZsObGssf7YTRCJcyv6+Zz+XLr4AXQ8iZHF9Me8+0G4Q09edSf9aeC1LIBAJwiZs
KbsQwHf8mzmQoMiqdAGmrclRV6T0sYcEmHmx/sKvjLPqRJjuI0GKXh05yyGjnf2z
xp6KywfndlpoFnWwoSkDF2ucKDr6h2Yk19ENZRzFiOH+7RqXEltRpirt0BETlVhs
enYXDVX1M2eBS0LTnC3MyxJxo4+cZWQOdDFYBJBMd/6iy/N5znkyZj5Bq3b4pjur
pBjFV76Rei3UJsdO5Ohe3HSt+OUbfrl5m/vB0NMJOKADfJ5zZo02X+ivB4eukam1
ogesZJ9lY5SPD4eiKy1irfXwizHnP0bW73bANubrsRI+gZ/wQw78pgxp2HXzRVzK
Zt0/Uzfg4ky0TQCM+1K6qbqzOEbGOMZMExkeexPUsCuRR/Xq6EUU1O8ROYpzEXt0
j5FjMr94BqfDWgvbmPF2VahtL4PySZhziczHnQc+oxbyFAsS2tpybB3LN/kAaIhv
yXqEBLPLpLLoTdhEqf+5ZBrzvT5XqD5wEcBcF/gPGkscpdAFwoG+hVN6yll1W/1O
a9zWQLutSEjc2NQ210ydX0QKEU+N/b98pwrmwcfzvbMPrGceX58Y8GymQ8RUdpIo
GoYy/uhPKX4qWF24RDmdlrRZD3Z3GITer/Kue5v3OcANiP7K5/Jb0eS9c1mXPqBi
1z9/SrP22fmVlEwmUCDDviFmCv+UVzBaB+WrUw/FMAdePYEuCG53gjHp9atX7+1y
WMPSGo08oatcHK5eDksifgp7zv0CYOw+26mHoatC3ljXZiWABX0YA9oq6n2YDJ99
MbiysHISoDhCQ8Z1qDf3O82ogImHNaQYmC5pmv8NoLxQT6U3DT1ePVGtg8xfhTL5
G02L7UoGMkHRjXZKybfGQc7SPZYOb6/GV+OTGKT6Xg8xGGraRaQNo+MWyFaYcE/y
fFSGBKymDDWb6obvZ7BDF5tKJz4571y03PQDeVbn4roKKrJqFTxgQHxkkBQMcls2
IPXgZpSY/YouxVW/gwNdL2DgM4+iL6KyoRboDFbixQeLAyyiFJ6hOtG3Q/8Tjz+Z
3YY+9zqgS1MYkEEVHvzffTgCMy9Qc1mAEY1v/2jfJqqlEN4ZksHdxHfe/kvIj+KW
DvktwFxo4P7VQklljcFPAqxyLsFkcT3T0Kwl2PsnHwLUsV9AJqgN3Fr+rP2W0vwC
4Tzg68OtmGwX71s78cwom+3oC6++nHTd2YfTL3ovOlmyjduwMHR3DVm1J5M/+opg
UiRJb/4X9V8Znkk2588/jFs90f0vjPRTJqWqxIK+ewRhXDPIA9SZaJ708DVRGoJ2
tE44KKP/0J21IwqpkaT6SVOW/2SQryDwL3GoPTrv/SSBdXUFMK3H1c23ezYzqSJM
DeZLuE4tRIpPpUbfB7D0evJEGKLIfuBTC7eXbIJii2xCekASGAN2mryMeaXPF6wG
qxIwrTqiiHdrkGCOEPWDszVLqA+q4T/ya9zc6nY71k63mJ0RuCxhqwehPLc4H/ro
eFNUmP4cSL61zzVwTYbPlHi2fQp71364WzrD/PU257jddpgs42xDfSuUCM33I6pu
nCCP7k9gumZBl+uErjPEjvE5aBoOXZBTpPbdrA6np5qdx57IiX+U8FvRd5xoihiq
kmIwpziSq4TLM8eUwNpeMMBbvKUXNLND6WEyOBLef6SudacRlGel4/kWVRvC785I
jI7BzGAKcWz1WzxrG21vHUfIkbg0bSI5CeVuAVZfG65iCOmUQkPx3MwNR9VOmtr8
GGufOAes8a1VlWIvm6j2Lir86RYk9dSgMUhWOglqn11QImU4qelbNUdcYwm/5NGl
jEjWp2vgLDR1MnGNrpCKSiE953jXutzMk8IRiMCdI6E24MAuMNx033PHMHIM4Z1k
sot68e5mbdugo/yAexHvs3eVo4xBTrw/O5ND6RDNC1DQ+BGtEIHFfSGGG86ECw6w
U9R5pfTBfVWg7qJhvKoX8j/64EHXQE4N1a0WKVNAnc3F7QO3YCmDRZd8f5lTH2wH
UBxqyz1/TN5Bk/Yp28xmbqQ9En235TwQFaL2h1lD1gDVYIJsCenckA1D8+mgxEv7
6E/7PIKytdFOVq7z0STA+DFtRHoSrGjg0FjB5ni/QxaPfP6fHIQ5D3F+DM8j0XWD
2PPtjk6nk8MuzaoJ2MVLfEHcCtHg+GVyIKQwOKvxW8uv8WF7wr34mS1MJsR+HKkU
mX2XiJyg/pxCNm/N2ifH+ngvdA4fZNU/KpghBuPguU9Dkcy1KMClYmAUflezDJAb
+bGfC52Iz5y7u/66gh6PHLEF4wRe9v2vdr7yaMkYfUYHjHdXh33NoqoSku1PsdSU
dUI91RJK8h/5KS/WeugIRFu3+H0NZUTx7aiGZbvjv92IDZ8BfB5EElS/sa+owvfb
ezwTkV6ejUNXi/amxtsoSDzQEawkTiIAscJEUpIuv1L9A09QeJ6XsZyFDCIH271H
2SozbbvMjieXZLoj1kMdPAwXvrirY9E1TNEzCniRenxAhhHFea86aS3tWtNYng1C
P/0TtnJL0Tyg/PhTFBh7x4NGal9xtNZIFz9jc4aeQNuaLuBlaCz4LNcDgmceZ6uQ
TQxrzp27NA+Y4X/Z2ql515PZUg2PluxQK5PGmUkTXyo+1HU+tl38fvOaCJ4/CMOb
DnvOZFtWAKa62vPvmf1SyOih+JnKin7Cw8SGBYVa0oq/M9qxA/v/fn7KA2UtqOsD
YFLwY/N7IHMWvxO3g4XfJKHymlS1M1cBwl/+NPlglyIC8zCDSojdHcnCYItMinbW
jW6S+f95ltl+9g7U6esEFu/xr7PisDB4DUoZTlIlgB90wR5c5/TG0jtGVOQWlkqV
jJUrvSzltymnG+ivsf4nQxZoTZee4Tw/WlZVxcShUKCwnYO/flnC+HjD+ZyQcOOD
+OPClSpnzXpDKWR8V1fDR+C9ZKgg0FmParF8xS2L9OfMLVqL0oyJkmoTsAEpRqX4
5ekeJBHMyBURBXBpXhTTAkdmnXURhY6R2k3y9CfC+/nYjdoAXeaaslEBIvgVsod0
dK0M4+FVubfw5Hfs7El6X9qRbA0J/yXE3Wc6+oUsW0M8iuqTZIJ+FB5HMotcxU9A
pHBDAITv/aPzkircDPFMv4pPYAHUbyUqCSlRn0hL2pP85R/SvfrpCUk3Wxj8kmqB
v+ixZNDzanbsXAzNr1O6GczAlBT0/f3FP4FMt/n4CUQ7/gMlkaNfFsuCT50DSZt5
yyyZXxsbf52wQ2dIO8Z2G9lwxh2LRomvpxiupChjvRckigceswNgtMvdB8F9tL1T
x9Vlphj156qMmpiyWJe7BWqNeWqDpAbmoB/a25r7LcELJGtpWK8gDMLy830mCWh3
ET5HowVksDxnVgqVF6HhsvFT0qr8B4SSPUKlZYwdIJuScBXpvBEozmzvOsIbV1DJ
WJ99ZNfUFNK6ac4Seb5vtblrlKWLX3lKV0cJpsW8J0itOQuusvniNbFFpkFtBCSH
gdXaI7yNauyXLkLvYMkzKhheXqRaC8/ypWpKP01l4bkCTmCrVc4r8MSqlOzdjlHo
Gb7MN29c53BqfjOLoc+cwy8yq5P/mhPD4n9I97RUWiUazEe7MRHzavzIDaI84PGV
UXvVW+B+WueM1js5fnvUlvU0wILKreSpNuEYyiUH/JgqYlaH+QefKzts8cmvsygU
OAJSWpLxYYIDslQc7gfMJU57B2KaNbpmu/x2ILoCVFoLwdpmvf/Z062b+SkzNIR5
pYgWh2kzWiVTjmbqb9+CWeopo8yj0kBq+G5mQUe07K0NunXLxj8h/U3MUo0ecHdQ
bhTqn30GRpUD05iR8zAqFIQfm9p80JLQzpAiCehnt3ve4pUycTAFkxw7Y4bCt/w9
dD8DwEvHXwtkH9n2ymNaAmMvHRqGbZzBhxapEqaWQnWiil8+a++FLSHlnPMKo8HS
/6B5Ryb+lwqdpuMTQEoxtPqghEhk3mIiuDXT6CJVHhlwYkcdp2wlVcWul4+A4pmR
tyLoPQcNRbM5m9t+dAwaFc+ZxfZf9A+Tasn+8M7NQRz0FYG3pHcavToJN1NXnkY/
dYcFdm2agqehHEi0iHBVzMs5IUcihfYubNfFxGtxkzEtMwkCB5WXo7SZIcAv+JFa
oWn9f/Qn8YhcoIO2jArrYfYrD6AjX0TAsW5JlXvrF6tMIVEmJHdN9fpPIxUUb31h
qayShwGqKsHlTAoZUp/JrHoCkd5csnqvuExF9Ae07Un6MGA3t/cNQ2qsKRTealUW
pE1Oadqq7F/YuSiPqVyDyY99prIeTWZOHHzgICXAWe6NZ/h570XVvVrvzpYo/4lD
QPUVD1J5CNM4k7D2aJnPaRLckkGoO/gaRjf4flK+pEDvx/vYmMMXLn5ZvdoH4C6C
QPCr0HlOgs64WS/g4c5KL9yb9P00/+OTG9nCguDNhDDL+Wk4bHeDjXdLN0MlX/du
jGEFNby9wR+/IM6l8v8Ltc/waCIxEltKpWNA40u1DD4X6m7DwtWlxS8cn5ML8+AB
aRcBENTvs6UGsaZuBE+CKWpquOXnrtR5f+nSh8oNFBzyE1WMfXCYCJJOxs4yaHnN
15pNd1GUd1sKt3N2W1MAeQDDLrU+b9ifJcRiEOwQBrf24K4KxwxjwWmDKKK+yUsx
yuYgnGBsqAD7VFzVhjhpw+f9ZQraPlFIV8KBln5InmsO7kglA1GpcFENzmZj8+W7
7c6JF/2om9NyN+Nd1Q6Obq5sTonKGZlTCGkd1py7/WVW7sU3QxJ/v9DPHXv2rgHk
0N14oKT1x1IX/BZNi5wTkTQ3BKAb61eyNv18B8g6CTzdspoRtI/JMQdDoJwTLkXD
NMGv380n9DuR7C0+iSLzRyyfEC419l18mpi6nN8LJb6dM1s2aZPy7++gnv0k0rHt
Otw3H70Xekr/ij4qo2ZtHldcE5iP64jeZsaWsqYSA3dgrZnrlyaf1AMduzCLck1s
aJ+Vlbn72nKzqoo2QxpP+FGPd4vZsh9NGHvBGYe0arxyRUt7YnVjSj2YZeSjxJMD
qbUZXkCAPg3rxNLuNeH2JsvcNzK9p7BmVRAn2L3MELFa9zgppzPT7fjpuBIHQCxi
iOJ6N9KqaoXKFWHyLunzpDGSHVvpULYfqW3tEWx/BW2lAzHAl2luoYGLjEcD+amd
YpbUunnlCNCwUKmW+Vvz01oaQvGep2SWfdSEuyHceh7QJ+LuUKEWnNp4C35mEx6n
n0bi48yRhjojw9Aw3nb9aFgKK0qKTee2ouTpWlxdXtRalE4OcVXog9F8D8N5wxr5
wfODOp60bY2o1uog/0uG9AtKXG1djKtDtbsvYvRvN3tk+NPP0JqOEwKTWrmnXs0p
AAnma04wptCBb4keXCNLyv316bomlvBnILL8aTCiuZic3tSUI73gTazldaC8jODL
56fdFeNdgCThjVU7rdaAXwIqZwpCPHAl2atyFCeH8rPmqVEuqnMAwv5cKffRbMTu
dmBQQGRbcuYj3h6A0FmOIhVFgp7lfGH72iy0zv1ZytJkwHc/db1viHr+nO79+RyW
/JPkroa54XDPiNBvkSr2W790dDxxDNbxzp8PSzsx6aiUqcis/2bp09QUg0zJkBNS
X07cu8ndoxVrNntm4WMvLkEjKqt+NnhG9NSEKQkNd8ZPDwi/ltuYQAznV6kE0p3I
YXWdyur383bmACgq1uZ2N/xKpExdSTHnuBkwdciF7A+rmeRhlyvGqf0IH4epLb0q
q1FcWQzdGp4eaSWFyLxGjDCe+oeoBfpicGjb1vJNriQfqscZy5P03+y0Qs3Wd+L3
Rpo60BL654AOhaoqA21WKt0w+qoVxLt/J4KFw9FUGq5zzWjoKwmObT+NfSR89wfU
kU79qDY4iyrBTFazoGQC0Pmh6KDDjomsbKYwA5i1oiPxF30cWMOLBa/8Ka4EpWmO
qmfhbKQZ0a9XuRKgT+Vu4aOByZdOzfMRS3fiCiY1nVotDZ+JdsQ+E2sAQH06xwaN
c9uA7HDqw9wiqddOdcL+Rby/XSl0YvWQ0RHIjCRX0ML9J8ppi76vMhH3uFcUg3Ag
Ok5ZeLHjdVf3j7oIhzqL9R2hmxfjpOzMwmq6tnaQ/dbHZNQBDEAZR1dOW2MRPhtz
zDN5LzbbGm0hxbeFHgzKsS5uTKzrjKKnLO5c9Tud9291a07vFGQewsVJ6YUQC+YZ
5ZrlQ9uwZbJSbK8u1lKaLVJtSwpUttnsN9VgrLaRFlDkPHcqfsk0BOlTPVe+Zg36
V5F5aAyR/LJ1F6yeE4gbbuVji0ftbWN9Hz4DU3nB6AolRyaSaAftm9lyDK0pH8PX
HnrndVoPBFm/jX7jCcK28zVi8h7h3AywMVL23r3GlSDMUpAo6TtopBjnDb1AExLi
4fijoAK22PPM6Hqj331UdWPxfv9tUoz3HTc8ER79hXoM1Qoprt6ZclfypMrYPAr/
fAyqVhuJilnLlmbWvhii8oatYoa2IGs84hRDhAfH3D1udj+BoEQD07Zhc+hXf7Jh
mPxzYTw3quuGM+cTd9cSjy27i9Llt1mDxcg6225FOT1bu6adNraT7jVSGauJVGC8
0ClN9O2txldmPzoNXiZC0ExHjMIriVKpLCOwBwhT8l8pNNiDdEGyc2cIh3zWygiX
A9Ci2nQ6QQL7DSZ4ijdVmO3Lmv0s6LvQwKfZ4sucX/tykBM1DfNiRHGsEphqJW7l
sukuHrxnSGkLYzoIXc+x3ikBABav8nnyObbBkf9b7zFo9DUs2oKxl9fuT+gLSrn8
yTIYHZj2nzggRVr9Ml+21+/qSO3lGDiD6pSfsXzFkeaYudySAi57kJQaA61yEp5B
BLyK+G9s1dkBYpv7Im4kg5WLQ5wwSkKuS+2PwzfxQgeBg2otpUfILiFKxB9WiLQD
alNhNuzMHKrgv5bgI3BUPxDEagK+uKBUfuEfT9+0FRW06P6pzdfi/WOW1culqlNh
O6jljN2NriMLyYxch+2/mmpqZehNMFfLg+A5AzpGJDjRoThVm+UjeEiIxTEJrLVm
lSPamva2z1GOy5tffGdcj6ObQC8ETWHbPnrL9jSxPbQF2XSGBY+nCE5bEuAJkuzC
CuNOtuMu/a+zLsKKzemdYKUPuMpPvYiiDux+BRlp5JM=
`pragma protect end_protected
