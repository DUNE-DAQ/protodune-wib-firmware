// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JGIgYa3Dg6qS4D5DI6cazFlrfJ58M8EDsBMau0SEZiANAobudxuowuZKjB3LoQ3v
aFoVsmOlaoal08pwEUc7TgO624phUkG98i1BLMf9t1Q/G87mjDNyRlwfvXZQUfQ9
6OsL2iJ36uUeaxOS17n1nK9cwe/PJoLFm/GZ7AWZfFE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
f7qOjwQpgjLaYmz4u9qczxfqlzN+d8dsvDyWUvLfDTttoYGfs0+7WzN8GL8iIM27
Shyf16r66TRFb4vSxgvdkDqo1p1ZL77vHxdekrH2KfkkdBgkTerh5KkQahFgLAh9
GmFxtNtWRTfuU+KGpqgEYYnEbkko6DUU3n3ZPRKed2gifkNba6T/RX4PHQapIO0V
V89xuXvlVg5mUq4qe2ZSqeGqCUcPFKWEp8W3Qb5gSqXCh0Av6IkFbvE53EJDArqh
Ra6ddo/fBz5bac7Wgq0cvXzaY4Jbbi8pJIFfmjMYP7+vaTwHrnbr2PSjgUwQYwyL
iYIvvVTQdIG8LNBoetIaGdzt7lS8laJhxEktGYXfLZ9b8ey3IH88MfaB/9K3hZp+
ZkKnStV02NB37916kfb2A2HREfxIPC8bouJ0dNXLruwb9wpv2DwiSrMCsXp2Benc
PBSRIBSbVLBCInergHGw2Tyvwb3nQnGLdQ6X4GAGvH3TLiQJp1LtEXKFvRpZQG9A
2zVhK002yz4XRP+Ql96tX+pJ65ID2AKJQRruFxgHrRmgyMnLbHwNkYNgtfV/9iMu
0tAhQ5YLEmzYL5sXfRuW2jH+y/hUqAE9qj8qWUgqYb9JIMJ0nv7inhWocwvJgT9N
+HTiF7uG4r5VwE3y0SNiG/uBg/3E5C9/YJBOB6VibL87MasUwIXhZHI0I+kDPvZ6
Aqy9/C0tvMH8OC7n0zqK06NhMDB6Ew64c9pjS5LqODr+DQjwj0ZKGuQm/iGch9tf
GRX9zKS6oswXZOODpfIzHdORkxK7EU34EhOvLnjsecIl0UxIdhbs0cnGoxOFwnDS
UWG0r8hSQ00MV5R+CdASJFdwXx35cgkwyQngMhkYLqWNUHxZT15grb0/v5hXvksE
+caVjRiTOHU7laWEFFNT9swPNu4lzoh1KslkYW7pSkmNlHNZADmU0lwCOXMZaNM3
HjM2LknO7uMkD3u5BRXpe0yFrtI38B2agCAOB/TV9FtGbqYGatilxUvAv/zZIvvj
DwmRxFn7hDrRQR6y5DKmCRsY78McAI5XGEKpnzFsAteQ/TyDxArQAD2qDEy8/SX1
xOQSsY5wLRfO4ken+nh5JM0mVlKIDGs0L37mhunDVqP7Uh9VTSx40GlROYOD4cqO
thj8IsnbC82rbfTOwbqVuR9a7j1crD8kwVdl80d2u5VtH4aw0FqMgk34ejK9/BP2
zvnGaVvlUOoqpV656omgGqLEdZRA5MpGl6jHN0k9qaxLI0rdwkwjqyI6ehkHeuB0
I3ES26ouuLO4EgEu19igxHl+o09Ua6cJFtC3gVqkf2vBd/C8g2qmFrRUA4ETsw7j
iHdi9nGzZB0rv0hc7ucz4VI7a97ZHrqUl4OcrlTfslb35jiX/YjUeqw2esDW8vbP
GMMxHqY0JFp/DSZylW+P/uu0cs4qSjYbX6h+IugL5st8xLTAYj8v2eaUMoCx66U1
WyXX4XeWYuADA4XgOTocS2l0RPoWVesUyqC9l8LUtlCWC48v01t1StYJZe8Vj5Nc
tB1BRhHDzdQdEMUscHcwSFT/DFi4HbGpRjaNFsJ2ovpxAR/s+VDvurb7Sno7sWar
HRDfQDQgAPUGFOWiCh5b5ZaIO9mkJZB4lNRAUh3FNjNgTe2Bar765+mtiSu1Lu72
T3fzsOoLF1OBip5Fmwb02G8jsSFroRsVr+K9+rME1AhPcVwPudtLSH6P+hidGx59
6Wo6I2Jt8Ty+7LRhC85MKpz8swkw+8mm/CsF0pHaHj5B4uQWElQ1Z0+2oAE3/mGW
xYfZk4geFcUTbE1psPgeA2ckRjErXGLVWQe+28h4tBJS5u96PxxPdqkKf0MBBRlS
a0lgt9K5HPRJL0Mswd0WGEhNFxigdKpOEFoXTYsueq8Z9/sGRVymM5Iui4gC5BfE
m9H6l4BUHLaWnHEUmKJKVR9SA1y7hlXdK1pvlf7fh0OM1l0Uj5xmZYWBGX00OH4/
XAaxTBRhVj9mN2kYLdmmPTGb2Znlh/hbajZeEA0XK+POjm180Jwe6lTvgGZjdp+J
swePMsBNl/jSrwOztwQpW78iEQJnZKfn9a41hgHLT5ZQwF8ZR7x/wqSq2n26PEjs
/3wnOKwq+2/iA66xNT9vIxeTAcAm3EQItAYSxiEMs+/3g9+gyKV10vXl4hxd8MOl
O47nfiRE0HX53Lyd2hn6NGML1FVvLkMhwNQJe39l1rQ/DESSDXg+ywtecWk/nUhc
LETHIe7kIMDyHkrYjILcHkJmWQWnTi2wyauRZoIwL4mE3soYAy85dC+71D1AAbtp
PB8KsgGHkvMcXvAaUctyVxqtV2rkTz/ZCHOi8ztL+TWEol0RNrHF0C+u+NwYwEeY
7dIHQHq9SYZZEpVqv6aexCFPN/DX/oMza2xRiC1zALVXGiW9nfIfCnKnCCLVMngl
6gkZhyvrdXnYTSCyJvRh6fhEqel1xPvDyK0DrusMdW0RguAfglUncyiezOppoeF5
8PTk3Bz2a+HBVyDLt2trF4z6w1tdnff9iNiQaTeoibSEpKU/eEtILtiIbl9Dncx1
pwlMYMx9joMzsWDSXBBIISntTzolxtTGKWNkq8e/bE1O+dYCxbnnEVxlRPWIJ1C7
uHiyufH1+7vGuhsVBhcAWVmGbwVmf7gX33SuVf1AaVfSf8i+hlc73ti0O3SR5wM9
MSwRLI8w1CCR21gJYHJvrxan3PtAyUqj+ugSYNa0981kMFnTD9DA664Uc372cYld
C0yFPDt6cgMnDQA+zaU4qe/c8u8XkeJbKI5DMlgWdwsc6wWfrLxpbwi6JlRAw18V
WkDCz8/795SAhd1CK730/mAergXWwFucxUUT2QcQc26pIyx5fcj88CX7pZ0A+/NY
ml4VUIh8pZTTInKDnCIY0s8hqGYIKUer2Rrp/W7M2MyFKpAh+uqCJoTHDqH7zeLB
ng2bfB9pjSxEB7fM71YDTV+hfkw6rxxgPiEXDos2q6WDBjffAVD2erRD9kh4h9lN
OQos4yByGvPnQu22LAjycUbYnRtXCcOdRIcn3zuV4ab/2L1zJo0FjttcqVdHkJhA
auxwOOiogVZoMlsoBChu+ZDlkHjp06WzcuEiya4OrLVXgWi+7Yp+L+lOM9T167sT
t+WC9mqPFeW+juU1ITVs7dRI1JTQzeD2mGWhdYGPk8QZsIKXy6zXjQjKrDm5CNEE
aa+3ekeMcnZwr3/Hx3sRzdNV0xyMsIqPjrSY1tukwpTosYg+un75B47gifmXEpmn
rxYhTp3SPIwUmT2AOOhSQECgN7v+ELdE0ZzR/2Ccj0JqrlYIelC6xjqaFPSFRypz
zAcY04okvRjP8F/snoLYXQ9QmYI7v5jXsRmCm1qco9vIbd+ofoipKoX5hklZJwN7
H2F0B3FOVTwpBuJigeyKqbKnEyfZ0YLVphShKe2vXbY6nP7FRSBfEdgXayhu/iEt
+n1MhrT2bkm3zZAs8iK6ze+r/4Rk4ZNIfrrgcc2F5ROwVi3aBwD8iLIBo/oM2uNC
UOAaXeri04DOpQ5f6DKvoI/vyMx68/NTT1OhX4ina0jku2kGCBm/VvblOo7kij6x
bjAFWCLVNgoLRAKmemj89SUVbIDkb282kAeiah3SQDNlWzU2A6im6BEqEkDd/fiS
GTBoGKEkqeBDlSK5aEXhC7wlgTifgiV4bB0E8kMTmUuYJncrDNYtUmZ5rNstjR4+
HYkR+BE678uzzcywXZlrHo6nUm81ZRgwTC5vJIm0ZhN1Z+qvC7IuUWOQ4PSLF43G
Fp1YKwIvqjFKS10gl9520TNmaHfLXx6E6RX8kkDRp8G1VjQg3Ut5PSyB+a5KifFA
7e4of3EGcChJldUZkrSjoZNnV2RUmQvbkT8y3eWiqgCmzBY2IoLhzBS3gS/3J+JX
JI57W9XxEQ2I1LeiYyQ4io51k5FcP7MvqWtQkFn6AZh3/plFwnJmoumxK2rTMJ1H
RHwv8PZ9tkBm1qEeiW3YRPYz5OCWRpLCifwY3d3izi8ORPM9Y1payqbEGnakWwys
i23eHwpuCWQJq3e9JGxZmYPsu0VJ2BbAuKJWcejSrXt5Txv7RHh3uYMRmaxgwPRa
yqgbXs1hQWirtNoVzDIH3yb3H5Ms39lwR96cT5CQjv2ZQ98dT38EJglL9vnq0WRJ
BfZwRt56LVOjS/F/Ip8HfF7oOBPUGwcNFcyYQ8rYGCKbcG5XbWiVbxQX61oEOrd0
EP8XpcxUSJPBmiKk5R3hOsoO26aVURPqsaCb4/mihhSY6Tq520wlB5KAEum5Otst
X8MmZeByc0xvnBJHo4XC2JHWQprtztmzsONasssDsxBy+yH/zPHl4tc3BNENyBiK
tgIhNpnf/iTP9e9uOtIk8iOcV07CtQNGs5lHRrHyCiWNA8cJRKWT4y21/XvMIMwP
3Z4ifHMo+zB6IxtLTwT+/rOuWBebM6hi10UCgeMQ+AkgvAH+YL1IAWidhJ1eDwVj
xFPdECc5274JDLgdzZ/i+bmbeooPasULUmxg6qdkCZ7sy0JwX55EmK3BZXxZ2Kog
elhnLUV8NI1NuylS1o3xDChWD1omOznL3T7rfx2cbInu81oLkOb+D5NQ+0OD9M9q
1vzn4ITkptF5Tfe0jHST8cgoCZgaSEDcvJqvxqMOvhJG30QfUiImZ38dYr68PGuV
6lOyEYzkLnhW1YbCd9Xa8FOcRKN5sFRNNyU45JpgS1TCwKx8uIwUOiw7zJsxkiyj
qrNhFH8C/ckXcbxJnsN5M2aR31ioriA2BM3mbAt0zBBGNEJuOU1HvNic9xAnUm5J
0dRw2hzJDDbECdJjH6uI1l8M8fzRXGMrwyP3G0Q8jXh2QyaGYGn78WPKskFXvu87
ohDPpBgVZTECxkEdeNgRPg2BaSeHmkj+pV3rEtMyi31kWBceCf8wXVNhDp6j8PUq
P5Z6++U6Xd4ETniJt4HI69DGvJhHOQYRbNilKO94meNI/QgY/Pl0ApaOhny4CJtX
wPq4aLktD4z0RZDggSQK8aoaMnaNmLh9dPUEJYst1DIp4x4P4o7BFvetQ7irv+hr
+ykz0KsV+sXv+OXLHe+umLsXsj36uN77uFUjIeyO0lWCmdLZhdWNTCjC9oLFw7MA
VRh3XKzO8AU+Cyh2Z9wsTZXvQpnEEyaZLSNkPwOXb1ddime+poUCX1PLoJfFL4B3
5spYVd2MxkLmPEuAG61MoVuNAqM7+eJ3meZlTRmSEeqqtH/VDRCsjFmg7NMtf/Xn
Bv2Uu2IcrFgAm7nFD09Tmv6+wVn3Qq45WA0vRXbEJviKUb1tIssY1JV+fRfwWq2z
ZhIsVgszTLsBMrkUmwvWLMMsD0tu+xQQWUsQ1sQnJTTNMIJESVeVJPAtBKgGeY5u
aswEMWUCiP7KiNgW/M1Cej9wA7I8cqm7bprHX2aPvAO4OADobUfLXcc+x1i0JI0r
zFWa+k4saBC8i3LMjz8VcvO5PnP2ZLiQLcgYJ/IulHzcf0MmCyTozbiZ4kz4io00
eS5P1r3cuwALzn8Y8Vo2QMJcA6x/ckMuoZR6yKnktkQpNoKqTPqvbQV/ejwIdHv/
tVpT9GXjJl9nTrwcwXbmAT4yeWmGP2E+JuHMCAfcaSUgzhcceizfuBCEXQEdO7r/
5cXE0PmZ6SsNadj+jwC8VekSv9f5vIKo+sC4E2QQ3LlzrsfR5QSzTKtU+5+O+F+S
A/OvtQxucl941p+2a24jCXSgi8P2Lt0cCm3LYFXetwSb3k0wndkZDB1/qC1px+5M
eh+AlBAI3GZePqwrWxspFjLu5/i5k1NqTlEU9gNsWxEdPsbKbE0u1aMugykqqfu9
zUceeNSd1p08LxaXl44gWRtpPKKNTPFJbYu24HcBMov1PLF0xHuQwkoZtQg9feHM
qkGyE1PE8Du/KWjbIU7pXWk/ZLtV5pghdZY1kolwYWKkbkaRZLafDo1ywaKEGuvE
GB887rvMZmhFToC6FTsIL8p/g/65QXjGfLSlOct6AfMV8s2wCN7NgDA55JuluBbj
Wywiq4fHM9751E2QWKl3JwOc18YDf8gGjcoKlba/Y8iRqglqCH1JqiFtLCNY1oFP
0lxcIPYeTzRV2hN7usIID8wX7pYAxb35zVE196FEhTIMPVilyRacWXegoSesx/+O
7sjWFTlO6A3O8IrUCKi2DUsUmnaI5WDplcgjC7yzJhUK9/0zJXXRLSrrjpPDhUMA
MwUvFmcrZR7aSGNHYSY91LgmUB6fi9hcmFGiG8wIM0Zm2zvODzEeHbOdFNj96yJu
K5ERvodGmaxenh6ecJK6eh68+Pmc6nk8Lq+oUj6rA8h6vre9zzAnio5dXuQC+c+Y
bF21ijvLxb/+J2jy3jaRfsU7yACGbJ12gwzyAy6nX1E/0SESsNi8OBLCRC3qLGxX
qVaIWXYYDMnwxm7apnkWyox3rrT7OVj8rk4cc58OQ7UAQSU63XxLDNqL0i32hcF1
a3z0URokRN759wTg9UIVTRena0tu+uN/EQWu6oFpmIFbgwtTyFJ26K135Qpwx2dW
7ASjOOHInl7wRp3+hcqRt0XMCRpThFp7orRY810UFx5ssoB0dsfcwd69iibVOjXX
W0trvCssUE0iQn99V8SzmiqYjqNeHqfrbfZnvat4jAZwxtRybsBZG4gbAzr0poK5
b4ZSI2yovq78v6EjvWYSrF3LpGmhzETPbXyeNMTy13gj6agrnvkYb+SGTrd1u31y
nFZF4i5ESslH+qoDkuxozM8haQc8vv68wMWqAFERlinFnSbW3CyDpM0eV7JfnNp3
rHsI3Sy2/hO5DlXlPv3z/vofy+YP7O+T6kH/fmxBQTQ/MC6A1PecmCXwnolHennt
zMy/GCazFzB9l4KOfZMCjwxyR7J0nUnMyr2c1yaz4fM0MAIsAj6ocW3/yE//PkSK
2/W/zb1Liw7dB2JJe6Bx3Be8PlQkRqg+sDp6u3fmz17RBph2UOrcp0u8Bco8Tz8h
QvLzsphFClbn7ndISa4bQ/+L0K+0+ogI0gKevUqr0QGqQMoLC/RiLcahCFEVN7jD
Xgezo4r0z1qYDloac3EdHldzfvGObdOlxymGMTmaF8PFSdyhMEJZCx0o71Ag+IOF
M1OD+f8YmTXuk+xM/65UtzM7mfpVzXjwbwwiyjl2yKt1yFxnPUCsMiZebrrFnNwl
BJCK67jYw85PvV2PDnjK5XmusiOXLozP1wnFyHOBr46BQi5bUzrOUe7jorL8Hnmm
XJfTRk7e/88UzMdqqKxggRjWjtdnBzvtkMYUz2AbAOfj9cfdlQMVHHX5AyHOQXlt
4lN3uN9IFP6qOsYi2gKl/WmWZwyF2z1Pd+zqXVaGNo3sSpA0JOQRbAYBK+ThcKNX
J7xlC1SEkzxG4anR5CoKZjaMJmRV66L01NCDM4fu1grbvi9N6eVo7Pffw7/Fw0cZ
F3Sy7nZ2at10pTI4tKq5VKF/2yFVH1bW9emK7Z4tsRXBbFyqmFBmVtTTqBKbgUwZ
NWoXqmO7O4iViaCUWtVouQ==
`pragma protect end_protected
