// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
t9vH3GanC8NSmXa8BSCPaqcXqPG0t8JUpzT4kV0h79LW9VI6yXQJn26Xx7VlkK38
J1pzpujohDeheJuG//C3keSNFkennJ4h5N01uwuKHGx+bY7anmyamHsJAEfrMvi8
1+107mC7sd5hAKjCkwWWN2iVpEyfKwNv2bs7tlEpawc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70000)
2yFvho4oJNBbXW5DiSl0u405njsxG8mmG2himERp/fIm/RKZ1k20U5ELuJDbUZMy
BQJ7PD08w/u5zUt/USsgvSY1gT9jy8rEQqOSmqrjOLHPnpDiZ0ileQ2KgGJgApmu
a6aNEAjpKqViemQeFU3MNe7/ce8L53h3ftDPrN9zYuZJo24q0U7HaIdiGKc7/k4B
XvMdaYBHc9Fatw9VIjdDFYGwtdzUxyMYoqswDBbp7NR0WVW9t5noTn2LnQBgPKQ1
hK1MY9K6jnyQBDkZGa0iOmvkakpbq2ERIc8RBNTZeQDJa5CXTtkaOcvjS5BQsJ9m
K7DrDcgVX8sTtBlRT5ytFSNuYgfBrO0TyxG4PXwNGzgROHAYv2WhJvqhDVhPgxHY
bw9B+EjM5AIOlyccvroErqdkQSOAH9WiLETxFEP+58yTN8FXIDJuMLUtdEP2DaS3
DCaloD52JvUSp6smB9KO8g3UgJv7OHBDJVvrSRc8mSWhRlX1hzcNkcsTmI9U27ai
h/6KS/C7s/ZL/a7fIc+s6biDh4oFzbMAY6yGfXIbosMSMpPSlyVg1QmOtVsK26hb
vpqYfGH2cWtm7CEpogXQZpkRn+1VamrhJipWADA6re28/sBIc/gR0Y2qQFWJUiVk
FehnzaFE6PKiybUO6rHgbgs0EJl4wvp2PSQmZh5QbUdNgMWqWsJ7Iqcr/hjU09iM
rR48tN7XhGu/LrKHQq6tteOFf8raCZYnCwB6RatjJ4ouYXNByShHkTXsPykEijZU
x/ZTrikI+vQSbO6i0VokxIQm+M8cYOVFrOi9W7YBFIQWebibdQS1g2tro5PkK72v
g9vALrzyD+poBIwkehUvyFbDnwGnfhTxHIewuHLb3zCz2GIBpPpWKyM1HHs5ppBi
hPhhCC7Dlo+CE/jdHfVhLhcgcZtw98pMmmfRjt8urbFqI6CY4z1VtlzQPjesJE+f
6RxmQWPjp1Bc1waXFFyZgajPT/xLBy8E/Se94fHH2gSEwGC6xGKJNv6FVR6oizTA
jqGHpWujz6iqwDZxL3aukaGgYeLVFR9PlmUwQzDP2xpJsTYoGW9hr4Zlur8vo8uC
SJFZQolMP+GiiQ0AKd6oACXQPvN8jmgS0U64q20syj/PGM69L8JmUZWlFU46QFXm
Ja4rOzMFw3XV0tQAjAHQjyQkcmhGZLZC1Y6fCnev7nj0kW+ZJ82NSwM8xJqpBMul
2uCL/2m2MXEcPqlbvJFODk9AbUatWjHmpk/U1aelhoa8Sj0z6PoLog3TYKkYiQyl
OlhwlX+Ka3ie0a2133vnmCvclU8T8M4hWWM0oQejNAWghVlCYzZ91juDGgMOEbcG
Q37gefs0s0cGc88zNldng2SQICBjGIZm6R71nMpUZZD/dCg2LHG6ddkcsfYTwNHR
qMMDgZQM10H2QYurp1wMtDuDishRoWoMV/Uz70lu5H+swErNHdvl/CwQerY3JWM8
xKydUvjAoT6Rr3hd5/O0wGwq2RjcoyDiZhjdi7FIQky8idXrjJYAyd/PNthPO7Pr
k4iSa8QBt2JuP+FLHmf/u1E9eSZpbNo4ZrAWAUQRiLYfsMkNlZzo9rzNLdvqvfus
dKwu0KJfFfcy4P/ClvZeTzhVWESnh+dh9I5xK2oqJLEENhzjyJZNkhW/xmInvw/J
8gmifQP8ArQsuRrEUvQuo5cQX05AFzd8ZyPXUoayvtf9iGffrRCQh46rqIFY1QkR
sgtOL5Wa+AXrUORQi4HDnd53gOC2xrhYn2reT1K85sO1y0IpJrmDle47ZQ4LBb0C
4GFBSb0TO3lFWLnUkLJXZ08a77gOwO045ANyNMj6NU9ZHWfpFOxsDkyrjgw7GNbW
CX5bded+eps2nAjCAgAViE8mUwm3CpR0yGRxlLHz2iAupIR/6MuA5lSZFlS9Kxro
RkAOm61cs3xfdHXYORLwPkHr8NhT0KdapD+OpQaiVkaWjB256/rsgqm+p+ahVnYg
Snn/RUKbgOFXpS2uLSGw8oFfvpUcZQxcXmoj0tHWwaDoRmXi2Jlk6tyzr+2uX17c
NIFz8UaoQTxH4atzAdbaVt9G6zjVNBdufbvU2j/KVfIDoRlxVoKBRNB7yLN080oD
hVyqpzlfIx+b28yK5F2WksG6yQrReP+UEGlyyDKFNX462TADHIVAd6Enw10sILdz
NDoqLgP6S/33hQ5ag6E/2b/ZUtqeqAF2jGUh2TrM/9h+0JAumQF9lGann+iKwQmn
EwypAfTG/4b2VD1aq7LK/6PMDMG/cuIYoi1rXspcdWEuuHBxVaCwo26l43znO8uc
3IWeuQapyLCRAHjNW9b5ZODUHAtTI32UjtLlGsRIBRecsjD78C4cdsBa0zmYgNnP
7P1Ivcm643lJoHkiNCGf9kcEqerj8zdcFiY5+7cWfxZHWZsJSTBZLPg6Xp/XUngN
k69maZlw8y+2ESehbC+2N4yXW4+xy7iVqveP361+FUYmmiaYLOK3YrdXVCsuRkVb
/PGdSgcUb5MKRV8zWwYGlj8zlyrfi9N4sPneJnvcPW/pEsmnaJGruz9khKX8k1+t
WseSa5CcKZYlfBT6s9K/iIxpp8gFVNo8fenqKvVM7DUFXRExUQwJMiOVSYZNEqHK
1USvgHZ84zo1vdW8sKyAqC8Ra2dBXiaa/jHm9gKLqWNkfpjEgzPc6RN64kq3JwxK
TMU3H+Ss+G5bAGMNKE1b2IXRvB1IA+jYeI4Cgap1mYvsRfFkQTIFCxnjbNSjocLP
WUxISEQkqIl8SkiSNAH2GdB5bGuXfwyZx7j7i20mww1x/FLdJGHUwRYolf8tHpA+
Ls1hxh/Q+GlL98YZhhHwiNHA7EGoQyq2W5FD+WXsJHrX2CgjuncDRA4sAchK7eM9
RXKF79hO3yxVq5CssqUvZz3wEQvOhkbjKXSo9tc9g58M33fjC6jdhacGhLkH7QxJ
hslh8tqz6eyB+HR9WL074gWpJIWFmT2+7DCtxF4WWpR03Tr+2zjusOUDTX/nDQA1
ELqeXVT4Fg3cyTOn51+FUGlNHP5iIM12ghTy0VcnW1mnXpdr4y+bO6Vs0XVhqzTb
GWtFkgCv5rt/qt1JEq3Jjgr1UaaGDi15+LpT+uyxHFDWgJourwBLuDNiK8CDs+nT
seT+gxOpPBWkzSLWSUbWxAgZuVJVh8vmhGG+AJERurvqxHwxLZASVI0dH+JHcmSG
5H5ENNfncZTbD2gQoHWxAZzHib3rBkKqe8gnHCzap7INGhsi8JmW8a6xrBW7hBL9
Ip+xd1yD4XD643yPAG5KXn69pivmxAnAFCFbyFJaHTXFnOWF8xvEKT/FEtUwNvgH
KHfvB4rRrZcwVrC47J8oXQ3SaO/r3R7L5uQkm9KBQA8+dzAR0Ze1lScdW0Kx7Nk6
dz6fAS9YVEcMAYzJ7izitg3xMm4JDjOlkZ4Ixk5xLCgHmI4H7QAASfkghznHAR7A
bt5CyN077SM/96OKYW62cbSatR0t0K61bgDFKKAvU6gCIiSo31yKIqLxyV2wKkcO
yKTA/yv1Efzx3ON9lgbaY8TfH/Xr/uBohT2p7NrjQBPs24YOWViWxHb6OuEAt5dE
mhq+LcxgORpsGeNH7969g/uTF6x51ARERsbYY9u1CSfwpcJnyxVeJ/3bRKFWt/sE
eEj23wVxRxNJ8vp07SxtoednObS6ZzVCfqAmGd4pIoSFDywKWJ8WHj7xYuLR57s9
mbjfwkAHimfgSOcw9l3aGM1FALSxvOVljCvnOcT3TJlMKYgiLKLizENpf+64bwHu
BIsdJKcrQmP+D1Kvn2ygUqW7CWsb665KTygaRpSEy5it8S6+jXLFVgVw+E3LmAC8
I3igeFRnQTqnqOKVBkOLrB5hcT2G7sJkmGzb1RORojEBliNhOoTFQUhQYugxkHmE
8KpnXt9ye9ed0IGtNkOgw4n9NQSM5Oig8hFP3l/zVjaLZ4sXRfV+s+b573tkSZki
k0xTUH0McLgB1pkej87cT5BPqfdMzCMvgEyePWLQTccaU4v/HuWFHwuMgQM8rKb+
nKhVZNcWh2QDlfi2o3MBTDP6hMS65P5/u9ikDhTX+DO2ovfm0IDyd0s112YKPCVM
mHyYr0upQkdYOG5V5sTMHbdeCBUPKnNXJokwoWq18qO2d/y1y+Oq/BxgB4Q8qo6M
0FL+GlKhaDWfpNoHQcV/g8f5pBlbkO1F5FTasRKxGEzfaf3nWp8KReewlJykx772
kmtElteZIKSWm+D08kuENA8haEnOB/y/ZxHGLqMY/kP5MAHEe/RzREfgJGpd9ZF6
wtkTlphzThNdz4tuCO1BmETa3O02ar2QzBWSXGDXSXUaBHoFqFVs0LilLC+6CAAB
GwrkhBzOm3PXX77iQli7E2GU+Est0nHrBQ6mgxQwy6bPHGzym66dBELL4i9dG24f
5T5VIHJmEbTMqY+NZ3Hw95DrokSiWJ3STdVFHXjl1aTylh8kE1iiUCuW1BgJmYJD
eMMb+3HBEH3S12t17WkWCzfUawY4LvgBW9rCj48aDyn2EKZc5tOK2/z2SW46e43l
SPKyPRZpRn0jR79+PwabWuvWBkqbz1ErvUOVkCfL9SbkCHv2Xun0EtXVlQ8NjLCV
gWl6AlaaBV2GVIE5+V20M1TPZzG0OsosD360K+tw7MB8fLSbsse5fBumM4j6UWfe
ITxD8fUWlVz6SQzzsT+Wuj2TfFYOJXFwneC387m6iPUEq/VW/48l0n+y4VDtYl4M
6llH5aNeGHdp1rFvSP+ayQqfmhLvmiBW+lpzUxksQ03UOd1iAB2egKEUo6yaUO0H
l59tBZl/Ky+gHh2xQoKSBdreeJvcy5t+J4PF91wuBeSJlfmyJ2eMoGb5cWnhrEzB
hwjq5JUca3baatPIb3SRUNCU0xkVUH/2NzNOUR0GWiVP9gAOi9N7VWjwCV82BGuo
kAcaAijc62hfb+UuqZxiSNQt+hTfxLKOtcA/Ko8VoalmTnycmdiV/YHvVVfF2brP
CwGpnQBMxm6QyQ5JiJv2yhlrahw1mIZwJIPf/vFzs7qFWaqMqaL07d4fUVxcWVoT
3qRHWYUjwui1ep+iFvIjtaJVgHeA6bBB/8MLWz59olXDGO3gcrttaar4FQfEJG8e
j6ogxiVIZ7INZwuZqlkMLgOq68xvveO1/eyKC2LWeffFwzKlWhijwRLHOmanp/9I
dng/+64uFX37PLugaMmVRbBy9B1aoEeMQBDD0qU9qsA7myyRyn6qGR0zY5kgweVw
1+N0MaxMx+ojUy5L8ipOqn1yFsSSGq6wN+T8YHr6ABvrDQsmlVKkBallE8WrXfSm
Vjw6bYDNy4j9cMES68kLihDHCoAGAaLBlCHvwoHcjFfgfmSpiJDlcyoGUXvYuvSA
i0pao+erubbGNwkK7IGWJydAZYIlR4cczkHoO5zwkNV07G9ue+VPvQazMGQAMZtW
pFKlhTeaYhUZP3DuzXhaC9x/KYMtbmVIKE6qkdFoV+QzPu1cLebx43Apbv4XkERD
1C8/FPptYOj/qS+OJmwfu+no7zKe1n0dtGUR0bQbC7/o0TRdhcTVG0Z0iNN6WSYZ
UwfqnS7Y7/kS8bs5ec98CDTEe1fT8k1vzGOfhWVLchCM6ZW5b8OelYQtFZ4JpC/e
6z/lwQ8KzkwxCHTk7bMN2KwPZKmsUyJYs8lJRLlwUZ7sglQJZnDKIrQz2JN2SM6x
NzyeidO84o8X44yqgkbECz9qQ3iNSWUSLhvaRGhHAY49PjC1xeAXyIX4P4tJ8rvh
7vTufaBFv6aWwGSTXZPfiiHSO0dYBHBFzb6Qpe2iUkdo2hTLsCjZz4PyfIljrvoD
coPpSFXrA9yWkKgqAy8QLXfYk7znPlZp5fbVASFuE1tmAO20kWdjN+47Tm/BtRpX
D/qWVCRZwsrTBJ0GNJ/ts/If6nMnuNvr1fTfsdpVmcoNOPlzUYcNS4G8Ey2sXDBD
g0MUrrhyQ6wS9wH/KCPXmwUKKo2dv8VRQumXK04k+me98CX8aJmAlMcCSwIELIok
aTH/zRIzOXZzYVT1T7YkZZPlrhcp1xR+K6q4ok1PL63+V83sa2KSPUJIZ1jekheA
aKzQZf++Tiuw3gML6YaBWAqeIJGfB5NdQ/x7xioMkBvyMiv395t+2oDV5fwcXR6H
qmLT+XZDEv6RnZKemY6Fj7KSoRGa5OszwgfoJoWI+lmn2zh3Du1S1pPLClLNpSfr
jABy5xuPIPsWL0YwV7NjAfdKBDUUSk2WSuyL0qk18IQamz+dP6hmw+jo7SzvNiLA
ifqN1E6LbmRCp9WWUqmYLGsDLY8B6CEBsHDAbrNfZImERhuo2RUmpFWtPAS8xt1I
KMz98kehPOqwtmM1r6gGUHE0nl50ffICJHuHUzV5TRW57toaG5JnyzzCj/zX69mN
6gBdIPLtk1m39vSRMokH753HRehwm2gVRkPbDUXP+mdVSYtrWtm3HUvgJMaCN4R0
xbYlI7M/92xXPKQSxbh9oJND2WBHaBOABzrj8qfoSlXzmp5hYGQuMmQch6NLWVZV
4glf4CiFpR96Nzssi4z/g6+vXcJGSLPSZXILOaxRCbqVm0hqHuRcZXTBp/ZHjtku
aTdGrRlND18Vzo1n8f+mOg0Y6n0Yqr6WVDDAVW/BZvcKzeS9JS8wUQPUI2NcMAtl
wJLc+FECHy0t+xnD+UegQK0oHtcn5MGn7FxacWvyIWd0r83/9XhgGUl06gnjABRa
DH0kaTcPGb3fk33JEOed1GF8PhYDToClm7SJOkiM0UhcDmKATKykG41o0E60+qL9
9o/RqxRERfj6sPCTaDUpfUSixpvH6S0Eeq2ZZzPzKLi1z4pdDw25kqz9Ny+ax42E
7HT79391JsFACJGMq3YBwaFv+IYYqC0Lr8nQqkghzINDqj3v3VPUWD6okx/MhN+P
0a9f8owH00alWn04x/YFKgplVL+SCnhamToOculXZqBgwwZcr/L4fB227pcODVC4
H5aIY9Vu9+9V8ocbNDnbr19haUdKzP/bQ7/qlO+zraq5DULYd+nKD8748/IImmVT
5px+Kf4GHoh0DPFdckB2kxx/LtqTmpl2eLr/sKKBsJZCshqkVaNJh1S2qy4aNSxG
Q0pmoDWeUce8LIglMH9TAt5EkZIwTdDaFKg5sHbN8KAkn+tLA1sdhIJXulFVjly9
uRFsqNCsfJOG62sOnjscNvEsumySOjYP0S1vplu3vFKMSlhpQQpSbVpD7XXsHqGj
ttGfuOV6jBtcBE3xGVhsbNM/kz1qJ+8SnkxxMKZPzun4JZRcsk5b9h0HA1X3oNLi
Z7f9fC/yeSIjDeo1fX3ybNbHslmCtG7fdqwNb0v+nhXasiX2b7viIBRHaDL+ZmzQ
F2gI88wAYjbL+1LBg8YG8ejAAQXPF6/z4GKzGoMb/DG49EfRlHwvFxwznuigBVym
ddCOimOnVmVq8p8MMc6pDTQ+agylgOcnSqJ+Ms7fjiBRVjmtYYHAgj6jZqBVKYtQ
NsBC4kopN24UDab4GvFeeN1fuzIuWE8SsK1Dg7qnHn5qUe1J8Ec0NHriiBb6JySQ
X2EkNAm3+XQN/PXgkVNERScWAX+6+64vf1eQeWs45RfwIUobrKvmANgSowceGg1A
7uAWj5Pg+nLP1O6uMZby8f7NnzV9eUPUfICj+7AcOm9KvkybPnDYMo9aOEFuMsPy
cmgBB5GPRiT25FLs24cR4bszd49Z1sNH4oFU0ao5qj/yYQYHJVGLsv0EaN9KBdhU
CsFdaKlp+ktZPhyS3AxYa69TzxWPMh3bW8dfsxoM0VdT9VhGg3+AASOpy2R5WSX9
QJoJNK/skVSzytKK0XC+rGBGy/q09Q+NLh/u1S0lu/e1GWI8wiXKM04hYUzri0ob
k+VX98czmP8dMA1I58eRIhUzApL59IpaoWzgZvA+4VN5d+B0UPEsQurAQFo9Smvj
RK5BuWd9Sw1LrGL96I/BvQRmA+zcbh9/NCMqL+VnxveNWGuGOmMpjD68J4M6dF9n
ZxMc03Z3hXOAiW0FRm0j+oA8dT+iaQ3Gfqa4DLAE6DeyBrqyS0OKXxYZvxQ3IU+t
pud+0/nLgowUYMn0rffh9RX/FSovjEv22KYqckYNEU+SXzjNMJuun/yCWkLprmjT
TP69wbAaNfkBgEy+9EB7rgvaZNsYB+mXw1NXqpWMgb3JeeNlv6ZMCRBiXcEA+Jfl
rmZU5pnGoptSiinhldQzuwQB1M9I8D1LzjqvJyM/u/sZoetSVPWaqPoQXWKknY97
TmSpqAUetl2A/Hzz32P4+JTT/Acl1qlHC4/K7CwGpIBe5s5YF0/b5cw9lEROHP0d
jaFQvJU9qJfjYjkxvpxWXPGpgv8C5so2JCp6GOnTFbLlkmCXjEbmTf4NEUJlRda5
esNl8sv1QPAX6CAQAlbaVc5YZuUwFPiG9K5qBzGEb5U8FFhBlGtyZpFs9nbAdRxh
kirZS68TdjY0cD7K+whBp8W5YVTDjR/5bLPDhi9xQDDacihrXmy6tesFkY36QUxX
gi4i6MvuJyDQyzZ3jsXjB43O8qIiluhquH73S0+YWfpcAInd/4QmMYpmRnBtfbrq
9B1kIao4mvFJHD+eXag/pauv2jsh4edKdVPJbC9Um5Y2/lzoDzE7KF8mxchEbasr
Jt+sB7zZLwTzmQMCEoVGQ9bx/d1eMN1UxZDQGN1dYuQKKy9eR2v0+jCxZ+83f93M
OwN/MobLVQpTdDww0HdD28xx/v6lvIVJ0vUEfsbUp5Y2YBIkgLkbeN7oQrwsdkHJ
M0Gjl2P5i9t16aCboESfqmptPu+gbIUE3Oeq1yGR9O8WIEpBb5qaXmSz7SnNcf6D
1M9QCIaYnCoLTVxUvlwnXm6GTx6KFGIcWed7vscOmjKHBhY/5SjcBbZEOk8umrbX
tK2FoQMUDBbxRuHM+ZkXGcVJHCoeeK/N/W9oqEMjqeTre4uiw/iYxoZV+9WX53Q6
j3aJrQEXBsKkvtvcICyb5AwpRooJx0S/w4v3c2OHRH9opyf4iKz/dbJxftYcIAlK
q2i6QHYwclBpzOXH7RzXpxHoTo1GTu3Yti1lCG0xZPur3IPgFs32eQqomSZzXaIu
il3UWkZP9BqyJqsFYlBu/jUSKnsAjM1leaVI5BRF6G/nrZpFEpus2UcEVygJQ1vY
LTclFDTL/JWLC3kRQFyimwz2IM4LuArD4zhQdAGbKtyfBFf4MhEDAL571yRvwUBB
jM2SB/VuRfKGzYPy2mFOrQv9P40Rm6t8Pwe7dkaFhA6gRgJqUZc6BXsZ0HqhOLHX
StiSc16ejgVSOlie7oStmZ5Ilnp+mTyK9VqY6wY7IIWJlvnwVMWbpnXkXvn/keMC
x0SbkMlIlvg7Hj0tumpE2BNEKjNv/icnCCeCUZWkhJuSTFi+Lj6bZxZu0U63oLi6
kQm2u75OKI6iQPRdR4d7XKN2eaA0FoGXnO8rhgYuB51G9LMEhBWF59EYOmI4Pook
sscjUEPSXdbYZlLt0dYO1XnI1gQ0R4mcFa+GUfP+bpv9dmKKxsfdKOiCsNEHilz8
HbbOPSqIzwAY56516K9x2A1Hy+ICbP7ao60DcofJgqs/w5UMZgqLUBfrdA0TN6ER
9HJaTfPTTiOBBGRLgHnWrQFdPWmZX6Z1/O769w+mpIKpB+jt+Cfi7pQrMYu7NaU8
sYXUyBo8MsUrVQ+5xfo+hmeNAvZ3evAcDmaPBD4QKTmNzYkFYIqzgrwbiDg1ozha
CL28rBt7x4MIfx2Of4JjZovAZ0AnN3W0FJay4E33fDWoPkj8m4cGlidn0b2xpvGw
Ip6D91xehFalI8dKjYAJk6sGETUMc7irEqm3dTgUwT0q28GQIoJY8DK/nFXQV5N0
t80/JrTPqjE9OxgdnqYcc8RHg5Kfe2FXvwIItjZ1hf/HUtogTRC7UjBuZYdfrFjf
b7xJYsBqKBdytXdDCqNBoZ68z3zrfo16yjokWbTvMvGLR97nNhP/kjDrFc0ANBgR
BUe/vXmP2sNOEr1D35Fz60k57voNE1WZffGTe315lELYviYykIeIRtYXfncIdPjg
Z42RoUZDFcGD/0qwD41pdYSkxa3KEflWxl9Voro/JJi+wCkP/VAFySjN5Fqf9UJj
/sBdbQ2Ny1Lh6WTzA6QigiNUy5X5JOXbmpjSCnKkKcmb2dNAXZduH42O+egSYsUC
r568R18hb4I3LUQ/L0FQO9lyvBCzVNhIyEg7TceVZpH/ZXFHF7PTveZFDdrqaj64
Q5X7k9BbHVRfrJIkUVp0Kh0lsYqE8aUVndCKIdE1kBBzLc8ZXvF+HdRhNoPlQJPw
ZSHwVo92SQnItVjDurtTjj2Kik+pYYCZ36jg5lpmpC6VM0dKkbuImSw34I6UZ09q
0iWY8q3bXnj23qd5/f5fRqtmRZS89SxEPaIUxhOxdaNTeNLvTRhZjCbTNBr1Oq85
lBl/mcH2lj/zZXOqdnh3iAzuxW6Fq/j8VH4XQ255N3421854B4vP4DzU23DvhS4i
5zs0UaQsE68VykvJ2AGu9BdZ9QCPeWcvTMnoL4blLhEtUadm9nQXIsiLtkxYFMIG
fF7gd0ckMPSlu1zXqzKicnpPyCJP+Ti1vgHaG16x70ECQDNPKitf21ZVaNXuw9xs
3CU+e2jE3xJHDN9JkSaethtrX/27GHMqPvoHkZaK7tohABelEcO10cuKiYQKIAdp
QgyLUaaShucqWa7X9Mt/lZM2py9Pxt6zNL52UiLWc/SLvadXF/ZlcPzpZI+rTMJf
JTD+js19cuVEhMkTTZv9cJRGvVJL+k/mD5l90/N/tebvDsCHZmRdejRbkf4j8XV9
9D/YQX2c3zg0W2f7TzmkviOaOc/eZBMesJ3GwbmxHXicrYg81R8ePVer8ERS+aDS
g22m/eQXGe6kVzhuoABPB9Qb2rTO3Bnht+WAAbJd2cBFt2SyPFh0ptcX9XwQQwBM
nlEAJ37kcn7vzHraGDJxB/Lmaz/p/ui9UvrgHsf/zITIqeNT1BX51Rh7qDivXlCQ
Fr+08VmmgLmfodyaf/mVSqQID8pGIIhlONct88A6ofagmx344aML6gM4fjFrOMBc
FMdGEwKJOaMKyRm7piIAoykgfmYjiIL49PwdfLsV6Xg88iq7oG5m6pmQ7M7PIQ1l
Nb4MRd8XUyzra4J/e1V3OpLH4fFQgxpC9v1tn3SgS0pX/Oi0BxgIZPMBEy5flmJw
HfdWFy3vM9Mx3viNTx/tN5omztyvtp5TChxSzpGm8D/ZCUPGFngztiiY32lGmWzP
Er+mc7UONKfKY6+lUp98JQ/g8jR+Ta7dF9RQVqPuE0i8eU3vTJGQU1GW3rGh7OgV
EDSO8Zw/pG7klZKW96TGrIedTeQzDDuWHdAfmogqd/VoTFP5a4CPKmPGOnax0DAn
z2BOUTsLEjuar9iUcLd0buexUE/zTfyMl94lTb/zxQSkVdHMVlPpMEftFmzjlFkS
wN6bHc9dPWrJIIIV85qrVVPE5yB6GxmVK0bbXA4neshvAsVaSp6JrP3xnOQXXbal
WXeB05t2WSc+qwXn6PZGQ/3Kt16urKiEtHYr13MlaCiSheQAfGObZe+wzRn8Oa7s
TZQ8HfO1cZzcznKlrUfBAQBVZwgGWAZ3EMHhHLBm/ooeBd1ZjRm5fJBwryMF7zXG
hTvm0OCblfhToCg/Da8fv0vMKAyCs05WRtIOUYSJoD7K3zFGp49jONkR5RbdtxrT
wLP+7rsi5adel504Hg21AhNx3ovyStGjugEdmk/KxanUC+1Jm74JVrw/zX2vywGf
KpMTR7bE9Jt45s8QncWsBpElAP6E6Ft3w9tIOntUXAdtosY5IpLgESeNGkHIfASF
EuSpksQwcFbNbHLPNBEHlooQKB5VqioqaPBsHcqr6O6YwGXfw6F0dSHOektxAEP3
5r9seI+/e44CTdFuiroS2/WzbvQJUR3oanPl6/z8KhIpA7kiMzugFAzI99WUXame
ZSY4umJwZEHsg0xVEvxR+ZdwGsewH0tG2J8fkg8iOlz2IQ2FA0+VRyNsGd3fdLvL
AnkQdBJGBR2JNriLc89SuR7pm0dX+4ZAauk/J+zpfw4Jc6gIH+S75UZLoj5PoLzO
X7E4fvm8+jDlkp/+dib6/bSgYMKAJb/3XIcyQjymxiObe3AU/hUwuBNa/Gj/4jgh
4jrWN+9NjAhdDTHfINoI0dFYP5S5+Bs7/OysIHoCwcj8WjB4xIbm8mZDdaDabbB0
HIUTEOjhU/CFP1Ffllkm9aiyzr7MiPB8OUSaY2AGfSJlCLLXTc9c9f2qSk0yMYMn
lCEv2MQC54gEK95sKzOsdB2+GrH/w5ZkyseO/f/VpVlUAlwsL0Ktr3FU4+zNQSNo
R7MDAXB+hMkV0ABAAPUsgRJuUja1Zu0LeDbZVsSQHpoc2IG3NEaQ2nXghvmNl5lN
VKEZY4RYWKI7t7o/XqoC4gdyugtDdY+e2uE3yOzo5GuUTT2xLx5xQ63eqE+A9eP7
aNewTXYPqo5rLVWO7Q/XSih9Y4HpD/bUgZHtV+9xwD8eBvLCxVoE1i6NVO+UjHwD
oapMck4xx3gFPEfBNDiuMslBi04f+++sr08M+ue8kwuF5oLTdl9Nz5V98FSiYisk
5cPqLUhCpfoflXfDTaDOfgbrfj2py7hjFF3E9h+OO9k7Nuf1Fok1L9HAn+WKz/qr
AwSlhUmrDxE3GGPSHf+CMuw0SEMsUQT/lyIMi3yymIvFSl39/Dn/85PKP+sMPDP/
hXT/xaec45nukJ3ddfB9vx5Iqiny6qQ9N5Ah7zbRXz057JFXBrBvctf2agi+Nynd
XiQ0p7PODB022oK4lKmTeCaB8ID/mvRPLnI3nN/X0HylX6R/BUSOHQyU5BhTtudl
yAeXBo2AG+IKUdGhCzCQQP7qXy4B/g8k4lwTmot4T/Ugh3r/f5nQAqSir1Ak5gxF
8ye0xqfpFJdq5pXyUwITdTlaX9TMs1eFO2qNo3et3wDGSmDpxLthomH1qgAZwhlM
e4lHxtNeF8OeRd/BQ3Z/UWr1J0XdEreZYI5xJ1KadeXhJmtAatFLX+MsrNSaAcKn
NUnC/hCIRr3KAF1H7p+v/8oHCApB4oZAZtRwf4nRbZu0ceyCM51BVuIxXLOCOGWg
X5MeOYEBRCJvP4id7+qhFRwsW5wJKefIoN2Jwq9tBi8N5egxUj42rLcHWDBoPPGz
5cpMzyE3iAbGoOd1UVTVrm8dXFMWnW1Aoora0uXq93/uioIYWr7L8ldQ2gkk1bnp
vDr5vOIftFcZwW2gz19vFlxF9WF2hesQTYtE93E858oU+o71BmrNtETSnrKIziJo
Tb3vw/pgXkDbAk/2AfR+gnOOt/FOmTFpikNFhTa1D17RBTD5UHIZjMmlK5D9+Uva
+VJtZSVmPWycm0SLUHeAU0aDY/QIABIVtVjJzeLW18cj8e4dr48tKLf2RIEMZr81
H32Z0IwiZyhde6Mc+igYyvrYEb5awhHnKLt8jQygwzrnlyYMpo6ycqc+spwHS61I
IpjrIqhyyDCAlW1lfU6/FizJT+HIUkBfXCDQdth+tms2105eU6frJP2lP1rS0cJK
g7Hrl+GgMlZyxcpSEtVoN02QlTUe/i6xAXNLXW3l1mQWAVmvkCS9r/WoP7pYertF
D6fM3JyWW/NySTFayzjXE7CcZ6ootD8AgSkGZxq5Q0AVc+zQ2/r1DmPuEblDvSQD
aQiIT/KjBDx8a7udQQAk2TTYBV05XkdFwf34cTCLqvM2VIsjieNmEfDv/22AmrE7
sZUc5B2W2WyqGmmo+nuojcdTFQp316Cw47Ntd/vFTHKgcnoI6/mapj9YHvdXSVgO
wT3OS7QyjAdaDW4DMMj98khrLP6wD+i+AG8yjyKaG9/EDlYYpJSfUpc0p7js73Lo
L5WKCyOFY7MpUO/5xaGvF6E0pdOS389wW/N1RVt4Z/bo6W7l9kSRXH2nDpTdIM8n
dkafs09Jh/qitm0XOIu0TnjQ+iBi7hOuXOzZOuWpWM4xOy5xKw67RF2rRV6OMeAL
Zj0JRZPkhzjYtW536ZIdLqhEj2fPn6cdD7efJGKqxNxkNq/I+uMRoznrzXiUJTpA
HKiaBYBHdueZ/6s0kXbPgirC4J7PntbdYYhfSbES5oIuoif+eIpZ6p+AB1d8zyhD
uluMfPScM9/ITcfVKD4d4+TS/i4y5/KSZSn5b6gonRk8UStiBdlQ1iZX0qFsMn8c
c8o0vfz42jLSWZjR23CFVm0BFmJmH2v68d9OQoKGpnRWf2Y2uMwEbkOn9YOhmnup
D3wdJmKMi5yKr6ZmTrkRJsN3ov98QFYEFjQ/ijtZFBygqzzoLoRu1nRmEH/6giYA
vgVk5NtLahCtBRJTy1ogbg56vBnDf3WrH/afBK31WKRtL61pLERwji/w7sqaltNL
cjJiYC/ovNpmmaTtLbjpnHxARhdqkarw7VmLmp7OaBsa+3wlcgqcWc/27hxH+9h/
38balGHomlC9Ze3T3S09bSpZxtXO6XiiIaZkVXHq6w1ov57yslbA24mGrB03XcMw
G+5Ucw3q3EwzAhwrbHwRmIs22sqO0qVXsJUrbTcyrxM+ZQGQ3Sj2KG0ytjqVahKg
hbn6tub6onLK7Rtdhfb1CbvHguX6syHr19n31G0ugVRHsqqu7fqsWE03JPDsZSmP
porP2MKnKfl9zWJXMEJUICxPLCn7gBLkdXbkqdqt2aFKF7C2MXbVz2Ll9VuikyxT
eU9jA6+AX6jlFlhEc9AyUZsslILD0izt3KKSOM2Raswy5Hcr4gXncTqS84fHNyAF
fHBgfpeFhrDDBv97kwLdBf7zp8tqhTtilJIIVlGJSZTEkkT6iBisvZRyIapePJbG
YAZbkQRl/thRCtJLBLHgekUbNPsX9DVtJwbtnQ940Oy5ZoCELIO6QgIoEkcBtNGK
ZPtSYArvm9RHEMJjI/rEnJoLTM28gmZjge69/dtTufYCNAQ6hp5HNOGC4d70P4ow
dzLKw/fGHXmhlTqV/IcGe0zrSorrPWqkvknIh8hBs1dqj69pRbZCAPxabuqvUmBr
Sj6ISk3190bT7ESOuC2RGF31Us1cQ7c7zD/6C1qQe6PKZA9UlKRVX1GKf4pXsvaj
Sc1H1oQ6EPaSF9F2bbBTowcCaq0JQRGRcs8/YmAMBz8pV4wHwztSfUYh0IMYTcsi
hBieNehrJENgvxmD17TnGdj16W/YbAFI9od3IrjQrti5TGvncg9QKls+zKBhbEe0
nUXru/arvocC+Dh28Qk6DuFZ1pMygk2zmybUKXl/p2wfmwj3fdDChAkV2EueLtZi
OA1pC+CAK5HFWX9Kjw1XOZFnpY53ZnT97b8nD36Y7NHyNqDLSboXFRTNhJHiKvhF
tVqhoSWrrQz7sPbVzZZiwA2HwT5qxauRdyeYvV4xzpn70ztuWwz6viGjyWtMTEMA
UGgz1XhRr9kJ1v9ae56v6V3FArmJDrUiR+ps6ODUCm98tiEpae/AG3wL46OxvD0K
XcAdN5UFX+I8WFAs6M06uEtosvmKGnZ5OAU1wNTPiyK4CWq1a6zc2JQMR50ryLau
E265yRN2pTrqlF9/N1fYq4jBVcgo6GQzpF2lFt0zVoAqxQ4x5Wr4weQ400lvVL+d
CdtggaGbCVdIeFXb/z/0u52biJJA7orsCXzODlLrRk8d7LP1zwpDotDLu2Ydzk2i
UNZZ0pXQFheT3iX57yczw7WOq1iuEKr075DQM6kk0k+floOxgOxlrARpjbGF5Iu4
8tz5nmNjo58/u/+i1wPxpEDPQqs9OxfwOQqCEGZl9t8ox1YhJwghUVeR+8WkG3w4
ImbGXcZWNfw45ywURL0O/qT3LT7IYtJ0+K91IGUJrw1dNEqbZBnGzs8lkEIZeH2d
1shdH27K8VmeLSKxfQxtsjl/4XZhLLHuOqy1jw7fK+G7FDVkl/D/8YQ63ZWWNEyu
o0pbqVSKablO/0CB64+qeLxqBrq3AdskBvYqzFlSLRenXVodpFDTWuj1ZEP4Le/H
b6t5SP5f1/xVmOG1XW8SvWiUGqvn4Liw0uG5Sw9gnq7LuzMQFPitG7R5sxCU8LAQ
fb0nAvvt40a53T5xO+ibnyufhOkvG59+DvqsKDR/4HjxKkmS38nQGeMnGJ3zum44
VbppEeohwAVeQFYLRzzJISOJBMfvR25YE9iCt2CnTmcwRbGyiBM27q0S3Ip0Zkui
WMod7t5u86zymJsErYyunjloGf7FeoKIWRFcA8j3szOwXar30fRMuCpU15lWhKf5
bYJiYoD65kwJpoql4PEvmFxY3GHmtFh9KXZV4KmNLfPflzmndQq7DsFrv7OOsVGv
bUNT8QrG2uBdyZMv+8V9QAokShLQwD8I8j4HJ53Wc9yvOK6HLClg7hfbJxKEIXHe
KXPKEWMffI6AXapjel0LOTgPGnj03cVbXUIk+78def+ctfjFmXS5rakSFZNTAj8x
DsyjTf5+wBKAi8hTrWT6pRsecd/QS/24Ldvd/c4YSYOtPCK8F7036rKj9O5Ql2au
RhIFtqgKRWY0ottloOISpR0L9z8etWzl0PowEkYJEBBh7cIIcW50snphzV1HfJJI
5k2e0Sfz/jchWygKTn3QjM2kWQmdZ/ctHOZ1w0brvRddeRYmgZWpVzrVj+ubU3qn
2XDehie/qznVsqP8xWjBKIsAMCaxvMcDXm4axQsbQXRavXcVn+OHrCapcy0Dlrv9
/0zx/UvxtwcMScSxBGSYSZU93UustHWudbmLuFgjAPAPRiyVrbqaD8oB1SlYwxnc
27iW++7stSDyDkIp3Ko73zrWt6vYahR+S39OgMJWghCHvXkIF9dE8UABp2/3IkdM
xL/omRQxj68YXLQxRz6L2hZRGj9dJZTgo0APS3g/oLJWdK8NNzK8rqR13gsP4Z4f
Lnp2SGCefrKfUdGedaZwMvCyOoN+wiAwYBZTTIogUnDk8U58ALS8ZVEA8AZJxYaU
nCNwyuRQbZiBhfeVLjPoFrqYO7dwZB4JgtdJvfdG8Z+LsZ74dbXsIMMOrTBxflpq
mEFRmJ8FKOy3XqcXn4oqSZ8zcNFejU6DjSfE4WHEz1GONSGoyoRRa2zrA9Kr6BPV
WeQmBYPn0I+QB8Z1MU0bBxzeJqznmtP1Z2rE5kxohkLNfGcfL8/ocQopzMzQ414r
8qt4NdEihqcCDk7/bem2rNRjXMWFezMP7KG9yrXgB3ACEVppLrHEEKzydMkrTBFG
9LouYhirZcTwCsfaigkAN77N74c5PonrA51u4UNgLW8bvdpAeOTSc79skb1qknIa
i2XiysONkLhn/9IJcI/zatppVkVza1hxQ+FNHFxEl9hqfvyjUaZC41fRdQxp5N47
6rWrw3FX/7L8LigXlXRWsc0A9O3N5hAOrUbXH+zqmyn3F4+4oGS41WjuziXjO5tf
TodkbIAhUqoxCZLMU/b6Az8HtTUCRtz7FRCfeAP6HA0IFGc3KIfm4jx41betf1nf
9c6UccMvDFmW19b/ADVKFbRjlevi0drUHe/MlXm7CWYshzsqgcvKQ7WBN4/B8+WY
bleiIHNYzdxakyctGUhmiKwrWsEAwhXsbBMK88vw4L764WHDxVwRtnMfCzZbStr+
pk9cSqkYNHpQMHcGupr1+Qi9Lcd+nSaJSMI5A1LuosNP88SDgoPG5CQqgaA5iTFS
w1K0lT+kqmcXiO8fwVkupZEDY5gSPdGCyjMZ5GHbEcweBPLtZSaRFLb+Z7RpOvul
Yx3DHN8UlPEzt/Yd3XaX8PlnyeJ+R5wSNiizTUH8Kz1gA6AiwxzBV9slcG7U9N9I
sX06IsF/LI5ImSoKRt4bVXAHIN5guQ0mRyaJOuVVRo1dOzwDgdZTr+HYQQa7LaIX
jFPyHbKTw7mNP3Cb/5zJJPqBlftsAl39FyaGNioKpB78LebXBT8NVj8gG34Kz3Hs
W2PJ26yrbGTkCshwHjbNE5AndMgB6f/ATVuHyQel5OBDukRcE0eLFweeGIt7nHSC
uJi2vH/k+YXW3Z0rVQ++qVIyde8ucM/eid+qPBkFRLQ8PsG2ogqjDbTbkIgfbGq2
jRLRHZyX+Mu0M+hyPZhPrkWOJNrCMGlsp1FU9Ap48LXV/s4leUQvAUq7WunflzDL
dbK74eTYIQhRHEMMzvR/61ORyNaZ4u/xsIwxGtxqNrG2FkzA/NNWK7jRzo60CFXG
cS6cRaXMoNKsRxn9tjLW7sSYglnVck1tNbGM6PzCZjzHEpD0bN5/6QwFod1q7Aei
eqhYSpopnl+U6IdQD750x52fH1mLEqLmgUd82mv2MWxQ20nsecKx3GcuxfRhNqJK
7+T6jsMIQ8kI84KD4vBnJv5iRZow55+OmIBkEYBi9SY7rrLS1LbSLqM9ricKvvv4
sRwGA4WNX9nAJzQAN6na2Vgjg3CfTCCU42gKhMWqUvaimFUxhHl2UaEBk4hUGH+Z
Y4nYxA972nZWu6+Btvjj8Ivcdm2o+pO9hO4LsN2JNMKteVi4SXZ6hZ9Ydm7HfnIs
TERdX8DQCpnB3Ciq+wc/pDvVflQ3oZzs2phaqQsoXacxQr1A60hZOcgk7B0olSYp
RsAs2mrwAIGs3Kggx6KNAnRcyVmIIv8WYZ8j5OTVhnYW29MNBJiH5v5m6lPUtgkx
Pda34lXVo+hf/Lc4GtvDSl8SDgHLgCXPC2myVJj8VbNBJFuYxW63Bcsl70VDeMW/
spABof40/6C3I9FLl1TG7NCFlt66EIixzuhtgJ2TORnH/L6e2WT+YvlL5MIYiyqT
Dmzk7NviEE02TMdJcmXLCRAOJiIO4dinJCktRvxHFQVIEV3GyfirPQbvuyKOsbDs
KbUQ3vgXOTNV5wmNHka3Pth+hrm/xsA+ZfacvsYBTKoCEWRKP0bdotVgWHf3kGTE
/ZWHasJ/Z3g6Sm4uSA9Rf7O6VhzFsxeVWeHFoxj8PpjhK+5xQlQcyk/YN/owXyTF
KdfVydCzf/MyeJM3cHh3KxDabrNm+egyT/676zTomL9tJlTu+BN88M+zUgTIlfVa
iaHUt6xoOvsPy8SJ98SFk5zb6FGeCqzbF+95y3QsQv8B2SsgU8Tiv/IfYp1ezC+3
dK/Ps7gGXzWx818FlU8ySzhOk77yYfuFBiPdwb12WmdcXfen2t9DYa3X+h8TsezB
Qj/qFMLtOJyz0YAsKM0ROo+I2zHbyLcqo2oX9b7r5xQrmdcR0CfRuflDPHPUs4u/
EPQAg0V8Mq7UAjrPr3yL8xN0e7sHy3wYMkyoSSyqpgchAIqbiSHa0XTEI148+JKK
rnHqBQBI7Qapub6QsW+q7TCqtRdswvbSvr2bNM9L7buFKYHUWkvW6qJsjeJxnuoL
1uSYrdF1Ub+WobncoVStoeB6T/WVvGmfbsDQwVIOsm+AX+UHmeYIaCVrJuuNFOwC
nvUzwJPDY5sia3CSOwTuizsZ1Q+99UPRuE+jw+73T4Qalt+H3cfN1/Cxg91I7pct
sB/va1HkVqlRLuXVETS9SdSyOOZXtyRTEpK869CFjjMaMGc/4mVYN97RSfTSwFmV
Gbkq1SVtyvQkmymAU8pndRWZZaRQus3gqruYM0BRO9va+gZSw1pthPZhvtvEvSCo
0xbKRriQCsD4jLBnJTaEjJl2Hn8gkn5nTPdQp0Q1V3hqpnzB0BRHFKCkSe8DFRBC
xCLTXjAQHvmPGYiecBfGMXIRe2a5JreKlFMJWSIXvCbIU4K9wSjMaES/5aTG8zGN
mypSxra5b3Qrwid+qkY0Wjhs7oR7KZ7I2A3m/TbN5CdcPXymI7eRmvp5+clPYHY1
Ema6D7CJF3wqn05I4R0CfRxJ/gy2qXbOsuYryJ2hmSUth/quimF3oydgsomz9twq
+nDdRYbI19k7lZC6IbWadgrEzvUr3mPsQlJVVYOGHjQB9whfwjNdiusEh6SZ98p1
tN9DULRZlOOTf8Qw+snyRO/IIUz+q95rf1dKBkLwSEEAOSj2AjjNpkq7ZPfxbEn6
Z1NTkNNInBSez05OPcYtb//14Btct4lvaT2QYS0q6f9d89lk8gJ0loe4pgATEjqB
Ma7KkWlsaAsZs7FF2/5sYdbQJtgM9Yk0UiHt5YP+RamfdyvrFV5x87afOW07Y30i
Dj4etlH8iZdLDUKhqOxThEmj3bk3Sy6PSyeylygcJpXfhXBFGoh0A7aYOUKEVlID
g0yVG9i4631zoelMJOinY6HkjAMBoD+B0RuaTl5bBmE5FHSnaQjbyfiklVxQPd6r
jEyNuQCaEYCSU71j+gRqDPyVZ5GX/RRi2lKlTphMdsO02LeakUcRJGxbcvEPWx3Q
UeetTVNvzOvt0kkBDU2BPuA247R0NVJpMbiK9KbfY3SiDqFvShuWVNac5lGKq00j
PZP7uv5VEXwurftCjhcujX60dN+siKjiqqt+9KfdwnJnfvLU90tmtSe4gKC6Dutr
YS1sEaM+76fuSYjCBElIyE/U/Wmk/9a06dEKDXiZw2248rNHW3ytehx6VT7HGruT
2Hx/PVUlDenHBtYAIfW8ToNGJ0SumjyaJB9IzLDdBEXY3BHpBYbTrwlc8g6qcTRP
Xf2gU8Q+28Axxt4sImiMlJl87NyQmaqmzeM0M1o6+WJoEF2OpM2EZXAx/+0RNGkU
yjJEJA60Vx4NdSbX8c/47LdSFqtbo0yRwUukKwU8nRlZO0MWcpJiRH0TgzMGeZ1Q
F5H90n9K9eGtznA3uePpdhI9cVEI31jSORbrJDwDXvah4fpo8yQWEgFSvTn0XxSt
mbW+JNWFCnn83lyeCRLvtGrfdZqscoUBpWGfz6uFHlyrQ4M94vuDQjPbtqMSjOB9
g9jBZRoYF0sbn+z9EsWOkNTo85PcSYXil+M/mVbkaC4AQsW7L5ax6Hfx2TYVhXzO
pAxKCnV532Xar4dvhNGCybfKYNMSw+4y+dNbmr4MtTLnPHRINUTkysaG4jcayu9D
oCnyao/kzzQGSdScrG42LLls8wEvLkva1Q+0cQcXFs+OAWKMqiL9YGAGaj+IKS3V
EUEWRiQFqLRE8XBupEL0bTi4NzZMiPkxeQqvK7M6aWWpjbNmaAMzPgq1YilGkCcu
7DNzJNmeRV/cwbouBt/7FT8sn5QZTjvgWQ2DGAGNhBW816DBEmPLjGqR+jQPV7ci
rfzQYOn0Tn2ro1WmZzozVtP7KfmPv40tcrb6XBI53DXmMTmnfygUqMAR+uWgqgNI
TTN34kZmY2dTGz20PY0Y3SOyWrzVoXMtpKz5iKUNa02NjJyKKAjEDLF/8Ltp4Cts
aEX2VrEKnjEV8p8uIllrau3W5xijnaWYOFAmvhOV07X7WoF9ceeofX8SFn0rMYlY
/iXEYjS0j9H0gP1hqJMfBgOCEZBcofXWywYFfWBM2hPHWEtoyb0eX7UGrmszvQ5i
zPEPqfbW/cbyCFMgtuVF6ZRboT/5Rps9ur3lVtxuJoh3IL68/nia8D69yMyTXZJq
0qx+5r1K9eU7dDkl6128ZGiX+YzT167YvhDCVJ/FC9mT/YCHynJ63KvJVVCSdpz/
1gdqw3SZtfp3KYvj/fxQGo/iDGTBE8SGwG0Qbfaevc/o1sl8XsTHz8E2vWKkcaVq
BxY4nSFVwmSePr7MEzewaL9f6vjFYBtOlXa3bta//tPRLD8diDtEke7vdW6V0qdU
p3B1bnXdtzGWSY7S1qTU2naJ/LRRVC9IL7iy9sL8d5NgMNnQKdYiYOFbKEsrmjPs
qTCPhXByMUsqXL5Y9Dud0WBvcow2vJqZR+DV6FJ5T9dG5ZofIpRiLPcqXOCO8ay2
TcuGzzGLtOrWigarbfzbgh0qrf6DQTy6cCGN69VZeLbEDcm1w7zOsZ2K7ow+QzWL
Qn6dvIYDz6UbccQClYtYhqmV3uaGYWkCt+Gs0boCt4sK68kYOY0IaC407MCwmPAE
w+9sJZAo5YeaVd+Wn57LDkMZ/0Kz0jmW6gyCB2sVHbsUjxGjYGxdAN80KAcrOTuX
sbweriCGmCY64KhZ+gv+eyFWa1VN4/ij07pVbLUAU4Qgeiy3ZwWB6z2UAwkEQuce
bK5ufEk+ZvfnXkxyAyxz7BqakMvLWWkoXYoQHGHfACLykWWLrKgTcNdXppPFie/U
LrBXJmpKVucDaJNU7g9RAaJM6yakEOaEbgiqsseE0VdNjpC/4/fZwoyzh8LikQcI
KZ8PxWAsSex8Z+goQOo8wr4zrCNATLcyv0T94l1yQ1XNiR2v9R2KPO1e7L9NGTsT
60D+bVOzTtMilijSfTgW+EvlJNLuI8WVPqnbIMfgFzT1KtMMja9aoRLBj2gz2vhR
qEkxtLyA+MbG1tK8pALNRYyZ633MajQrRNW1uwApBMFcwOPTyBV2uUyMmMMqTSbE
GhKfkuZOhVaVmwusc1js6ZuKDuawxOdL/roidy3246YsLBiDpwODVposcceG3sDE
x7vALWFv9TCCFG3fas9hu8hzRUa6LYM4TQc9gBg4K6wMWQ4uH89Ns81TzvPahpdS
1QiNLqYpGQHAHMUWHauYcJj8QX/rnEcpSWGMcDK6m5Sv/3fNQgyRQLxxwaTQbcF4
Aw2VhUKhBsj/iNX9+YGYD2QaKNVANHUgWIKmx6efLNwB5U+RtwaeiN5kXwlPxQhX
n8MW69wXHdMB685JDaeueuFblBoLDX4nmSsC5OlcMDtpIW8AhtuKABoD1vi1VovD
yPxSoYnJWYQT+MmcWhBw1+X0W7I1RKbg5idJytCNS/ghsXgGtWUDgGTGrDkaoAAQ
VzuyxgKPeRAA6QML8x0M01pU9fDG2Za5aOyhufaSVVLAO1mUFa2G39ZznkIo/Ldz
Pme4gJLwa5fcvZRkUEP2Amy6YBTC2vLTckyO9j1NHsRh+7FuHJiz/nv400XgnOsV
pwavOtaS/rVKNyKHyXFLK8EqXobqeH3HZqlVFwreG3Nt/8b9RhMAaYy0FuORD6wE
62qtS4WL5MHZWj+b3NXYorTY0u9V92M3mFRHz1Ep1bVmwBj3E7+43ZuY0VgJsvQh
1PRne8tU2Ai/5gdPoiYklYAd9cFl2DZQN6svekr85rO5JJRZrdzcCLHXL+Fnhk8Y
Mj8lgbfeSqvJdCogGxgWow+QFqEX4qCNg25e35Uag8LvdNjh3qVhp/hlYwsgiW7v
yDTNno78brc9uhz0zeTXBQ+0VLEfyWPujpRilU4qyO/3yxO7o/q0k4kgM967jfBE
9sVPZsTxLijl/ihju3Amlac1Wber4NBbzfV6eXEXOzGeSJpc9ZG7rmEwgbgyR5Np
C8tpBmij9KYNzWwl3tUPAispRWLOUduMSZJO/pKPKHNcxFo/UHPXCnzM21B7GKKe
P1iWRt1OHkxr2aXk258xaS1ft7iQ9Z8zYtzvWUB+ZDKCZIj4ZtI2aQb4zDI+oahg
9dkTL736eSgiZQfgKsR5HQRd3hKBVhMfFR5jCuFeWt2v3gHfeqUmJFJkQ8eJwCnl
M332vodHOETzz4Lsizm1mSI5cozv+wPu5e0O2u2QzXxMhPLoPAmU8F9DtbwWWsUK
8GXn1t+66XnPRV4WPJmp1zWoTExh0JpUnRePBWxBLFZy2VSt77ssmPCqagaqsXth
imu76+UluhF/WtrVE/IejDALaD45l7xuYxGpIhGT60+9MnWIQKZFlKNV701b4GhC
82TydVNZ6ITT2zlolc1GnbCQW67VqDZb0cFrNJqcvcz7zdxJoaUE/fTz5zZFGaHP
0HGnHSpj50oQDeBRPlOSwxZTzq4HBsIHnrVAoqng/4cUdjfYWTzKqB5MKMhIH8jC
glbJ8WN1YkWDcHiP/KiswLtubDTJotnCZJmWJBtDpZv94oDb9rmNeKV3f24TGrRY
OUQk427M5Oe2uULOMIQGwSFzZn+uCYJ09TabAV6bMlAF7Z5zJ3AWICWIUI6avIv5
UP5DHryxXmRveUcXitgS/N8XNdBBXTKMhk8gI/PGFg/ovtzhzdsg5aEM4RjCrV9I
KN+Hm7Z3o0o6tPwNJd90eXgQVLtY7MwQr8pNbbaGEZdblyjAJERoAwXlDqti7u1B
0U5eTF4E4KRHANz1lRlWE+lAHRQrHdvUisZpcoOSR/4TFFC4M2elF1qpUc4j6MuP
PmPXB/1PunG+36VmzyKOcqNkustLsFz6Ivlvkbdq6EWV2/zyrXGR6+13jhgK1rdb
/I2GoY5c/4+ZkAML21td57FUxq1EMI0qHAnrqTh8TgsYqgaOmnQdbPUaxzVlZpN5
sHy0HWCh3AMS9tg0jRCeBTFV4eTQMX6K/jj/QOvmlYsZ/emaDRTTfpBB0cCMVlD2
Y2e2xUuGae7XRr4KxU/1uuxZaawoUbL1HPERl2UWVzYYr3vFb93tw2hCrZFRV1Yl
mFmyie8qMHpEI+pedMxLjTg3W3nuvdd9A7Vw0QvlVAJLdJ+rNtAR1polOZXDNXuY
7j87LD5N6Kz04sjNhKaE9heYwB8QHVNu0TqLjnPXrU85x+QdVHhmbtMvov7VfYsI
exBlHpe0jwKNVL//YopQFbX6ZX84iq7gkk5RU3FLX+XFezHku3RI8MiXdWNsud0l
dIS4fYqfHGu5vaiVL1sMRzUknaRTNk9E760ClcCYibS7SkGiUC8FSHTZuxVJI8vi
Ob9Stfo8xdzjZbWqiNzTbO17/iYEePyJlAqLa7EDQa6ENNNJcf3rLg0ebinLtVF6
Y6eWy7YSyjpBYL0U97PZ9jiwRixrMPJF60qOGnDsXul/nNade3RsropQpHxiYJf+
4WhMXF0RwaLSCsgXzgWv7KmWRy6YsYUB49MokyZWhSBsRW+iwmy5XWOThkkZDnw0
HgbRuEFeYzil2DpSALD0215hrdLUCpjPXVY9Ge9etdy5tzXvkr4DP8VX3ngrTwV3
TTp3f9I5ljZppOXUSrcaP6M39x0Vs62l9aS71mxw3Zzi/LaeMx8PFsaXLJeeFskI
LpJDfhVgZ+0PXYg0X/Bi4QaH3msMabASl6CvTg+e+zNe+Y67UmkIf1zPrPJBI1se
a+XqfqT0z6NiBHUgWtcrjb0/Hzg5M+nhmtR0gAu5Fb0M4O6D/4PqF9hEkPPk1kUb
yjgbV+Az68hsZUANW+blcGDa/h1IFrsUWKsE22+/RgcnKqXUS6Kn3CVdGaEny245
qeyUsvqqNri1kE+alyfkYm5goLehKY/KOhNQXXBhDoYAemtNwYylA6hpJJnCU8D9
Rvl0UW0dcsYmHE7e9DUt/Lnh/3TgeRyfUHcgv+LwRUlhUDpXw1MMjFMImFmWuWoG
Hjmpjtw6AH1W/h6j4g6cc5Vrkp5yvCulDJj2oIh2W4M0JEbrCDmSwVO8dUHBswbn
0IyzS+fk9L3ZJPhxr9mNMbuX9/bWvdWnvRd81A1anGx8W/gle1mlCU2wxFcVRJuS
hV6or+M1vS4562c1xN/XwgF4ZzqQfd9rmMl1XzO119f59hr5edlP/iKS5F4ehfMB
EwcV59Oujfcp/p3eutrykbLYPLbLb03xSXG/KA4sc6B6ap1SCY3efeh4OpE2BgHv
CATavxGfrTLbte8XtxxX2ANt/hVG9USaLiIjN0AZt2jzDKW+u3s5IhZtYqPiM/u5
d9XZoGaUgsmVUSCor9sjI2nBALQVMKxcAw/YlVDuTW8WG9Ynf9aTH+atxakAwASe
zIWDdIo4DYk1egqW24K/Se5QeLK01Lxg77pdVhxJ+ldfpaM4+92EiOOZ4ZA/bWXG
njSOT+veMsNCt57IMnd0BuwLyr6XHqgO0FMzbLDKhBl1E5yJ/+VQxEnMZdFHGsGc
fvSfVmMOICiPgFKRTPQkP3ztpyl3vlXAvsCn2saa+FFMG1QnBTDaZajTgHe972vj
sSEsKhpuYb0+Pk6NM4ayExeDHoGtyqT3W5j+Kd228xfOCP1gy2Cd4P/BBVxqtq9e
UNXx8zRSVJhrfX5PLbY1+rb7xmf/ZQa7IjF04gbdeSZP47h3fwybIZHWLs1Zwjw/
+KZDkVbYFukVv59tOkJqvXQ0uSxBtdiePwtnlPYkPMSd8dwikGXeKMhWaLP30TDR
9Q91ZX84jQ2WDU+DWXaDNDUlWdcmmSUjY3gjsAP/bdQkp9NOB3d6c/BGATdYMyF9
tUyuanIke9ACtXz36wSu3LJ3cl/8TTjZkBkDtt0hr0XeNcSMX9FLMDchysIncrOw
jTqRF3NzMW7lUEFTHpNPmHFJaVfkdthIWIl5zkK1OawN56CAVxKYrROuyrBguU+c
DxcxG6ONoiEY0OhZxpdSOzgUm9jz3rqe+dg24mZtNDmUXCX59xk4PpfAQGMqzh5B
8hrE8AnPhOUoTL3ofBV+UqGrSjdLttpRS3pOHjmuLxU5yJ0mUZtSSud/5gVmVDdC
rLvV72+vcVfvJswZBV++OTVaeKb+5is5IRpZzmXsuvZyEv1fKnZPjTSQaqUt3HvM
GvXpuL0zjqKR2wlsyi4NokyBwpGJp+K0un9pHmHitd7HXD+MAq9Rui4lDLsNwzQ2
Q5A11NJ6JJTIfwKcw+jzEckyk8I8i3pO5QLlHUssDPlCBGvG5SRErxYsAWZHz2sW
AEZHsuj2WEh7fj8mk25wwWIekiajOoogHRhIr/UVcYqZU34wwYkUp6lUE9iYXOeX
m/InF7J5CLpyBjezpz++b+ngciH7FTKA5h1yo2mevIJseQIZURW5a6yZbzUC7IkB
Bx2oJBl/CqRcPUan0hXCGbu6fBjtJaxpUIzBnmnIRgFhlQUIOvf0G3fQmjknrV/l
VQlVAU1fjb3/w4KPEq6zlpJnpxrlQWfh5ZIqpw0VsTA84Zj06rNq9NYuAd5LnQ2L
CDarH3ym+DqAZ7tYBCtwh4iUSrMEDNM9nWLp/MSRGUrdwrnesd5yDZpexa0CKlZm
uZ7fNkFzwtENq/C/6tRDtnvICdIrGUsvLaJPpvFcQe8cOIH2geOw1qmJov2biI5S
V6ApnHPCx7fXY3qDZsEmMvlLeoqWwzLTtpqgaB/R/H/lAhDVzCFkbc5mIsURtdzs
O3Z6MAISCFHNjKgoPgBM3uLHDAX4cUDcC+IiBIkeNkb/MJcJKs5QsvFBKHd3q39/
InZBO6T+nHCK0BbfRDFioDMSOWuz8wKniFteUKobvM2MNfMTvILTNsYpSH6Y/1uk
vBzmrdkJpj1ETHfFBookXNQP+JfumHbjWWpb582VgU8GZx5oiIkpJ0zhTB//N/LH
wVJtXwSvsfvnm79JQVj7K1Qvkcf1likdf+oG3z0mfqXylQxfmclFaIlPb4opImYr
5ZiGPOBpr6WLctwfC6VmTmc9LI31eLhBopZ1bBOGhryj/9VOw/b8bgqhG2D9OEAd
8ZSXUaTzY8yX+gVmsQcjYyslV/mwM7GkjWOZbddfawRyEpK+v/kU2sNOliGmZ0UQ
U2c16vT1boDMc6JwcHoXUN1p2H81CBxrYcL2nzIacM2nlKySxfyTUlDMBLNQLrBC
RuuaqcWza6uBymZxDXcY2HUaixizZYcs12JxEMIohgT53fpJjPuz1B8haIR6gAju
Hmg2flKDjVMxgML46ZiaPwxBNAoTWyjp6mvE1fVekTLGCRaio10SdP1NPt3ccw1a
CuRJDNmpYgsGa2HZ7t0dXntsSWBS5BlnsiZszejQj0Hf4gL0C4S91hpA13KP92Oa
VJPTELtZZouTzJOcY2NDyYnsDj1eAtrrfVDRlXwYkD/WDHOICzSx3LeLXmc9qanl
gQOBKL1zUupbFkyGDKPCziiCeyXYgHTRCxzyaJOh/LJy07ra4BJFXf88YsqTqn2W
nr8Zml0UnXvaFTjD52n3cVr6rIFa06Fjh7wMJAy32OhLww4xfHsvtKNuNvlkxvIu
HHRxAo/8Vj91H0uSIqNNQDprA+XfiHGCxECNmdoM4WCuYRVSeQSVpTWBjb7vuPS2
jDRH9cdzbVkiy7XxuW37Wt2+PkerMO2Bw4cGUo1vz0lngAyw19SbwlRX9c/bdGFN
jc/K58bLlLk0xgakyeoix0VRYAWmjTiI71DGgBwty3yCvrTS9jD5pWpmjnPsdH1S
lhuHvdasJaxu6gtIIj807IU3c9EiGcaXKVP9Ch5eH5183UgxlX2KrHmr3gSu35aY
yx7Tt/OlRHT4n3+YDS5YvLbZjQUwIMwcp3sWkUZDUQABc1b2KBe+BzAXZrTEpGVA
+ntafkylwguDUWgY+N5gDFqwIEhzp5R+EUqG//a3cLNgqo71aducIBNyx1uC+WgT
XmQP1OHMJf3GamQN6WTuEeRMB7ubhgyYKs+6XeQS810njVm3PHeHTx0GUWOEqIhv
BcuzZnVQtXKAbORunp2Fhr8WljL3iKgQicPtxKxTeJfsCn1vdy6Njri/4rQbueoS
OAB38+R8Ut1EjyHYeMSpaHlJ2JnWGib15M+VegGIZzP1ySAOIyFnI1QpfoiBXuKu
TtDqRGRm9K5aggdh8k/jkSPzehA7pBO1RVq5p13Ue471gJpEbN04ijNga0SMoPpS
W1KKoNsCq+3qzRlWMckuV7LLuvQvDBVEbtNLXJfTYbJKBvXCPKoYZkaeGmxSVx+r
YprMG5X2uzgsLZGdodu+3AgTqImzjIqh5/3SmRYDowmKmD9DScE2Nv5JeImfcWNH
Z/2EdrU9Cg/JYASJzbe9clbrsdzvXxhwR4FmIG6je8xKRiIG4uNE6mABpnqNozeY
T4fA3C5v+9oPHoYY3elCxt4dgEf+YYSqA9t52eHaxnLdDBwD1MLE1thgFgBohLqw
KRXUrL/3SeD7/JHcq+quwt4e4MkdnyfOpLwnaNwwJ/u2Z2sO3/0lDfrYVJI1h+aN
meJOc/eawhB+JEY5pn1B+RcOFwiT7k0VXI4QlGpm0+GHJdlQQFcG56CSFsvSOXMd
7iK8Mr82aFbrnY0z92Ec5fJXHD/cYkYpjaVJo37ecoKoXnJm/ZldCUzWVjfa8E+z
9uZWrFpuaSbLdvS4VnBZod/TfsK21oQlqq3saYPLYjIJHlI96gOQoyvSx4Han4N5
KNbGH/C48831HaZ4bmooj4WGRe4dvysutpW+G1sY9OSG9+9JyPtAUeODmVbNa2LP
+Nv8377DWKQzCEJtzT2j3awCUtIcHZTCOtRsPrzyBoSZVXlrnrS94vAmeKEVe//1
H38AcezrdzJPmrJ3JX0pksKUqz/K9bRmzAMU/WviOLd8OyL7WyZeWtat8WsZ++4X
Isdw1L+bLMFivuP3kdxk5+nM2sCDBVvLS8VlpwSNX9Ge6hqo1byItPwgz518sKtf
hYPtwZh0MSai9pNQiG2ofJCktTOfv317apYgiMiiOnLNzXtKZr3qwMsPLbo08IwF
K+EjkZgPrgiN9G4Ph74R746IXCbvQLKiWhl/PoF/kQKplfiN3jTqZqQF28pFc1Mv
XFV1ATJmFmTYfLaCgIhQNVxsFWJ8JoX0hNWr9P+oD+YpjYyWJYKgpUm9SU+Pb29Y
6PcR1V3sM46epJxFF4+DYtyq6MTUbeUzlO1EjdNQAgm/rVnq1nL8IUhFt3k5m6af
gn7hQJZhKT0/S5/VekApic1lSLRH9hCdwak8zaIJWkVZcqcAIkrhOaaaxuWCRrV+
21LPVhXV8B/D5z7TCbjlU8uySpGWV/dxN2hJA70hJmG6AeQlXRypMB8yw1Wfk92q
GlpaO+kIASOV8IrGm5BNTKxRusCFXpNLasg6zuAuYvGW8y2lxmjz9bCLUjdqVme+
PD2llU9Zpo1XOqSTG0HVczSc7VwrMVxa24JH7EXjVNQPYUqC7Ly5xZBPXuY9KpbG
3IIMtrjm1RebigePVrwYQavBF108FsIahemd38YbDft9v+agrZfDPrdKJUM5XjJN
SH+/Omxdbqk8fbeE0srMqGpwIKhmhXg26zz8WtMTcX1JyEOoBT/lPBs1B5R3IfSk
m8EV7th/PNLhW6l4CGKXmd1zbI6jmu4nr39/m1otwuHU+HKrC86s/JAJkRbb0DyL
RpYBrH8gdAdkGh+BbDZL+fNL94YAT1pDqgCMd0VIHN0Zn1Cm291uAnrOkahgEuBl
wX7NAUNfY8WKoaUl/a5oXN6YWXngx1/9hzUHJA7wiv0H1e15+oHFrMtZNbdAfB5W
NiUocoqYMC5jKYGMGbif8YqwF+u911sqbYUYLbIBib+q8A02MxkG0KF9cFr5bOj6
EppIcvYDDIJp4IDrL9jAyY8mGAUWBOyayZx0wyJXpkGXzWIBmt7K0Ojy7pGWZJrp
enlZB2w7fXt7I/56AEkY1XaQZdM11wqS6fkGmacrr8+2EZUMpp5nCs2UjwLSGwSm
BsMOBVlGrR85917h8ZuesEHQKDlTw7CzMEBWy+/ey9AGJjKfnTtrKgvTWM1i5FgZ
UtvALPXuaGmr6G8WFC/hjddg525XxLd32fD/J3ffe8AbR/nt6Jd2bl3+NtB3Uv7m
7u8zdJaU5/MiCIFaWVNoU8ShHRipxpgXJBp3+M0CuxBvdK/QjoKhao9rQl20rpkr
9xWOkX4/2ehzr6QP5UZXJeoSRb1k16p35VDfp9KtM0g6bSB0YRNkV9y8AZvTkdJ6
m8PfyAAHyaR5cPsBJdd6wb5lW4vjrUimX7fDhZRPw/rkqU8+1z7sRDWWWH7HHiC5
RXRYBQ8NzT6QbegTH5oIh7smkyhmRH5Oz/mnecWQQjo/P0/hjdT9Ztkxgqg/70iI
kHKI4Y3LevCLwBC8vUu4oDT9VGG7+mvfxptNNchFatERGVfuXzRo8TRI2SZloxmI
eP5K3gqSzDFtermAoRvkQ2gXDyEchpA1DpETxQa6yTNA8RlZFG3NouWdBOl6oT8d
cQ6QpNgyCmGDzzrGfuFZdQMUVYQV+N60H1IUmxrLWhMeqU1M1sMQrROF95e3m1zy
1L442Wj3WY4+/RIHw8xiIZmIUmb6Xw+eooIPZ1cSZ001B5QXGEKqZsNwNrgqpfZV
NNHVJZ3gYysz1zN4p+rNJMDzBB08uKBvZpCsbYAy8q2hDFlmYsrSsjlZ/ao52c88
UZTic2ei832FT+01T1IZM5mN2WqFfEwNutcEplygHUYpPXyggfs6u0MuANbCDksM
6DJRe9fjWqLJul5JFOSCc5vHlJJmbZWGDvfPFi+rDSkRX/OmhTmd4S2ouGcfEUxl
9wryLgp1Xl0fdEYTKR9B/UgdPiesGOZXtIysfF3IpJGsZ6qNn2jdw2DRLw4nBpC7
4NlTQ+h6c5xYigFfVCmznAqHGhni89/g9QL13kRrqLQM30o1jdxaJYjdxovpJkRQ
zZZoNVoLuYgLiHhBXn2lOF9+NHG1pPoOdpZaYDpcq/JtQDefeb4EkfldZ8IoP0/M
+QgMlDpWT8c6ovgsQoJuYrhNdkoyHwPAz2OfigaaMobaTOLeRlHkyBaYR1lIh76m
erWL5rw+DziT9eHnRqHCic/Rj9iKPrDoAWwTMxxLmzFvQV+ZKIEtcEELnoQQYAgJ
UrZrZCqzJ+6f/Kr0WdqgyN8dKiyVgyXKK3cQoJuxYi8e5PTqkI749F40mJJrGeqr
lfKm/B13+RJjt2Ex1VWgtlpuvB0XxEf11awFx0V6DJxsDkQQuVwkJnK+pk7IX63M
f9r8kB56ZF39Ht6K0XY+AYoPMvcTDhLOKXFVOz0d2dj9SeeKZYTBAIw4vWbDqFN7
0K4u8jOszcL1+opXevTlzIo7byvFCQ19fv5gf8E+6VcaUGjYwJ3LMrQhA9l0Wyi6
E3u4eNQbjnBkn77CfQKkQl/g0u3QCcVb6AuQ7znjeBRA9pqd2gKw63lzsTvbh/xs
fsrPkzPqRAqcMSvHFUgseYsHgrVJt/C6SnjiprJQ+6ZrGUeJv4/g5OE3VinqQgjh
0nh6bTqN7t0dh0UDhHXdtmABQBhPQqp87Z9Wak3bwNxOClAUBvWmaNAdthexDWlt
fgr3/xj1Ufe74Vb1oFDj7UW8gUljWK96heWaUsSbVbViJc3x9rGHjYAkhlrRXxxk
gZK+cLr0XC75dEBQnydPJPFVU6AJqGS4OwXQD8PYRjHkvAWfODX6+scYWTSWhgID
qb/OewFd33PF4D/N95cz7sJV0+F8L3zCFXiFXUwve9a0QIUFtICTgK+EqwVenV4o
ywC37pudqriPpXDt+6qTGTw2alxfs31QUTtt3nqfTtmeYpfcMPyegq21/IYwxo3Z
uWuS/yQ5lY1xPGO42OU87RrCTYtc9yGFRRPfiMGnOTw8gPSbU06fkZlOs0sDSJ8b
ro456wPLDvn78JQKwC01rdf3AD0QMheSfynVFdinVtCfqbFfv6oLPnyblZ0tI7CN
rDFrjIpmUBHndzGC7ZVv9NlV2Ap7Jrn2wSZ0PldZ3B/zTucyqJav4ze9JIXY+khw
XEElKR3PKcxVsq0b4SE3oublPe063ic3DxBA47ZY4YZO117yVGUWqR8DTvKn+awl
le30HgdpnmiymMJ1JcRIlmBN0FUv76QO/1yib9nTJB9pi2HVzGKnuICoOILaXbeM
VfbM7bkjDPau13hVCjYvxPsGAdmF1500m2vRO+n3HRGMxgCVzLa51mgA5wIIWzl+
L+wHmttGiH01gmKaSKVBZfDQSHuxvkQOBt75wwg/rqTRLFn9tcLGOWNgXxXtlr03
JgmeiUOEQbp0fHO+SqyKLFFJkPW5WlcrOG87be39fIS3cwIIVYR/Y8TrCC5zbVQT
cPdloIyhfXa47j/iBPlU94HPV6LwX7vG7Vzpkgxq1qx0w+O9GcHEKKBpEmxlesWj
rjd3Fpr8Lp3lcYegywqLxl6s6yqfnY+25RDF9HywmANXK2AIjT+GHZQglUhybqt3
0Szg29+YHQnyLDkGSW8oR/BUN137I2yo7O2Z2spAsLYEBQ+ycp4sKkmSElhgdQj3
nwFH6IyLh/9n3JlQdUSvX8gtpImag28wOAiUcYClIKh+C+YdRVLdZg4ddoX4bnWP
OS4OpCY351CkK8prZLuyby5Jd6qYAtyBbmvqPyA9+Nxz2Bxd6Q07QtAqWgZKX32L
/vgN4XJD3nceVHCxLY419R+XwHxCHITVaXBlBnsy0pKPaEw1FRSZmgQ8W9gtW+hF
VUvSDRw6UxgP/P7H84FZa8mk9P0tRP69FVPj4ev53QIkzBFozESW92eAqy85Ymiz
P7yUQH1TNUoRj3CG6mGZouIwlbpJWadDZFUEmaG++xi4lyOsYJomEk4EUMNH1o6G
9bqdXhPOfVeZs7xrYsdka54FKlPhxktOStS2EXlIWafDXB1/K1sEIqfQ7TVVuGwC
LrnYkEj8+vHGYk3Mk8lZgMCQPe2mndetgQf8Y9zk8mKTT67USY5viyjd3YouVocC
vnvh6Rgt0IwlCpdVMDYF3JrreghdcEc7r07XgCLHgqcdW6nGrmti1NLUeITWFepQ
nrNU4QAcxh9SmRMBpS0qc8qh/Pj+ZE1+yQHCOrH5oFyTdTpL37HhDpaUivWGHE3B
+NTHcSzOxRvatim8vK4vyCQF1P3Xpq/A+8EwRtVE6jhyPrNSlvRX2gpLxgMG9zb2
MzTzeNj/YnG7ftcJdzTuFTXDgKKaQfaOvsepjgI/cU84fgckXFbgdBjgqK58W+kN
CCaFxXJ36vOCIfH2EbQN1dBzzmy+GwrFtQiEA+B0ULkTd4k68+89o6X9fYOJmSKK
8GiFkF7nN7FKvB4O5qvjwC7jLyuYhMR4etsSFcWDj4Ul9HwStxe2Dx8q3NhQwApA
U8fuxW1iWb9vEJgszmefXAAFUhtrQeCNKGi5rkEQ9M4mo9Fywp07K9Q5JvpQNVPw
a90IdHpYZh0yJa3XxxACcimt+HyGNBQhQ80jgzk5YEdFHi/AKFhVTWj69HJESxCe
zAZHztxQDDdYXyhHI8priCvRgIxjRvGadYoQRn4A1J1FFtxeklNWVv4JyeKiLcyj
epDQwXHNd5dFIWeIYqcXqfvnjHUi0aL0nnhsyrPbEJaMz9IssZ0xlBUSXaxHQNWC
rPnNjccluf9kIAV9XyQyduHvp/jzVQ0LepCFRmvLzHNJZsk+TPSqdqZSqRRCSo9v
/wkeRFg6mo7IAxdFaNeWnJ1QhXqIsMYcPc8pfUUfE+r5SkGNPIVETeZhKB6wsbZN
gtuZAotbS21FqRtY+QaS4DmfQs4reUobA6/pgZnUmhBwbK41Q7ScjeLZopZodBGp
yGIIDvVpG2mmGBfV1cACJZpiITMZ2iEaHqixjng27t3OzMAkcHCJ/4VY2OyL+tZJ
wrAopspKHcv5kwIB27nX2cKDtkq797a4TovcMmhEPMjBAT67HnnogyTS9hdjSThq
mN0givOyxpOdUZCVQsgKrldZKwUNZOlkO/DgRMSX1QG2ynogph6scJ7LHMZWcyQY
X2jYEXCpY4qBqqJM2ozLoTkHLpxyDTX0g6A5XNce2/SJ2r9yJZE2vMPweaTyn4kU
XArt8jeMF0wbFStwBqE/hvPlaNTHe95+Oav1e7TOdQhHklmfCq/mK5uHXAczQMRa
KqSaRltkoyMb5NnjzJsbD4N5xMD7WLJmWWhT+2eHmEGzQhrakgW3KamusI2w0kAQ
V9/hpnIMlep3hz3jrzPgADe+jZsihWztbFdo6Who0pRUQ0ukxd48SbjtHuJOVH7Q
L5+7CLY5M3s8ef7gRKcJGuodSc+TFF8mugaI6vEOYN7LVsVU/gCnHRUjdKIqKDkv
7DMSp5x5qwfsfCQDulWsDaiOjPiPZw6nOznWtFIJHGJgKQ0MIlGOBCg1PeUv8Yth
+ayRZg9RzdkVawUdyl2QqMtqNhZdeSaldjJgOhD8hMaGdSgOnUWFZe9XECaZdGui
cb2+2zRxuCXcgIcPt/lsYjM3q09n7MP82H97nyiG/DuewwoZzLYJwxCA53xBXMUe
QF02hrocpLtY+nvzgXP0dCxaVg/UhOTziMBtYG7mCD45xS8oyWbk8IZu+pJl8K6E
jVr80hyksxhz2iTC9xufYlTGwFAPuCRMZDV/vIE1KGm4/eYp7ba/wrblOvOyWhhR
9arzlVHSzUm8qAgLPC5I7Ms1mk7KC50x9bALoyzGKxohyNk5U0C81KjgYdfsrRle
J9H2Mo6vajSuVu2wpncWw+6jJaxt/2v9zKM0eQgioT//IOnxVOAqK4nVuEcnTYe7
85BhI+6JMy8COl3ApfcAo7bkEiYlkO75EhSDHoTnh83keQvO7VekDFjfKqwIhKEa
vTE1XEV3jG7dRS4FH3GKpKnlnh6+wDWX0FHkRT/v7rBz9CohlYhMXoyvpk4CiThS
N+cwXJkXi+3tp5SSaU9Kkh8cCyoXGd5RBbcr9qCbW7o2qaE927jQMd2Ohm364LLh
qDTi8cW1662yFpf7dzaB+oFEjOTFbGq8z6hqK1TjTpCJkCVmfrFGth35vFOwOH/Z
Qn3IYZC9KHZo2Nbq75caRvnSys8KuO0D0GNXq2fM346AIM0utDwytdhoPJfUpyFC
PXN/KYuSVBuxJWn2Jo8aXMrO7r0hImGFeuOSBmiDr4lyQhFlITGduP0jz6yLIpNM
Q6XXDs3m4g45i91vbsvD1vg+sd1k+hJMCrfjRBBrLMEOHxvg+p174gAnGxJ3+s7+
XAPXNAXiapya7nsEI/VEikAVxfL8Oeje1UL1rcetjnDFCk3mH6TwY6emC2CX7FPM
4I7wbpyzlqSwuv+AmuQGeJ1Rs/0cDL9qMqMRJBo3tDDO389MwuDl07UnyjyQsgTn
wxjpuh0gENinChTFPLgaur4GsEZ1xmeNDik/nLzmSP0ArF3qb/ArM28n3ulZijrV
YOMEdcc1gacbNpuBr7+jZXKC7HA2U9g7LIn3zfV5YE5Pm5v3a4Q9VGlDPILGmz4F
BUUQltXn4qP4X2D9SnRQfL6E8iBCLKE2zAZ0yhscXYkgsgPcRnEMk4Qhs5QprH/G
qfC3k5MDI0ms29Z8roeBWqwTchUrzzmFPEvAGlZ8tQ11GdEbDAcoHxhbLUuV86Gd
LWaL/0929+SEPjTjhADMSYTb7p/GAd3di/+D4+wodZC3aN37+hWFKm0UXJbJ4iHX
LL/f9xYdTjew5kRS7gihRiuC7msRgVY25YUQR6cVpEaRO2Ss969hJxs6xwvNLk6v
a3dat7XsuZ1lqba4aKyc5npO4hgUipo1TBP53S44HNgqUyfk+Ax7YBbdluJ1BRDc
ETK83yHoUp65kbHKsSeB1GFLTshXIV0bBZUVSSzkN1/V1Km/G/qnqJeJgZU2p5pB
z9FkIgUdy8PGKxC3wcQc1x89m0xWLrpza0XJMvwrMakLjGutAIkTZnXA0jt49prF
Q7kdtB/AxH3XgK2xlGWsd2qUIfRUS/FxYeVskkxJ1TN/gmMTr7zgjGIrlyhxBFgS
7VMyuVoAHhf85jMdvepvEHQS3Itw+hDyREvG6vIFHdZrPOi8G5t+BUzh/qatT/sl
1q6yhFm/5DZtbwgaUC83XC+jTqSLjxAvxCKCi2JoLvwTse/yPwXhHogYuZO3qJg4
+NRyfwIUXqZg63fvJwg8xLaTnSpwTAA2k+viFmEBUg8Msg6hbKgnI8Ayo6agXykU
crOktgbwlqjiHY92W5/okoaUc330kcK4IJOweGBrk1mr6y0VwBQ4SU01Fu8kJLTB
Fgw0JbF8sAEyyMF/mrRs5tobjvwy9FpoTLSMqQwR50bdrXgDbFKnHwRtAwKLc27d
gQPyKFo4jjWnKZDcaRtvbNPOJl+6ZnU3AQP5o8PnEd+w5GPWSUm5sLoASnLfR1HK
QN3D5mUOS/cS/yN/QPrSkirl+0nimXJco9EuTW/LNLaRANHyuZ/38F+F/4Cy1A4A
Yeodvkc6eZIdwTB6uS0I3Ksqy6JnCedmDNtcmLY/v2oyKG+u+5U1LLWKZYsZo9Xh
6DtAcsSTcrhYUopKjelJgIxdpNxLqfoRuO/Enc9GYW7ixmTByx/iK72lJOlEhfwQ
N7Q4527I/qOoQWvI2Opoq6UgDccqC5FnXn7LsDmjXpqB9ySK7O+a0QJnIW2xyC2v
cNxpagNh8itCc7qCF2iH/+lKpwWwItLkZkR3necYX0hYhoYZbrp17OULnpP0D88d
+mOOkT8hJ0xU3M+d+GuXIyRgO566j+8rd9axPjUmWv/F4uDeRfQPFQnNAlrsns8H
rYUidkg2UlvGRUUnWozHqmoVafBLR+Irfoo/kGnIlTC/KjKgLe3/ciH/AYBTSVX+
xatMDT6dRU/KUIo8AIXE9bvUuUnJSy7lDCCpWe6KYRZwsxANiQSn5R4KVOj1XRip
pwXTi8iFGgmXt3NfBGpzJVt+O/q0vyab0VVlUbsnwKCLTJUudasp1q4XMIpTd2jL
Nb6bO8/X4Z+MX8fr4Fh0Z8XgDQnqA4okYTEeKx+YvSLvexvNHBHM/j36A+Fwzhhb
DJkegotvW0u+rLpgbUpYDLzFLcO7Jd9AKOCnGWjOn14uimuGXKEQ0G5QgpmUbO7e
7DILRChY1JAfeF9DFSLqjUNWwFt80lse4ONufo1qfYaO4Mw2rqEEmFGcidj8uTRw
g9cYj+ici/wPQWxe23h9Yu1OSo6snZOCwohRZSaCOQGSJlw6OcY8qqrzOnBSOjgw
iD86agBZIL8n2ewkO2SnFTTUMpc21jZmsAzYI/llmCxTfZQ8OFYYSnOs1eeYH6Pe
OQ7o/hIIhT66QRhOyp9zzOIHNyeg2e1mdKbPFMmpmkqcPiOWzgu/iIGrPIdHGlvk
TUjdXVQCpiYcsmTLmoamp+ivIIeRiBN7smgtfU9QXH1p9SHx37mPgvbYBAe9wTUZ
PKaMj1ljEP4qzE07jwvIQUDbCEP9WoFba2CX8cWcIHrHwnxymKoqd/SdHS4iN6nt
aPHQweNgdFXjJgvmdd2BPWeaaGqRzXMWy9jv0kPx5gvctyt4+weVvQYN/GcpfawJ
E24GfDk8oV8KdpYT3XLUtTbXIbmYjcA0rueniDm2rZPFo1zwX7Ky4jUzD2NfBRSS
P54/ZH6GPuKOM16YDiBYErUweRvJW156AP10sbKpdAtEm10AMBq9MrMNURaUFEwD
qSi/iBe/di19htADF0HvoXoKbW349qJcF87j08U35/E0KdRorE/n+QzBw6PKKX4S
uRCNGLKKm3XxoNIdH/fcXuZ48QY6DQZAhxnsJDwjZvNJDXHJYP2Sarxpv2sRnzPk
SqyjIWzdEEwltNR7mOdQdnNq9noQhB30wZLclwtiwDRRR0tZZXW855t8mtKMPsir
Iudf9PKoXPp+XmpHtJLwHp1tbcVNRUQrRmGcERaQVBmKQs4LADjgJAGBqqkmrVBM
p8GwRBRywzna0YjrN86+xU7yz+oG7LSaQEwCQwoD7ZaZNBUTlGYEXmqQJFO7pLII
TIwLGTH5YSXi0wLr5yNRQMRftorC+TKwfru4R4dCXrhB+3hhYGKVA4GupssXaf5C
EHeZxci+8cAEZmobRNQap6ljDX42WBynZMSMsTHFG4coXsxR5szG4NN2XEkAqsQl
SVZIQlvXchyoTb15J2/bXjAYqF+jz8YHAvGLVtvXrEAleEmwlZopG5sXkC9g9S2t
Fm0OmD1WeHCJ1mSkXbWn9sYlq3mFXxUSbvVzosFfROAAk+HiRKhL156TFjRFDMaJ
84krHFc7aK3L5iwVf8KdxCODJc15/1Mc3vp/hlSBhJLTWj8jpnUbVYOTh/jSZZu5
EliNgCdfGTa6P9Br7H36BSbaCEbY1TGGdMbn4z+RZED1FWg31vWf2rv9Wf5YfaZY
RYKWMWZvZY9mTgBI8W5k2hA9C1TVCaVvkxt/Hu15OI8BuFa0lswTL+SQwou2Sq2u
7vdBiAnEUQz9o315uHn017euV1qGCPHAmeiJPhZTSzzhQL0MzCQAeVmrQ+qSlkMB
WmALHOF0EB2yYy9+sAksKgWebuiiAIXtENhL6uXoPC8zm4NsIWojFTBtWgBVZZc4
gqv74CXk+LWLY6fSVbXsd9OPAUbAG1Mgm3l955U1aR1Rv3RQvXdoSpQxUMqZOSw4
lXbjFm9Twdcun600+mijuVW5RZ7bdJNFrdAr78qwxLeVrYHmO9H88gsSYadhG1mT
BFU+fg1HjHhVKZunBJ85tfnhT/J1dXNT5dZK1jxFUOoJzzIWlOp1KJPJYyyx5Lif
U9+NFXCJTF4b1GVfG8wIkducNSJNrffSADaCXwQh1qvVwBa9vxkVEetQW/0GvQ56
wpOMyqJL8fCKcIMPeXaVkgNtpZeBNXrp/Klf6VtJCzPTnkcdApAf9S8XLgrK2/oZ
Pp8ZZ6eQo59/5CI2BjAb7UVg0IktjUr20jBSEcRObXPipkM0AQOJWWhpKGAiE2rt
vzdG9xPDhzHTAE8TR6l9H9JnLOL8qSNv6786cHQuvzequ78pnBMbvbraJVwcOpvV
sXTgEDR3n9iTgnjpztUunJOehxqGunuff0o7jkdloL0/mEUtpJ3KYdb38C2fEErZ
JYHfQ87RQZ9xxQp6mlASTiNkYXjOD2NEhiOpoXNnGvMzmzT9s1YhUZb09I1Bf37E
M3WXPIOp+HOosY8G3sJ6+pGENDhneiDlfquPUOauQhCpHpqZlYmNzpV5MDIlgwOj
/rYFn6LnWyIMxl5pnD/OAhFOcvZxn+hXV7qwzUTZodyVlxfF3ujcRlLqrnVe7dja
vcnVRzmrK7QeQDe0dZzzxMLv3MsWh8Os9TfohY4qC2zdC3zrZbPJesurLNpEq7js
1O2U2L+enZLnJAHSbSZFw1BGbCD2Mn1491Tw6mc4p+43EZTaZ8DkHLPDvj/rIv8K
ak641ysLB58zkmJoN18r9fslgzrhYVmGoBQs11s5QSjGVSGt5NGb7o7R/ZFJTJn1
5PxK7T5oA0zTKcJuRnviOPGiw3NE3Mt0DiZItDp64YCxcET/CFKU/bw4l7qPuENA
/JTfWqsoIwChX6R0CCYCiTS08zkLe3YqG/48cE7FyomfC3i6TI5EQgVDNhS4Ek4S
X8QoCdYHiyIV6OU2yKQo2ZcB+XJcF6o4Z7XzcLfyl5boVzbSjF2p2CgtIBbdFQrp
ybQ6izzf/EU3QYefo0xyP48xYA8lrC9KAMfs1XxHhBI+5YQw5kAho6aVP8+/4orK
mak5YsIXqzgACNIDHAoD/4azp7Mn6UtWNvbsu96dDqF1S3oYqND0QFwJN1ry7fg1
tcIYW2faJS7AO7aF3ZhteYMR+TIBRVNp3aVzKkSl5Qetuu30nzjiM1Ki1tM/aoP2
7R3/qkogzqadE6tS9zX+oyiPquM4JzWrHQofKPgWtiHlPWrOiPp23AQVRdaHa5kl
r/yNzi6Ijk0p30MHkfWuuMEK/5cAxITglB43kHQBWUyntLuww/7KfaNGBvVFi78a
b4pHucJvgFq15gFM0RkeXQHnHZE8KpEnW9yQB7Lwvdb7xpwBcig+Nrqjsaeo620X
2JbcqLCWMEVfxHz+77I7/FrAGL9N9QlmrVEOI7AnpU4x1KNkEOriHhO6hZi5/rDd
BzNurK2oSzOohNgMk3fgZWQiabx2KSs7y5m1wr2oBokpi7DTCSX0t6Njkf870TDV
5MpSd35Xkj/BuQXEoPgVogfsceApgFQlglAWQAs9IK1fUab31z9C1NTdRV7a6RQb
lvoUfwkSUI9gxQL7lvwi91eFNeqrr+HITSAgfXT82PtXwREWM9daTvP1kk+hntge
CVcCFg6UE2tSklsZTXqTxxecGwNlWFVxKG1/FxQfqd2vwKw0JXnaqiVVzDVu4Afc
9YsqOQIJPQ7r41KRaBQLCrLKNPC5e2o9Qoc8Tq2UEsrn0/LIrN67PIyU/oonB2fT
HI6fQcLdPXJLnq07cNYjIuCegavoHdYL2ek92zCPL8G7P7r2edC4B/UJplpWP6xA
MNIlk7Sc/Laf5HDySCStEPzNWMxdhNKkw+AXTZLXE9aGAXvzxWnQgbUOqLIUFs4z
H4snqDqfW2dbgkjGn/CN5Wp5wwErS/mxvsBt2Lr9tx5tmKQTjWFCe3D6mwkkhdi+
LnbZdGYmTuZBdet0rIbJ/furcPngOt1/CG6BDf42xg/yLJgca68rIhC4jUICzN4D
YZPznw7rEPTzOADQ38T/WPcu7KUHB8ixaHgH92+0PUlV8nFtZgPem8G/0YA2Twuj
ceSYS+i/qETdJC9+VlfsImVzlO2tmbaiNQF4B8Nrb7bFf3ta/3jNO5Of/cyMSvq4
6zeEumI4GKL95CLAbAGZsimO1MaF01I5o7wH7WC7BizW024/t2JZL7PGjTbuzLN7
p93DC5wVqyeZNt6cbaKOKe3+MQVuhP36E0M/NJjQ6kYXSNhkGoAZpULyIuFWOWBH
rhBcCVRRCGd+8LZomT1a2QpDoWb5451ctyXZQQyP3XEaMObmmeNyit3DtvSerOAG
YZA7ceYoBqcGYZlnNmorMNgDlWngH8LVi774XaAoiMC2lmK7n9G3NjIE8rSdwI71
5nZ/jkXb/6Xj69LO9Lr0vt7wnviLCzjYiBjkUJQVzgm72yhcHd2BHwn/EZTlGWzN
gifirwKWzUGRoWGR/dOUYvPSchkbAv9ZfE+iV00ZqfiqzW1XBmuJK+GgUd6i5REs
pmIEJxRhGFhKQXAQoKdPkOVDo0OKBlFjRzg8L6PEwRaNt6XWvToWFA0104L1h1jD
9VUHaOD/hk5Otmvm18g0nY13DaadllNOYq5j6CKd4bmb+9KWv+xY5aPuUl4/oCT0
AHJ4ZbvnoPAwgbgL0YdNCFc1PZVKWhdAyhl3Z1YbATvNyPVp4myZdaw2HBhgSiAx
hwIbD0E7DhMSlBFokd4AjoonXEcOJNDLvtK7/uehDBrK//sbzWu9q8VMq3rin35B
nOzbQFtRz9Q6acyhe3O4++8WzObGiE1K1c1fBe5WXB2ylGhnQ2eFeNGjTJBDL+YI
vW7JEO/GroeZ60UfCwjTfrUzSrS6+yigEmRFBzmz2HHm1L7SHtoRgRhMBeYG0Jgv
mJEekcy8H3Wgfm5EaIXf4xLu7WpJOp1YD0NTbQZDE2P66k4+OH3I4ggM+03+/11r
5DMG5HSzv2Y7g23cI+/S5hW+KiGGVrxh6A+MJ4nRBKTuXP6fmnkdV+2SJnNjWGyY
xqUCV6bFfYJ8AVDkmatrVo/mDML7aFWnrJQn2Zlh8wpuoCoytfM1N+p5lB0zVO2s
BF0WDWeDA+DBH6YjMiemnXITdVzvqzELFi9NCRT12GIHQSj+3jX5vbEVhALp29CA
c/ygOHwBO/JjgtgAM6TPFd7+G3+/DLECMWOURSHXnJ1S4gvBxOtrTgTsWK208wFP
OvJM5yGkA2+RRC15g2Qh+a2VnnpBr1v9N+gwZd3if3mgV0kbF7RFXUKS0+Yw2nc9
Skr9d2eIcQkVSFFzJ//b4Dx2x8pND4GbmO+U3N/s29Yx6IwrCCXplvkjIUR1pSlu
OVL3bWgWDhIY9R3d3gZ77B5alRHcdMTd9W+mdV365R2ZTBa9VfffV9Iix5dbOmiu
TlURar1kVzMmjkri6x40LFbnbIYxyPSmDLmnQXQnbm2Qyrq8SBfdJrSDabcK9BxN
RbF1td0MI2HhKd8ejzLj6VwrdASYYN0xxh4awDwOiIRlUk8jiWZZEEX0DJPCuSRk
AyW5ij56VugFqJvdeR34ZN64ptyMSxdgSrnUKMOc2BILmvEJo8lig1o6xPbmkJf6
dCSwXv/rtHN2spWDUD4Q4OPcoh4H9OuGyotU0qOHTElAZeO4RE2Zb94J1KM5Pt2L
b4HL5Cu1n8doTw8rSYv0zwF+Azmmkl4VS40mprW0TsHLimmwilhkmKTyvzQw4T9e
EioNJM6mt2zMryHM0Q9epBeNIixFPRCnt0i/QHemMrCaBR9hy/TXeCvp3o/V5j1r
OGWgCV6v+qwqPCvIgVn2qoeROBH+vmMF90S4wDtLCXUa7iyNsXUFMdpSw1XiC9GV
qGE+upfV/a/k960LecUWHQx+8/M0Dc6Zsh5SM7BSfcYcT25evNWgUKnxijHcc91M
BgAVI3CUMXrveRRmG/m0PsaH6AQokGJ9BEWtOSX5eLN9AACV5ZKd24sd+7J1OGH9
o4FdkTinpUD+nIgDGQ9AE3shx/0oALrhtHGBsHnpN92n2dG2PQeka93iONYZBHlv
T9VBDm1zcPBoM9AxOoBbKCaeke3nQOrzQPIVUH3WlXm0YyKymlIH8kLIHX1Eqrca
J/kEzNWWjgmi5EfVRM4felf+H7QfjitzhYU6mgjJn8CJu45kWjAgKse6OdD6tEk8
kjUoVP/7bDOGkDLq25LSjj5GhZ/f4bgGazBba/lYVY1AAC8Gj3OCGWVoesqzMT3b
sfMXHwp66cgrb460X8nKYe2iS269XMFIx1QhHr0PPHW0S04uBoCPQB/eSisOX75Z
RPSByWlQLTiKsAKD8tr89HVz8pTx9g4GMUizP/F82rW0AM/IMKQc9wA4EyyDhNyi
X/QyweuBoEgO3s+m1KbzX0PR4nbqb0wiBF+ZvnHTmF76KzYe1bAUYI8ptVI6q/ol
L7yJUMiq0NLicdw+LJTXrW/+C/KZkmA1IjVfLi2Fmc5lwg4tJCkJwVlheJUVYWZJ
OKHALr/qjbM2GAP1klCcKyYXOawpHGZfOxuSMhC9RK3lDzw5kjKLJIQ0Bu5Ax3Cw
1QkXO5xLUl7HsyEVXTeOoN77J4Zh0kZ5VLAsQcoudmVWWyyDkAqbm1mTfqm5tYbw
5d+9Lxrm8HxakTSmRXc/2riSHRPxbGeVcSr1+xm7Jfc3P/fNoUodIYaMQKuWLbtf
N5218MrXKMuNU39Koo7HDOV+f9+bwxXjOPyAChvJ7QcHIfrkZzEJ7BXf5F9Jv+JS
Dip8YmLkw3mismagxFZM9vQ2SICfaZgIySLQf1CyGC0vW7x+3cTbCpiI6/VtNs5a
oCHiAqXDr/Vvr4232ck8+D9lROtQe9CyT777Pt3GlPltfMZiTlEglkqKK8bQf0p8
f4zTbnuBqeou8aQOSbZadJhjwJx4OP213AwlPrDEVEhAJeRr+aI9u7QSBzpPuTaC
00hyN/g8gPuWJxIh0EcQJfNWyfTEw9Q7PqG85WQDxTbUs1e99NWh02aihFZfD5wn
QIUKfRbu4P2klmXI4HoVU7iSQpU/5U0AiQAJIGCIVIaXNsgejBuFDIdE/Ylg3X0+
RXHzoKEOE1t/tbhIFd73O2OTJqmSMQ6gDerXsZfcyDCoLQcwgRb1lKgo4PZDFMlU
4MyteWJ/mr1rLpNJocKLOdKVgdrL12LjNU+HZuAZgHIJsD52tf6BW1ZZNiXm6tmx
EKH2+TrLOIRgdOqx17PbVaVDZeqKPf4V6j1JdNklKDN6Emz5W1wHsRwx4P8V4yyf
tdxIfg+8gcJ/rvM5ul88FvxEieInYvPaRVlpstDeyu4HHbsrnl9PBSSgrXwCYbxW
V/K1fGyaLFhHIq1TGw362zXv0RXuT4/5mIj04aCiPt7U0N/pEGfH5HinMijmUQB9
EsFiBuJsHGIUsJICDrdN9AIljXwxBNimfxWzVA+BaHeRX4ivSkpXVIHoQmaKsknf
MS6EhKVmbjJBXQvhVUcIwuDh59cLZD/9B1ZJa6hPhDf6gX1WC5oeZxXTiPiPWTy1
9tpJZm9u1ruCZxBPaGYHlfzwFlV6yjOgSZdUYAXKCciw4YsvTrKxzW5co90g4hMC
sCoR6lnEcLxOhywHUDdMhyLd6Gcjq0oG2zoqHoJnY3UWSieW7Ln1Xm828gC8npPC
OOIN9AziR2EvMgaOLmzYNA6XH9BUhthml0aYnNPb1jDimsqvSKCMp5NFFK3y8WPT
3VXlJT8UJvAGXHyvG9LLYca92eWOKrq+epldhQy2/+ydyOZ+2LMGeasZ+aoX9faf
yVBSzg7TXDnHJdTDgTueB0e4ezPWxERBffbF8hG3ArqvdPEd/eIUAVRoaSo3FXAN
tEegQGWEAZIbZCpjNshKwS5yihjgagTWtMha25PHZPAYYKWCqz+GfygvmOEU3H7t
qVliTATojp0TjjZ8YnSVI7pvI+9e8ohcbI7x3m4GPd3jfJ2byol6HwIvsfTlgH3b
Vk4m/oiiDyOzPzHlm6mca3Q3WEeYPSEiDGKD8/uqxIDUN/mr+i645W09PXaY3VRp
MKiAeWmAKe07XV7crs05igInbUSwP1fwaRJv2xhzvPjfaDTE2khA5r4RsR/14v7Q
mPCCvBv4zZugIN9DC7lKn97Tq+5EsFfvZxqwRcr3uvzKpeyMlTLpnHEuEh4Ww31p
slsTi/Q7tB3ZPtIgY5q03kXUYQ1TtjiBj5ck1+s1rHeHeY+5HVclV/egF1CXzHfl
2+Qp90qxmmcY4zIXKx0a/l2fCkxfKAjwF16FTFweT0UvySBj4saqtgla+8UZOwUH
VEpdmW5x9YOuRExlcTeqpPdGtVnAs1d2RX8JoTfwsqxF9f82HhuTV6sgNdN20Wfr
bfsR6Hgs788KP4r5ZS6UqWV4o6vsp/9QVdu2L7hIa+PJnrf21AsK5F52OVmR/BdQ
5gUpKolLjkYMsZ77yv40NLlfk9sUBCiYOk2QZMZYKdeT6sPRapwkXJCJaYx4h8lr
6FJjCd9JEMPxydzt+nDFVwgLmqYE+VM2ddOMCwG5q86LnlC+i6HcHmNmtIFuuwLY
PA6jklLYuTu7B2EDObcektVIyaigpVojkHHeY9ITwNSFcHx/i0h9/K2W/hlOMmgQ
yhIlmQST1nnGqfkTp6Owg361pwfhObHeajpHZjFTc+2t3faS3NxvXro2oxpir4wg
0XkuBStFQOrZighs/IqIxhw8PQBLX1xgdtz1Mc/bs53teH4R82LO4ZFZM+5/PGxC
ga2+uupSzTAWuoXUwBLExsj8V2NC6XvtY2IHUouSyAlONHC/xhE3giM/+hkyBeR4
SOlAARj9zjLWCLXnZIYQL4kuiIdRg/jVaxNp1wGszJ9QeO0qWvObcXtzQmV/MP0n
7ADG48iJXizsK+tqrd0lj75s5ZuKFRfK9NlR3L79cQZjNM52MwGSpkJ5lUZUkXBn
A3gt7lD2cH8+UL2/3fRR5v5djNPx2EF9ZDMbi0nHaQWHw/vdD2f5KoMypqUsiqxk
SkCGEZ1noL0kPWWRpTBQJN2QZd8ruIsRJN6O7z0qLrOCn4BiQ/EI4lilntz8H1mC
JZrAR8UAP+6sz0NB2CCwP0aR4IWhQEtImkWqS96QpOfofI3UR99vVNa3PBU5mSFi
4ILmFt3YtfF0od0A3LRGO94rOve81fv3udxHHGuIZ6fyaQ4q5SRxy3Qm9GfsL9L7
aaXM9umsuhwfUsTAxmyT2umzxIrg5YBQ9nyTuDpHAcFQ+2bq5WPKF6FheJ+e+Jp7
PBIyJTqSjAbuqgWl3FkyZoXqvWJ2M72FzInotIadfDc6rJTccfCeOml6fFsTRn3P
zI4t5GaaCXHu2SzEFLBgYBT121SnLMIKCMh5FAZiKrCQ3GPPT+/9kfU/1NoT5Xf/
eWVBhVzFyd1eFFuPbuxktcbKvSJ3I2tV4YycUXsPzJtV+EkbnRtZdKGr/jv7rVNX
Ge8ygbY9HYcFpmF8ETDbywfaZZiJz2sM7g6doSEYdjD9bxJ08W3hFtb++LlFaT8q
F/xGCWTM4QNHLNqjDaD77tNnN1VPjL6KUeAhnoyAy2wukOXD9CcR/o2Iwt7S5rIj
rcm5zBPhTK3knw3ktrf14k3aytQzON2zPsBnx/oHJfI9QEnaQswPk+McXdEFqen/
Un7x2hs3AJlx9a9UWKcqcxOgA71X5g0/wlXgR74cbL8vmn6aRe+Lb/08szswJgoF
sgHxbkh8GfttybBuMpUI1Ko5NjaytVj/H9FAT1QsxGSks7QX0iPjBpzYKrhdMQmg
8Q+nEM9NcklpHmu5wUELHcZjXDnCXAmOT8foB/SvWU3/EdgwKYBQjsUzJQR8iyx+
/PYJ6x1gITTWZyn/sde0HQZMDm87TDD8X1BpZQ+XNoBVnIu2U4/Qb1PBD/aFr9qx
3tREE1+YQq7lNdqwK3BYiBvZuSp6ctTfJi589vs/+Xr78DrN0nhfMY8UzbrfJ/Hm
fHwJwkmx2HeeIpkm3zRbDBjmXwzl7QWUpXkUBBduOiv290d+F5nls3x8UDV5IiDR
p22Kyy+rSZ+1baXIYtWi5+2CAbDeQHMnBRDDSQKwrkM05FricF7Ln+W/pvFto0BL
VOWpq/RBP8qwt9v1YH5/eVz8nH+RqSNUKrhDOCzsf8GAPzbeYfMG4cmcT0CwYc5P
pKh3aUQxr0uBwydyCn4lVjaPQv6+Zj4fz24lAUmgujmmsEoKWKoUQ70PLzPdi3P1
OEp28ZmDYl37kk1na/6K77bjve1zb4se1r3T3udb0I31uSebLgmFwP6tNW37N83J
Zo8td94bBDi5ppdkcJSGiILAu7xtNlg8uN8ZkOSTdS/TsaLjgqRyFDO/zF65d5bg
YzMGvhmqiUeUHnGYcm7IxQDyZH9nLP9jdPSAvS8KnjHGwq6jMQ6NY9Np+2dQuNN1
zvEE/QgZWEkcPkjGd90y86C8gYtusXQxVMYU5uWeoan55OqG/aJv650lLNxcjlga
KbgpEEjGKi0go/wtaaJbKAckOh+pzcWfVY5yIp8Sz45vVmfilChJKdiaxtP3YbVY
/uowoYeu+x8BhWnoGRcBf6qzJamFOIUQeJ/ulkbYsqT1/5TTyLQuR7NrtSRQy+HE
bdYlDXVj2OCvLrSUcgyVg/iFewi+EplQBGImWP2ZBDFOQblDvG2GJFl0NXpBGkXb
Fa5AeFbG1IJSgE9E4TR7vHw8ogeZ6mNrJYQ5RkqMosvBqfCJOSoHJ4dM96aPGB0g
CV2KfRbl/SDz7kpG9vmZQ1tic+XOUtdiPdtlXEejihtB5GJ+dhfkZBRXRz5dGzQ3
h7qhZotAhAw/ysL1Lc0/XbIphLFgaC5jmuzkoccNAnmOMt3+8uJ2/o3wKsIHDiMZ
jC1Hidz5lJZAiKUdpKRn2uDQFbVOiGng485+WrmIkn5IB2xbfglFNSutnSk5VQue
bYhODtDZXGVYrRpgPoFGGoiZoFtZCT/iRm15cfIlQVdCjSNQmEwP5WNCQf91axoa
pOPA0NSpYPG0JkMHu3NAx1THhGidXjjuHdn2DBpAE49sxZCtq5iBF5j4qy3cQcGU
A3wxyK+8FAgniW54d+0TuOc46jGU1HTzJoDE65dtBzS266lJMUK1wEJQcM0GBwby
gsFkS9rLz3wcHpF0Iskb7xP8JMdhEQaiRafvSRM2OqV/fdgI2GTCPiK4X6SlS53C
6ldwlwe0cH4EeovMp3EOJQPsGtcdhU9ImhdVs8VXpTz6j/I0dJ/P+tf3qmMbSVQo
oyfAcqa8j9NAmY5gfY3WABCCn9RCIpYsKRXS7qE+yFPrhFQSid7D8e7O/m6o2s0x
ilU12RXn72BOKsqK0bhg7vHhN7tdMzXf522EEDY2cOthveLBSPXb9xW88y1ENssh
C5FFlhtH8iG0g2H9jK+YDqceCx0qp10sJ8+9nPpNNEVqHfTgr19w7TGSOip9gy9r
L0EC65nXao4ARBcitjjVEVrMwWDYitFl5XtVoKSgpF+495QU4FBlmLRJ+Kx3IegA
j+pT2MunecMpx5ekxkDMhG4vgyDyn4cHQtgQJEb4QURTxkRlxDHJ13f6yaU30k0K
+j5dSupuzVnw3Rm4SRMSy9HENnBU7J02teu2UjzlJbKEXLX4TfP3X2Zm+nLcP9rt
LNZQ4inAdymR0yqL0B8sRSB18N8fgsjI2W+Tdvvj6hTUCelvcocgDnZyaV6CXAPD
L9FevfUNB1aVWo+T6X5zA0CBUip0MuiyuxvjPQIVSpIXQ9qKa3MWs/HAzXbp4f1G
j3c6+yOysthD53bLEHEMEMIWllFdQdfQhpX+MYuE4ZyjO8oxeDexBNX9Gy6g28RZ
WDuCJ0qN/Y0WrYH04Hqr/m51kTI4q9IC+LZ1hLcFOU/2frpqErUlZJSpgUiV//G4
d0+cSM9rUTSwesO0YU6Rx4wXGKGx9BK3SYz40sXbx4c///BP+jEA0qYJUYRd/q6v
hejRoyi+BdrgvxRxNUBQEB9jZk/RiQn+L6wzfymwawKVf46Lc6d5/sSwp1CzU6KX
4OcFF00Dst8dyHlN5MlrcGOwPWIkxC8PWjFm9cW3ddW5h/4fKRuyOfPe39+dSpPy
ce+KjR6BA83Covmm0vLy+P7navnmRR17eC8zqYQ1EHukujzzoHMXBet1O5424z+M
l/3m6pkb+lsKxXyl2ndYSRvkeqc1b1qmlZD2tjkDJJ5itL22HN1eKdW6At2Rsj7H
Zo4MtfOmyww28HYbRGyifzHuRAXrUXuecVfsa5qkdYUBTXKjfdzrkZtWKcr1w/Cb
PSeaMOmvCYyaObbSFJyV7T44xt8ZcVVENup+7zTFEL75iEIqw9YCfaLU+U2tt0U3
QYBbFu+dKXKSXx3JnrnPRZn+HL1hfU/Fa6yhFD7Vjeoiy5/ExnwDXHsl2jp0NIG9
Oi5amHq/ON+DGc/cH4/1SKTwahBAHkjv2nUb3bIp+4xU+BjfEhn6fF7p6B/R6vLw
4lY1RAbrVV7f2OkMfM35SNasd8QSvsktBPXaNnxwVrAuHnw7UKZ5bNcil/YXOAH9
tC2pfHMjKd7D7MTps8ZW2+q2Y56928ysxfzOq5YSWra3AXFLw/KR2kGGllyVl+ud
TpNV2OhOHoBxLKRGuzRDMXnHtC98g27g0YNdNXtG5iSaSaxjb9rEbL/zaYiWhd1V
o8CVBasQBzqv07rwGIQrs0rtwFmYVB1MJ1EqsLv0m0au4KaEDQOxY6udmgJ65pF1
pKudmsigZ/b+zNV4z6EjaFZtyTFrjAJPH7S8700W6rky2hmbVSn0NmlyM7N8VUKK
RUivft9ldujAQCicI8f2m8XPpTkeJGdNwxaazTiR8SKcY8H3JZdmF8+8milfF/ZL
fVL+wh4s4GqNkgz9gOwtnuGL7CU14PII4TEvNSD2FAm3LVLpqbianX8YHHFO9n1g
Jt6dC0P8GsYThHK5hxs1VFsQiv32yU7nDFlTrHDCY+wjV3Qaf2/EAVu97+a7fLiJ
9BNUah+XfkaP9Qr3Z9jFjtlf/Wlvvihlp9HSYU1oco/RAllaHveyG1DUgZDcUywB
fHyHx3J+FANw58qb81MnM1WgBRIyKnXBLyWv4+F5GgK4LQofmNdUYrHfUkxJ34Bd
NWr4uqNC1qG20fbqm1uXaEQdkT5xC+qlYFXkJnTo7FIOk2yvf8EpWf41gJcxZdM9
rV5W9kV2Y0Ki+arFmjMd8YS4kbJAbmJ0TBo/KjnnC+PdUOKRR0ngp6L6/5URugCu
7wvJTU5XK6lmWNFOzOAoLGn4WqKK/iwbaNlivLMFfapgelk6lyC330Tfr6QYe3hj
r+q0W2RQU4gZ02ouo3BpdFDxshdxddG8s8C0puaqaleEKZmFpxhygha/1BcmLInt
BkHrcgIdJSGxuheLYcvX7dOblt9xTXkrHsBv/QcX2UWBjuCOseXFghAcVmU+GlxN
ybSIcQeRmg9ICTLvO9jd+7xOVdTXc85BC4T2WHQm0XSEatZKd6wMEF+3Q+PQqRqT
RDMIrf8xBA7usTBr2jqQySh+N4iE7upZxIs6Fky3VeVSueE1jSg2KoD6XlS9Au4k
BfG6n14zqzsfabJmPoH0g9kXAuNttnqmuVfYXii5yfvqL9qIntVJi5EymCgtPF1y
GfbIx60VeRzJBwTHQS0d0BBoUJVblWVqYAxqR/bZTj6nG2VLFT14MS+/PSHAYCdF
/YbWhAsTvYLbyJoliVtsGhUriB0rLbgAWAxEboPZBKB+5wQmqD1xOxrO6dQtGZ42
PzTcDj5OwEQi4vKFukmtRnCVuTPCIF4j2NcVlLCJb4jvzpmCmGKwbOJ0uxRVrvB8
d18lvqglSMQ2gGLl4nlukyCXkw4BvQOGaNX3yXAtQgxO7mJS8M/2xrmb0J2/CjKS
udvU8rlWtY80mwIT/B3ZyspYEg0fzVFlXvLPuhppZpya/F5mZw8yrKO5mrJk6Ra3
+gPXgEG5zbpF1dGACdH3iptVq0RENkGc4QD1YKDl1c9K+YE65GxTnioHuZHOh81X
Jp9SpanqGLCWbOJaVXOkJMhjG7td1vh4Di/lN+ngBDja/Od7SqHatt7H4ZtHcfP9
DBMGAHm0na7m0tAY8XFjIuz2+QwhocqxbqS+moDb2mnpJ6RfJqh9DJOoClzbunE2
sO2NrSCaGpL2XLEAkRwwUHdRr4iGajA/Ux9oDrHyxrmlioIQ7u+dUzkL/VcBU4NJ
eMHpDp91NfTNqzGa2+7E8u92j8GHv46szZwGLarfEA8RokbhocjZF5wkFCtAZzTz
WQ8e2WbcwttYTw05VAEd5x5nouaDtBQsSq3lyCbu69RXlLc5rYpVjDMvm6OBKNJn
IS4Ure2bv+0DyQrzOjI81Ef/yV9gOI47PtwTwiTzR+5avBVjDXwD0X3K1nToRC3t
jCZkVptyCCrz4Y9d+GHpOqF/Onjeb5rUirJGIO1jRovy9t1SQhstqiinrtQlojTj
a6r+RXKqsLfZboLU53AbmGCn/XCFbHCsUo8WDcBFv8SIGJVSkrgXwr8x4DkYX0NJ
Y4GXwuga+7UXISxZ3YFwlo4qey5AHHaw/AU8TZUjrYUggVeRE+dFhQCDF+dbnVEk
17baWCAwnqnpCChu5u5S/1xxnP1NxDegzzLEXEkmNYZz5apKl9v4KTslH4FIrOF9
H9c1LUEMQ30h8NSC2M+kvRAzYtfjqdcqOpy+EfZar1GCEBCsjYtsWmKXogzmvZsI
6WOkkW4sqbOBEHdSmGtFz97ZXICqD7xnIW6cyLVI6y1hIBem++U3F9hFHBP8fvE/
WT93Zs84LA4V6eCNSKJuaUHQdtEnGeOFd4vwBoUbw1mgI/K4ONsBaZAN2XkNZppG
SA7v8o/NNDq+tmghHYgQ4BCKMTHgmre+UjN3LJGgOYLo+MqKEwf7SJDmVcrBBf37
5TVNrGyIIXDjsv62MZQPlmR/Ae/UdCigRfKsre7szCdzjukphI1I9A3B5O5eU70/
74jJDDkt+H4wV36dhBNc3eExQCRUmPlIc1YrL3rxe/x2aaz7bhTWvnD482B0/KpN
6RklDGc5d6gZZbCZkWiooQOkjt7CqrWCpbT+rX4DpRxOBZXF+BaIQaKycOzi/wkz
wVcsletMN2Zy1vl63xOG35e+J6NS4pypPhOcdcZQsQ7MekPhD3K9YWj8ZrThgqNg
x2P+jbifjF/gO2rk8t8y30gbgbtzOxJPzJQLVj1OtXCtbyqdUPrbJHKmEs/TWqlQ
1idheMeuXeA4CSADCWlWcElMsLo/iSD6HW7+LW8fs+c620C875H5e7/eY2jO6b50
mAWlFePYhXF2zROErHxa4dFLV6apsUmjPFxP3oEG2QBCavV3sgoE51mUnX1H9tbR
Ab0q13SLlaY9w3MvyWArmgkJKgM/19447B4QFjg6CDuotY7lWXqiVan4ntWYGYxO
S8L+FuUyenqUBGYEfCzfcyWGd084X2mUh4WbEws4WxmXTyaglOgjHfJodPAVW2Ej
MBHGQILPP5HSrPjZJhvsZGVbrGLV+hbqKfyoUrR4bYS9bukOHC/fT8rBcu+xh/rd
aP++hyILCPUYF857lV7u+V4hGpMBvPoqQjS54a7nJH2CJ/thnzFy50SP/hPWgFtC
LLt8gcRY+2QavlNmPngyZ8wAUXzSZ5MQJHN7btafAN+aSFmlfibPrhPkMVp5aljX
YIMkte/nEHURiBPwvM12OexivRX9qsr2kHuqG8ubhmObMOWjvBjsnoepibnvQiym
agPd0NaoxmKMrLiUNqM0t0ofh6B0UmZASbq1cuRHxtg4zI0KSPXKRPPq+Dx16yYl
RIE4PGfK968FMAQP+qMLIc9KS6TKf8pqib3iq4BGg8rOrpmc0yR1CaFQ3y1lYGOC
EszY3lxG5jLfk4oS1m3u3nYYqlATyuU76+U6TE2J18DVaTpoBAGZjvIARn8vgJwb
QET4yz1wZa+OVkVVeYca0QPtTS7Xi7S9tCsLMl1f3cem1+ye7dT+mu/HRv2q3I0k
aOCPCpvsKyWNWhT9Opac/m7Z5Qx0b2DjRCeV2O1FUqarRuNITDTqpgEk7AZiIsAc
A0S4M4BiBS5U74P8J8Inz5sH2hq/1mgmhkbfpY1YxA6XMSAFUp0VTSiNTERGt+50
0RcaGdZnMah5AiGSPZTDqytvVBwlMxeWK6c0aCnH2KzDgTLhOegCQ3z5l8kE+l4r
wwhNTuLxsXZvIwBMevFr1ocozbw2/REhDQyOcfWBVtHt5SVoIMfEGXo1LYsXfUer
JusNf9hCRRIl11KjgFFJatG9UBH3IAXmoUQxOkPAJ3/aayVuzzSKSQKsWsCZJlxK
O2R2PPbrK9Na07HCdt7XzLkXa9kO/3FoUE0wPPuN0ZrpmQ3YR/eBiL7T5r8AxA/x
jv4unE7H2aJhAeE0rJ/Z6N7uOl/ATOWdYlGsATufXsxZ7datCZ/tjfwqOeZSXdvN
6/KIz3fKt2XrQSIqu3Szgi08VTE0hC5P1bbHkqtjrnvmfzQyol5xcFQt/ALkvzcA
QjRrq8aERp5xmZQ0aWO7klpkluvKZUom0tkW2GPAbPZYVZZYCyTHkz2iaOYmJKd+
i8CJ05lZGlzyspYqxYpTBbR0A9EqLX6QxEgEB4pGomUz7j4tHthkQsjkgXupmQwj
YJCjd/t+y0jCRTGsiWF4xLs+BwaIifnFuGKeIg3ab+ak5cnOpcLeihOl89Rb9wMp
VQRGbgVwEr2VG2nFGM4c9jllEEoQ//QDKIKzQ26oqgRr2EvR041yExXwghSNzIMt
wRSktqeVGS+WCqJBFmI9xAFS0iZfJtra4NINN98FDHKN7t8k4DaAqdKxILH5HxCr
84/7vEcpmuz8rmBxixIOhFmdFwBMXA5BftDdjndR1abB6lWzoSMMfN/0aik82B6V
qkmiJzlC728xnN7cjKm8XxtlSoUhwcqcv1OtDHy/tgibdEF5C4n3haoXEvv+f6eH
ZExoB4V98aI3gNK9J6Ub3o2M7AdUPP2+xh4CyOHyg6Acvo88N6qa9rWCGzDVALKG
Edp1WcBnAHWZGicERh+mZbbK1fwI+ZydblWdHtz6rHoNbPIxqL+q2j+JBB9e3RxF
JE8X2UcRYT/tKbfUkByhrGqOhycLbs9gMWKJUDVxO5Jes0AWdiPpLBH/YaaAV4zo
dvr39LhfFCZi/UOoN+fCnSBl4TjhAitK+YlT6746AKQ8ClPodpZ0NOBjRYwGuNmk
vOWJOPVRu2wQ4jgox5rW7D6tzWBZW6LZ6u2gBl3EnXEUrhrr/lUqyJdqEKjgaXEU
8EZRYQDMAdZLe9GObltEOfuhU6Ymk36uGNK/a/+paR3K0/a2CHF7OsZqLEMc/s3U
bjq5extN6OUpLkMQrsCgVi1/S4qX/G4EPCAbAkha/k5moEEl+E6KdBTD2Grlr8VV
pVefL80erWeU8eF34O+05Zj07X3CX793wXJ/8OASIhmumMtZnGDb4jD92i1/uyna
gsQHKIrVL1PeDj17g1G17l1CMNjwOO/BE39mwD9TRovjRWIKhTeOk2uhFjSW2gIo
GTLryVSLMrjhhv8xoA5V4swJgbUbA/eqrmP2ld6h97KoY/l4dRwvLXnEm6a4e1UB
lD0OAdNbNFlrtNImsrKLBJHIVoAROxl4LRnHlvziCMZzs8C7D/OhJIFHxbqu3znw
6gdN+37vLrMOqmEOTu9g1k13N9UzWWlpZRtjVUzlPxg1zAgpZQQYSKNsTFjyGuCD
Ftpv3D4vH54e8A9jHmmuxFuL17mQLE/qnVAW/vQyIkHOhgdng5jJbEv4bdutB1uG
4a9Mw5PP41Ai9XbqpwYNY0BUJfgABQDD6nL4V+nGEk3MZwD0rlHZCSWWjwZgIlf5
Rl2YijrLQ+ipIQxdlBusjdNyj4WepYBOWEz6JlwjmYr/pSCWYzEoKpT1tKfVyNjU
TenFgo2HjluYjNmbI8ITuoADv6BKmG979aWFqT6xk4l6Xfch2EBdLIQmW5KvCcwU
tQpu0PXpVU0aWqleOjQ4xxeCTlUIW7EgPJtS0qLLRjJ6z61jGF8JbPalZjKkxQg9
7zZJTEz3RX47h3xkXM3B3V57EVMdTRQ283NhiB10wJHeNmiwfSivVVg7BOTtQt5H
KUeQ8Zi2OwHZ1R1D0P7i4F9198BJybLj5GwnG1L1canwr+iN3OQHteeI9EMOmEU+
m3mD4QglcJHaIWVBKYg8TUy2uezHmnVNjf9xhIZY4wC8WwzZWMdkD1iX5u9ujtvf
7Xqff//Rl/Olk4VKsQfhTMMqhXglPLNmV6NUBk0r8wR2RLsto0IGMZQJvSAFT/0X
GFsGSYZMHdlSU023w5BCyACC2SD+II86nvzQIq7UAKm1geWk6BqvR6LjXRNQPhqX
PU9q6NQn5BtuzlVBwygW1EIlMZ57B4pdgsOvSyYrZ06t+OkrEGAIoPY9dv5Bug5H
UwlZ7deUB16ihubkG4Fd+TyeqkZRrZTYpzhRq+7Oc/saEn952efFhvD8cnwoHkwl
F0pT3sYolQt839WQwbpWpFqHQjSrwDIHNNn7Me1G1YEsH2GE9qq6c78rOBh1KDsV
WNH4252ll90Rvjvlr5b7CYsmRFOIFczqGJwREKSeQr8XH6wDxwtUKuwA15gokL3c
/XPYIiOHR21Ig7kXpF4ILgZGArfFKkMiWhBqB5Ja84hLIT05CI2SrCThzFjxBv8b
h2T4cERd0wGKgGm4kM7eqGdIVccw+mKqRInPx3T6I7VwNVKJ0PaIQwVAyMPgW53U
8iDhBf/nMg1fQykSwOaYebBnYU6UdqXRO29Iq5DOBye/DFJptTNm3IL5/X02Tghp
GcoWf+ii37kwF771htLi/AIgvp0SzkiXZioVgNSFs7Z84JV92p6e5KQGWGziIZrB
+PG1o+cw9dJAF0izjy+hjTiFu/iTqDd2bNOWZPEXmhQ5w4izXI5hsJd3x47YKEjk
foIQCSmzLTdL9odMaC8/qsSfxwxKBPVICdnEhmm1FQuYgwPoo7JNCygy3zjlJ1RK
GXFFYC2vixMF8itYDCiwyChb1h8eGcqjKkAzhjBwfyB5Cl6DnQpZiCEw5mK6OqLA
NL2TwJkqGWz/mdDwH1IQzTpSoAgFSwPdVFkBFAU3LzgA579K9UqtHxBPZfv4PhmO
tDcCcBpm6l0pGyLJXYypiJIJiFgSRAll2syL8thOZdx9FDUwPnDs4TdGrWhc2klK
Jl0N7CM8h25iRXbpBGzb3nFUuhPLFyfdp5TE3SPNzV41VjCIwXXm4uh18R2kVJM6
sJZxcC0uZ6d0CxsY+6hkLIOcow73nsSyWF6xiqMFrLxmVQ6JK6V5YXbrgiKLoptW
ATVMSeF2mIUJHHn6C2C5sOPtZOErbt2NGYEOsamM1DC+IFWLTFYYt0blodoEsuYo
Q6CT3+XsEuXapZfVPispwt5jyPvrEuwHYsZRe3yQWxrtfuI7RBa+o2q6EDbCkyQ1
NR1npcibfxbtEixeUwaY0/+u2GhO5x43AdJld8/TmGD53apqWHzgTAXuuJ0JH+UA
l9nW1In82DqXMRoNf8Zm/otHY0t9l5wZBQytQLjgbQq5nxN/1z92G2MRON+akWFR
h/55DRC9E7p3YuXggyuWXCjlVkVIb4iuNmop9cOLzeJ+BRnPTxRZpsR9YZEwj1/r
2b9RxrIWBh6Jw9YfG1M6k0JYgKkvK6vURkBKdgnSpnP98Y6eUn4gtq08rfImfTwK
VejJ2ENt6iXAP72DWkvI4Sq0MLDlpDY/IAyyugzMb0dMMaU03uqZDM5QzJxtvERk
Ul0RSNAOFP2Jey+6HbnmF9hM8XIppJcInynQoiv3JApXM2YAlnYNfGxKTFXO0Ggi
MMxBMQIBG8ReBx46SipwFQjYJ2i/hxCTVVS7Nht9E0sMXuzHsZhfdGei4WtNH5eA
VcMa0d959RYwI2g9ZYL1U/d4rZAjXImjZU54ErE+eYUzsgdYIjWC9iUMLdEbJjFh
PaQwJQ2rZ6TdfhkAMFBAq8aShde1pqamqw08r4GKwoGNeXlKKJGCrp0NuUutzUT0
1JG8heKnqNsznyrWXV8CswIkue4HJ/p+ZoWAA+XKwa8KB1Nn3tGd3LxTCXSjMqCh
ZdH1CN36vDEgTnyjaxugADClILatDObpxRkoJavuAGwPS+TawdkmuH+nxRyMAwAu
FggJxCO5WQ0H9PP0zOP+BDEIdUQ41srrVCLiz1jEQNb1bilgeqe6KT9AsaIbwQb8
2aiy6SdaBkcZgQXkxnDKKSaX9zP+n/UDMuwsWVnV5yJH+xAC7dwK8h+FiR7ZnmyA
MRIHSftV7abkH8VjUn/bllwjRrVmKX5/w/hdg2zoi9rqTLXrge10T6Iwv5SrY8ry
lRmCxT2/1LklnfCQrsQVyepeKQkSoFmNuS14F7rWGNVYxwKMQoClS1pYOR1YXAcw
XF3JclQBkSvubOrBdXJAcwZVcvhbVBGGUt4MgBZg1tsIF1BiGf/hBnSnjvMjIQ7I
QOBTI2GQtNK+EYQ8pWJJxE09DeMoiMp2eENumAPd+Q7c3RAVbfQK+D6m8F4MrMgJ
xHFnof1eDvItvn3tTYhJGFq4u2HGtpVYMzmYxTKhxdGCbVvg4Ag77Ht7P3F6B5b5
BJyHwuUVGmICIbWlaEhEbwRsgCnzl40hnywNNAVrNmHz9PfjBbWLeY9ESO8lFKeP
/qk247eG1bTqwpeed/EalNho0Oe296CBRk7plEVxHSWCBL1RsLdUbYq0t0mjOXG8
GFoL9qaOZtEXu/jH+OBP9yCQnBOkDsl9oFLGFy2I48Qe6vWER92uT8ha2QPexlO4
xxv+6zYfbRo146Pmbw+5ZpijbVyYS3BkMKzo3GDo0o0gpBu6yNnh9T3bNhEGjKEe
oM0zC/7zfRJgblIdWs7+sTDOfIxT3qfpSJwNnW2HGGTxNHUTQoW+zKKc/xWvADum
514CKeIrlTYSHTIqx+hOE6NBFTuqt38mshPPuiUlDnqK2pkiB9FgJz8nItI/I4ze
R9Xi1OKy67IjDw02aYZPYPLG7kjrGiYwWrZOwpQ/Uly/Eh91P4UPN9ZdlvPO+8Ok
IWix17C1rVn/5wwZMmJF5xVz9uhv0ImwXKCu9UEnGGg3cax2wfWP0sSYYMaWPpM9
2DmyVT2UMIG/AAC4XornALEkYlADlOFaq/nwQ72Xm2I1PyNZ/ybzwsKQVprU5jPE
BbkLniXB0RBLp9q65l77iQNbJYm2w0uPiwA81NGOqdo5PneCKh77q0xgZ9J8k9uF
puqCnfy/iLRdz+ZO4+pD68/gPBJfxpI7fWHIM93hEGWZRBVJYW1KDGfuA3q71HYV
sz0PLuw2d4MNFfJGqq1i/6BwuHG5Op+ew1pnrDXFvIGCY3SZRH9zGERwuF00AJda
7992N2kxBCLWvZiWZxgq/ll1nVnM8o1kd1YbjtuB2x0OX1dv8JD07ShIcFEivDJa
qRw9gxnspEo+qn3w6/rg5WppzMASq9n/3c588rdeBx/Fhctjg/bdtuCWkb02Ar6F
iIHAzEJ57J5pufBnpe5zaevkNg0J76Aj9wmnFA/H0mwo59Al0maBG+95wc9t6EZc
Nncw/yiYMXrSKbEY863+/Rkbbr4BBUc804bnjCTJ8uVkaHVCnLR8Z6pZuQrTglkw
tW0KRrVT6rBPkh/Efmq/B0UWO/T0NlNOwPpoGg23l948y8lLjdS8Hp3lasLdT+NX
MeV3+rgG2FOojuf/lZo4Xj8uZb3k4mODmZio81Z/TXK3OiWhXhHozi8ZARY0IP+m
daBZw5rbm841AWWTOL1wtG1rWnPqqRuYScZyTU8xwvjYoMshQRYlpOfqHWsibEBg
2XkWPCLLeyCyxsKxXfpoSvyyYDMMXvUDDVJmxI00VZy5A8FHaX4plfQMG9PP5cc6
cj/L3ZQnV0wlYiDb1dNCybkF8gDiZdQdxkZbNOYw0/HJICa9ABO0gmnjmgfJNBgg
L/VkOtkgf8jEIMdqB0ljVZRt4UAcf2fKmOxl7sHBNAJj6Eu7P3GSVS6I6u3mWYev
s3JUre9aFhr/ZTL9ep/nyvks1KCIEa/msU3VJYVMRDGsYjvL2y1DOKjbiLvMBzU3
ibL5MQkKdHLEl0jbb0fvKoVnVsY7tE1s+KvrYLT3TfGU1FtKXfx5fYbW10Q8LpLU
QUg/7bowppgT8GzwAX1jcphpH/VHZKMcvnO4BQvzVagXG14VDu6f5RMg1s0ODaDy
bNcFVf13FnqyI1pU/yh8u/Vcdqpu9MODCB4H5bgGgeZjidMCvddxiuy4tBGR5sGM
ssKMCGDDwQF0A/sDo+jb2VMPVkpXDJx8H11Ljj+k2WxiTNiWUIWCtumN3q1iTESs
WpRY2vKoN3RjgcXAB636NmFdYN7IyaB0osumg/523N3zxiCxbYwNUD9RKC9jtZDV
LrVTrYwLXiyR8x7iNOFndAdW5Q1RqnZjsjod4pBiM0lR58u7k5k80Q0laucDlR7m
vRt7vowdsT5mhnzs1Zd4bHdNZSR+JxPrqPpuqvQMXn9CdZzXxWvNqh8QXW+y4wxa
FEQ/+Jd/SlZZEDzViqWhJa2nZvD1FJhfs/JkrGRklw6g/m8hxdYvxnco2872cRqV
BzYncaouWqwV8EZJXy/84Z71K61DHZYgIR+qnRvpv/ewTGSNsGAGcDLPmtIwcuiP
JwWQmyjqRyjRmm9bJqE0WN//PlFUvjcsCItgicXDZMYCVBrsTrDf573WO8CfeBEt
AcVJM4Ftlud8hCpV00rITdify238JgMlIYqcNZGkI2/JphwwWleI0/NKckO3mwDQ
ifAiMCQpIlNpf8uulVh4CgU8LwQKrvhhAb6D7XkhLFR7EUTKt6lIAuGmqYW/2PZn
46ymoZ8u9Ag4cxPsp7KvO6T7BPD+dFU2XHX8ni8t0xFSUfPKbZAJgNhPDYAGlbK+
l4dCvS8hCr950gsMMHEYAMK9l/oF/kMkqax+0WXoBdbRCkwOSt0pbCOQgduRqH/b
IIfWRCvPrJc4PwSDPePVQkQSn52Sbj/CxNr3ZggpiYRVHQi/5zyBQmmAec0NvM1m
B2M5csEFsv62yT0wnO4MEgPhbGdlX/Fr8XyfiTYO69TRswzCTivcDp/QTwfB6FmU
Ux9WjRBc545euJTTFr1W3AC4zwrP621SrYSijFIgTwfKBrNt74Om/yLzmmfnl7Ay
uV8eKQSVdIJcY+Dx3XParQrB0xcAn95WR4xt28VkVh/qpfCwAhyQy+5a9RttHRnO
ACndZSVNGipIzeVq6HhkQO19JrUgBTQvAu5nVciK//pURSQYnyI9nVX4cxu7QKKx
tWO8LYLE5LNNQQ+xurdLXEaPqmOYX8XXhDUdAqAIMlO42+J8xhj6LZ7GRKUmDmTL
YJ+AAucv+qOQahfoFy8dB1agktrbat1m90aYUF6UKQEV772L/TvtP3ly2TU2vB+g
836hJ13slh78tZJqg2+KEZ5iIt8LZMe7KwYhnI8+WZSrOlnhiHKnp0g//KhVrubL
dcNBLguLufxCDg0sleWRDVDJLRRKCE4lnEZZErNXVLVbsB6FtogS8laarp5YBlIR
9IL2uA75DLEA6n0rjxUquEU3EDKBdQYRqmrNaGU1nqT9bDNwffSbiFXLHrof1Ul5
54blBBgGDy7FoJYCFXmvI9YQcihgaHpsXrRT3ghudfhGZ14otbfXftkp/ZBhDpke
NRMAOHhH0ERmc+DT+nplu98JxRwqWjFRS9Cm9ZeyLoucpqg55gYa3D4TN9mCPemw
r+E7lg3tAwuZtBccuTCbLPqIyrHyW0SuLMQejlIUQN9hcFx4PXC6P/5MmkLFTW3i
bOSFDY3O06YWEc/updjK8o70zFVmAT2gqLGdAH8LrkGQ36eT1N/WVG9EWp1/quUJ
eeakjunkl4O9cPBmeTsIRzgxmVGS2M1YhYQy/aa1wJt0bAx2j3fx3B4y8VATADsl
zXRsKI2wmsxU9thxkgXXGzlSS6zT78E0irK9iATuDuGFSKlwVHPzmAESodyjliO2
HnpubIidvv7v2o8QLF6k7a4jvrREbD6czLmFUp5HRG15GTaHYZOaCLU8ZEhnVgV2
c93cGZ8q2GzmRovoNfJ3FIUC5IZGVbFnXtjogdva1p8VlUoNHiR5I+ANBaakwWag
2oGYlV5kHiXYNe24xoYG6Z8UBZ0w6QHzqqvPmYZCOlQdMfkwNlQFaasig42L3uXl
7M4ModrJJ8o0MmdPO/T+4baBgrRpHzIrr+Y2Hy42uhsEVzpc2c/T2v0F/XlwKJcZ
pyFIU1MO2vmMT1pdhUtOKyWARLfcGtGvt4Gc5hf9IU+xW9jSsbPIfAlkK0H/169W
cZ1L3dVIidSe3pslmxmsznOdfUKSYioYP+rqiPXHwcNUyzCXWLoz/G7cRFVoclxo
Vl6p93mBXuA741tA0exeIIRLqeqrzc+dLKaaWEx6X3gP7o1l+QygbwQoh/B4kCRE
0d78gzgyC5UUWV+qdrDHXwsPbLO+murz7flgGvTCnHgFx6zq7aLrxyXSOvfawSob
qi36Xt2eFMhtFohn005ey5jlKYhnPAcQKlRZ5Yu8pDDETB8zNlCRlarT0b7Ptnyn
aWGA5sbip1dcSFlfkZbY7WxziAtTIaZqPk0otp/0vC6TrMhxq6QlYoQy+6Ch1hho
+E5YpU+thK5s0HKH4ZkS76R5Av0u7g/hJ+Yu1nfRgnv/SpDLvPPbQx8pad0UWf/i
StyqcIuW/0TH4mCLeIoG2OGPGNpZdPyh8vgpRNnSRzENqdykwVoIYB94OpfjMgEc
r+o26RKogEuisqkifR4Q0DULaO/rUlDgTKeoGu7mj5WtVc4JvPvikDJvbrdBx9h2
LXLLxLdhalzUs8ltrEERb8NOoUDIGuKLTKboI80mOTQS36tEq5Oa9VZug7QZVbqG
xskHNEibQ4gEp6qidVlWgmQx9rZRo/QSXY/lMWZrLrfJYLeBy6monD4WExVoCuuZ
zkiK7GXKv2Sim4xqsaX4DklPrIP0aN+4bhxLM2gdCT6Bzvokl7dBWZe83MwOEzyy
6oHpg+WKI5OU66ydaI0XzV6ZsuTlvOvkjJnz+Cpa45bU3fVjByMxb/e90LLcEQLV
dEJEcMmRh1RS7RM4VMfCoG0hAVeY88gwFFGtfWBpx5+kD5MnPlujrSfobdwBA5FJ
CH7eQitzJkT6Ckj1B58SHziLaIOnAomeo23Qh2TnzA3RkH+y3YnjZSJLU904wMDr
MJ+or3ZL5iX0rf+XMmxfuatZ1vUjFga5RbjpFtiao71mEPeoyAH+vDGw1fxdlpfs
MFLDssus9aFTpfo+To7JpdWnM7lhUbNhOnQ4XMdoXCXs1Pu3nj16A6UcfZyHdlZF
dBtkUhzl8U4uVR9KJsfTRy6ticVQPibZRv9xjIv91jSQxuNPvJPCP44MEh5aWz7f
yGhWcWB3v7ubWTqnBgyOeHiJdu7nUvYOURnm/I+Mxxmxw3zh8fLinmOAUPKlairT
0Kh0nOYXitKk8ypaDuJVX554gZVTYghDW9gDmPRtF9B27gIK6PtF6r03aruNIy9t
77j2//hwi9RoAc5M64TrtRvvwH6935mNfzJK7ad+BkO0YYEKWHcaX0w+2Nv4lA4j
ocx4+tqf3RM65f4/GGMsE15/UWhzQPfxTUuTQ2V1s0/6tUoW32p9CK+lkeRGYOD5
9TwyadYRX/8CiIL3wwT1Gc9dZq/SHzyo2OUfgnolqSdv3xBM37W0BN5w2ksTpHp2
XnT660AEHON1cAtMCuDAU+OvliMT8tQ8QyuFiVxIOPVbGkgNO1QKnIOhMdYE7WZb
D45nknsDdw2MAfOloNNSnalsdlsPribnkSLNWjpA5/BAZ54g4Trqo9ZjLRqVxjbw
/qv42cg7G50VoNJfKrqSRSCEi3zVxITcUObU3SBjl6sgcnh7HU9KKqGI3vAbkD+d
JakIzVxYd6BuMqJfZZFTrfM7ommAvt+5ZtWDtC8DlEHNPEhXQol7oFZzPYXfOFRr
T5jKAnp8hqWPnIpAZ92oXQu5JtExQJy3RWmn0yesqU30yNnkoXAfJ2aWeWnv0x2/
3XByLaT/DR43Lk+83PKvFsVOg5W5AKp6jjZ/YvBJJJz3k6RTnmrXnediVPbSONBL
FDlWnlxIrCHqLRItMtPUqMKBjtabnI9dd6/lJUO977wKIT4aR1yTiBxTMspNxBGh
t7EC/VsIMSG219hDfj0tKPqSBaT6MaRboeBcBXh0hUkn49wUJe0h3tJ4ePgtYytl
pSdMNuk9rGHt/XfNl4LpTGmSSxUzt+eiYqdqyD0kZe3MVk6dhb3NRP3+vkq5HEuJ
U0Ai+vjqGz3Y0tUx1e4o2NhGEivzP+itezIcKVJrC6IfRqtMN4Y1PZWzq6K3UFot
bDniv5hpdPdmizBjgtWvTF9zO73J1iLWxYN7T/gUHHdkQ4x9viisNuTkIIn574BN
Q4KrqLluJiNdZjHZGvqm/I/eZkoXrcNlJgiv8j0J1iEyEf6/1qfD2usdyNn0/Vlt
bcmws2UBrOHxjqMXm/D54ID0CKa23QdlnE7g5p3WkTD7KuDe6RbqEZqOgAkvZMAg
X5Vqu8VgXw1zGVVQcIzeCjQQ5BIThV6sELt3EhjNFzo5+R3Y12CwOkd1n8oL7KjM
V5PNx6gXiVigO6z+LXXylIUiy25FEjIHhwgi2umtV99UNNCxEGdho8uGujQ6SAQH
T80QqDLR5BLuV7zSljGJixm70/59PIQTJYLekH4o4KoIVD3bK2LBE08bAJbRrMLE
XR2i1Xxt48ggx+rtgbTy1Z4pd7QGujiBtwB++Sn0uxzh1DcFviBaERO2MFDQCN79
jc/fGOWCpV8vnJGc4D6zpSJhFoJTy7cYRTg2nWXCCqJKbLaWRcWypjXTHpnhXioH
1jII/OsiJh2ZdcIJsoGYqLAkehVUCqpAv3hMkOlZdIxR8C9Dxel833LzpeBMUhNc
AVlSVIDL/2L4PwSpkJiVoghdITtpPljrdk/j2ZpDHQBvq5cMRr3+a216to2bNrUw
ZpxROWYzB9EQRaH3Q7zYosFtGf0wZiF6KrKrGqckehqbZzQjVI5X1BjadKXJvrOt
mSpOp+2DXObKzpo5pIF4NCOStauIwM3EBJcZJhIBbl7//HANLBWVeZdPU6iw3An+
1FxYIA6hcEE98jCHGXYLCnK4ilWRHVoIy3nhWRO/cWXrEjts3p7C28rLumZsyt6+
PNHqKBtn9tuIXoIPnjSCKr0RXlb2rLBeYX7jmNDR2QmHJor+qQkX8ICkmkNXQEEj
PW0B+oVDq56iaxJe1aMGMZEUn+amDXaiWOvaZO8FPSdQRNZPT3k2jRB3ZCDGaXvF
hYbif4mLCQMQXmQMha3zWh2YlY7DPEzBndiUPrUvZ745cLCxNdL7v1mqsvwndMxg
YbnvIarzPWGBp57wk3mStAedrpbF7rwgZ3REcuj+wqUAilugncwLI920gZb1Ikb6
Ek0qqzKKgSU1w0Co4Z4C0Y7I4D4RW/zfATmw0bRF8eolOPtTUgU7ZkixuWHvHT4s
b6sfUzsEhIxqFfE+puDBLcrzxAOHQK0l/Gt5sdwcHQ4n33i/jT7S1JQ9H4hawgwf
ypKYO+Z0mIol42Krd8q8Qg+gWKjpFkrF9qOQE3P4ikz8XImBVA+rBhM8IN+IaK2+
atpen4laUtC5tW0FAUIMCAcgmOGIeMdZPsTc5gHfcm75ECn0/di4Ga5W7p8pty1t
tl/mHc5pkshF1fedwM1n/HVSR93st1JOB/+Gn/6Onb9ZsYyGvrMJ4dq9iROI7OOK
Qs1g06ibwIo5rrh6FOHhe/rixIVKu+kOMbn2MoCduLPWx2kFX1qVOrzZs4SkAPTM
ZURqqz2vrA16QY9NHqMzc2zZ6axjuLZzddxvp0xUn0mYA8YBaqNc4wrwcBmL4zJa
7JFsFvRQfH+EkVRhO6v24SBpga2s7f8TEkAsCm95/6h5CfJUlIKO2B2knH3L3o6D
Ts21uPP5KJuo9x9TqZ8sn4h/pZA+AVliNLwUIyK+shPMUEuNkGBAfaFSciSa4ofh
O0kdIyp/hLTnc5IXjvWQDVcSkxFD1Uc+aKPOCe6lrPtmyqoG23DZneudZATZRuhG
Iwhlex2BRhVWYPCWhoyWn8g7wCYTx7s/qMnPlqzG5mmZiISybzYsGNm5LpTvgd6T
exbRIOmHOJMnSQ101i5pMhNlS5YewioIsymPXJJwa9C5bMWaQEp2eabI9frb4MX2
BhShB69HIRjf+HQqxkmUXLGoAb3OB9PZt11j1hszPagAWHUJTNfkz0VBMuNaoF3V
oYnmcP1o8z2uL8MN8H9shUht2UBEPxply9S5ZAz2VgvnNB4AAFWTunl/QaCOsMdh
qFmO2ROc2jrvw103Qo4OzKVSeIIoX56siigjXHOxCr1MvQfq+Ym79TQLBokCSeHO
IcflAO3leJkYPBDH42+RQDcVCjZixvavtPY/isZjWuTqeiIUK8ou8JztWi8zduLr
EL78G3H1/bWMYQfcuMp6WsN60S34nvoN2yaZeBSpxz+Wy7CHfBHwTtr8LBYH1hwZ
btUnvm72enYFx/hg+wH7IPqcIVwD3i74XBaHtxVYAz+fIsX79mAVGpKu66tGRNcz
+j0jMnkAWvf61SoEX6n2gb7wR+eJ1ppKCNfvYc/CUivAFUxDmvi97pqpS6Vs6CAK
WxT1NimPbbLHbDG8i3hx54iY7n+FhDdNUK4rOGr23MGNhSfNLbzGOdbn/AU+h3Uf
wu5q4fVPVCathWFh4WtI84NW2+1iBfCKnoIiXFKpqwbPehpWTliN6lIgBaWoLdEk
KD8b742HLcK8ao/JSQkxRDWdkt+o7tElgrSS1fp7G+pXBD67kL/03/qoT+qW+eSs
pII4Jrx9WZUa6ejw+pOoPkuPU3dyxS3LemHctXcpNlg5n4j4w9fCU+Jl/eEqPpBO
ZwhNBKwFFwd4AmG/PjEK+hCtFE3QOslJfVsAUvVNVIKhDRbuG5Iv8ZGSEJ1eQJhN
o4BMtnnkERA5vQP3pUD/n+v9oC8Kun+EINObmMbPCsOfNN6oHxgsGlP2XKgQxL2P
VkPax6NJpODkl66no2DgvObUpGK90wJlF1DF63walvpaaKmQv2yt21FZWW62m8yO
ItnYJoGMk0P3stg0tZAU2WXJvthooHDlDLkx0JMR8/hvoAnIEQKUz5RcB1G7bIQX
bNuqx/Dy6Q6/XOEylMD07TIWfzP9kdIZ55AHbJQ1Ed7Z/mjOFejb0oFnu84PVqAj
mOSSRZVmsp9ralqkL5d95zXLzjS9VidY0APhjaPH2PyygM8TI8PYm9/tlfT8h3Bm
danSEmItyZp3ePGCHdhcKayIpwIvSS+Ndm3BNHPo2pByawj7r2u7F+27B8PuV+7w
7q50hIA71Sdp0stwhv87vGhWlRObywsIooovlOKFz8TrIjYbdXQCYVnBYuHGFPMp
fz9CpHrHl2FmKPlMFNeQioViynyxPGYFBxc3+LUNR6rEO5M/A9y0wPOhwd8o0AYc
9arAQ5Ood4gGyyHWbLVejdX1EsrO5loa+kwvnwqSL6X3oW0BdSiY88kFwUNydoc8
dwOTceLxNV8KVCB9ZEMolPh86rnztVPzSk+xi1oxL98IQKxO4oHDAXRc5yql/4iP
nkbIle2dBsX0WLZAuER/KWByMduAh3/4aKh1RAb9x+CsuCLvoWAD+fLBiPHT4is4
0prpmRK9x2rkRsnUSKymSOOAESvzOu6FomlrMz4i6FaYeGMBzvp4F23u9zmtDdiQ
Q3incY4/zi6li1MrSlIjhZtWXZ5HLSBZVx/YTJT7yq9qU5adGKgCqYgF45f1KE9o
jLo2CcTG19lqLojTqd1aMTAz6lAKuJXN9ObiNSeO4tH4fcqXtUttcv8egQw8jO8H
+78X/B00jrbYkXxr8EZpf4jDdcs7WiBSUoiGrcM85tVKrC4FQLRPrZl+/szp+p/D
F43+oVHTS6GKKdMqsxjzTeb2KcfBpMbZ7u8ghZlXPcn3HbsAHDwDvmBVQVQKdJPu
ZnFJmxe/b7C5q3MQPRQ32mJ3sAeiy/seZDSBQN89S226TcqGvK1a3GkjXVNXk2jz
5u1U3WqS/9omf6N08lpeyT7mUnybT6HJvmbD74Ty5cQmxSipwmnAyjmd5Z3VMF7h
zUQqbUiytQtrnxNju0y2FKgyT4kprKHcD2j8J7cnXamaFDRIvaNBNH/inRHw+78s
iLkffiJGKi3PnQM39XcvlKuc3ZaXCTyqD1kYEZZYVJLdolW04gnQs1QxajFcEQEj
Wu2HbnP9JY5oZcYCkq9kNHOrvIuVHZ4IFnAbRa0/Ppd8hCAOgzTbCjqBALjtjMi5
TLp8hcr8ADdAoX/Gff7kNFzYkTNEamR8lAYRxiAJqWwQjolOx0KKQTY1RewmezvC
M/q4ikq+Jn8rvhRC110d4G6lVBAwm6+diSPh15HCgUrcgi6hfrOffn7FG/PXeM2I
yzXIj6puu/h1ZJx5oNtm/mYEtXA6/blkkmiKH5m4345qmmigO/Yndx0vNfaO7U7K
Y9Uh+6DEq7BlonwT/251kAKSqkePWQ7FYxIF0ukYeX/S/3quzoIcB1THGmTVimWj
l6KAwvBwkFGdaPT22rGX2ep28LDJPMFIY5naMZ0LCu8GNU2WDpSZhfT4KjGtlFI0
8zhkOAHd8Ko9m/m4VAgyQjBJpkOVGdJPXIjdShQRfFIIVRcQdX7o6LBjR0YtrWxd
ZfxPyNhJyUnYvCWobjdDYHVugkfxGnQ9XW8ApSwm01sla/SL36OQMur3BGQBQlbM
SnHIEJjJPuxY4Kmkopco3u9CdeiVZBMyrF4jHvsKiVn5crl4wXtk6XQrCA2MaciK
R6nGmF+t4HO0HdIHtv5abLNEX1sgeYWTeVe93rfi1YWjjR1eti+4r15R9Z4WSg0q
YlmuohjMG+m7y06lZ7+URy2yWLTrEHniv29JDBt2FJ2wr9YS5NIEOIxZLS6FaJGn
/jD6H2K33/U6xqGGkfo03p3CL1z7llWEKeEuUQA+u7QcuUL3rLWSR4Kp+SLwSnRz
k0c5/kBH2jKhA8tIkrViVCxsCvh5dRgsco6na87tjADY5HYweRkSvLBxurjbV7eI
oXj/g25w3H8R7hVFzcI4mfcWYeqUfrP105HJmzcPOMQJljA8MNJg1P09EyQTqmj9
WvH/vBDBODWF2oLMAsVRLfMLiKdZ5pB+mAD+uOSwGRXLkr4S3pgHZDLjmi82JamW
78t3WZxiD+hrbXFjYDGTl8GTB7eXkktfu+SUx0NprCnmqkAr0p09YFCLxm8jpXWv
LIlvxZqwzlU6o/s909dSYIExPIaKNXwXXZ62hbIs8FhHUjizrFFqfP8kXl9yvX0c
5azwAzmJVyyTf+YkNuJVBdqMywEBxT1pjFSKV37gCnKmk3AukZWFDETkRmY4XQO0
ZbzgGHPZxJ6i3FFaPx162ze95T6tFJqXnD6+HQjfJwxW6VNgNAJ9p9tCTpz6ZW3+
nOsG5i4wNSWqi2iBKQM3iuWRGg50W+jy7ZTNNkGxyWiuIsc2i7KqwZO9gn4skjDO
Uylgcjs9Wx3uUMfs2xI/OLJIQz8TkJFjqur6h/kVI7Uak6m8dfyX5qB6eQcLe+Jh
G8motQJic4/OlDaJoVG5aW2NG2MFxFN1CL+00ppNrAf88RtVTJRlrjwd7ubCT3IQ
4DuzIr7xeDXgcUHdFwlcDpca8npIFC9Ea2OFSaQT4SfBydP4pRRmGx6SyQg+j/Zq
y01Odf6fmdXII/+NPHTfnHF8LAromgAe/rwNzQRqGUt5d5zUqiWHVPUEXI/E8MaY
LbV575hh5Z0G9W+CfOSq7IoxwTt65ctC2OAc5zF4CzFhWXcOSHdSApGXHomj/fwi
5MXzSpiojSFIBthwbj+B3x7eV4qZQXg8a4CdTrhoWSdLI7U/m5S/aeZO629uEjKD
KgE/q9PLwrSG4IjvKliEopmZM2NOBBurAAJ9waAK5IeVM1t9P03Ji2yw1CrZMgOA
qo7m+ZTylslEe9MNe/jx0CnBOKNqNlzeTqDjH5r6K2FwecwG7JnpRYLK2bBkI/Lu
qgZ1vftrmvI37IMkMwA4RwfK0JAphaSjmmQxU2YXDZ4WeGER8IbhWF1RAXFq/MXP
UoUiiEmBiOIzYhVa9lJHgXfxjGpJymY7FevT85WdUqSPu2axwF+xlk4H2y5h4G+/
M6Xc6K+bKkx3h/vyjfkmF6A1JPxcq3xjTvyDiql3yu96JtdWm8Di1C/ZxmoVkH6P
MujlgfQAw0i9kWqLfloyBPENn2E/rO6mkikLsuq4ZfCuzJRS5UuSHckvKTA+D+3g
Vuiszoud73FKTXXl5ZASCBoR28V4HHq9E+zJXMb7AFYpsuBELayiJaGCnCBPXX61
fCSHCRQIzLQkgj0i0F1cJ1nvr6NPQxlx1BaSJBpcZIS5sTuotHjBiKsltFSPf1ry
qsh6Hz09qXm62A6C64g0Q/HeI91CF54nbVqCXHBEPIG8f/Wbce+zXxtNytRpnOFJ
3u2TFETk10USLk0A+XgQy7gtieATXZ7415B01JyINe1NSEwC59J2reDeWMb+o/Ug
4WCfQKYOp5PC9YCp6GOzVri7/nctW9k08xLIjAsANxYBv3K4XAZmkO3FgjukHHWB
jCbxfvfgsi5Ql5LPiLPRJZCzRJYyAVWrc9/BXUIivv7l0bOj+zkSibKilVt7j7TL
Ga3Fpl5QUHP6EvPwnLgOMNmNYQMSrMt0ScH1SqPiPcK2UxVqNAV0kpEXt/j5AE0r
8ahkwIfF42WQnc4K1yUxEL1/6vew3jlrkRbBcC1BFmlgB4ydYRcnuRPPvHhirvcY
+Ea1baNuro40hJyj9jetRMXT95wZcAxbrJMdLL4/niQXSBfTTGpdcsE2v3WswdiP
biUeLylYUcGqQ1bN/Zyh4cdqPiqKHez2QHEAGM1JYFaP4If9ZGHYVG6N5cOVI2d+
FGlOURsHdbU9vhGzAcdq4MQBtS9GrJUmF7s8hkn47cNM7JMfQPq/uJGykOAyIN1u
mybP7dfw6MOnnTqlGfOdT2f571GMkmqe9JTXyDdMu+tGHrGHm2TAA821aatRk2Tn
TsvBTc6ZFbDgLFrf6z3ixeVqBbl3iC2vtP51QRxRvnDAqZcro7IZ/tKqLqVGcVKu
OJiRlWGka/su8GNLt7gF89+DaknNAdxPzDElyncpJBvkakqpeVrYH0ERSDRlFngO
YTeSKYhlPRoA4sGschQJKK4W2Aru7JXtp5Cmd7lMr/fRLzTe59s8N8nLU2btXtrz
yw3K+tcIOi3dfa1cyb64DDQWmSMLXbUwrSOHQmgeH6CktY4PkORzHbthD+Zk57Nz
Gkxskhr6y04URvm4ODYJXr7bE7NNJkSzjTomk7FNmXKxTu+WQ6L6t3VIu9e7kKPQ
i5gLk/PnGyuiT9+ov6QK5OeTgyL5uhRHViiXpihfGEyANnuRCSYSxKQpyPLd4pnQ
NFArr3Z+h6RZzRoI7DCOoPsV8xYZFSgrwlhirQpvlI4cSio+cJfOEeKDX/bjQsNL
EOAn1786civCe7cQ7IZFNU6pIJOpe3YRSQK4pYl/rnn39exQWRq8d0u7W60VjpVg
CGHXQPyV8O4NJiP55MQk3H17YOQQzHhFg+0D2QQ0CIFESaaTwz5yav/N8wXiWksL
ekAPqhM+ZKpTLciT/wcZcefNQJ7odlza13zGInsUHpoKxIPbcpC9p6+kX45NLMoE
vibbBtJ9/dmQaeZ0PFCAkTznjmwH78YeqhDyFSfPMH8ng8vNUDof/u6jdMHF7woh
tLBfzx/I4VPxI6xU/JWZRew7OkLrT7yHI/hFtviYUrrETfs0cIC6alrH7HsWbE+y
dwenn7BAKcLp1WLPfwBE3xi9TR1nNxNn8r5ihpeU9XeCPOY8oWRc1SFlpsrR4mjb
rfGYoQbDFtALzx0MYRwTObMPGQK93jR9jX5AgooQ9IUDjEz8VlEJ7oJY7Rcohi5T
cUZQt3/gpenjIyoEU7uvQrV+MgSyRqqte08Rweg/bOM9BjPi21H2GeaTTn4o8flo
GzqXCHOnBw8xw9ZSGrqAe0aFoMHNXNrtCMM1bhpBtLW4ossXxMsgdmxF556DGIuZ
SOfpGn48hOKlBkSJArCEhr7ESWG21KvUfxnRJZk5wH+Hsz8KIhXseRZFmbQdnsu6
Jc3ZsBvoujkoDR6KoJ3bHbsNB1tsjPxWTTz+edpG7qVZnej9X5o0NaxMXrK2XCCX
YKopim57ULoONJE94ed2TO8HV81bPzGZL8lm/iSPbAqOvfJKX2vEcv3sgTLgIpyB
vjNL2ZARHpXm086svnADYBLKl6OUiMyn893CB67vscpK5qxrs+Mrt49bE1TF+or5
P5AGkwzB132+4ei1vAlJTmS2d3RwfIQTWciEiPgxYCaiuitjrDm9nvNtbV5EMhi5
Jl3KPpRFS2EugbjV7u4OAfsAFKRnDHUkiBAEvCTMfToG1vxG3I/1ooOKgwcukJUB
sAwcrznZunXi7iI1Tv/zZJqN3V3YxlH9+cJNcFdchWk/A1uawCWC5EeBhgLCcUnM
rGhY32pGcqcx2j7Ct9dxGpYyejyXPT2RJMXvJLRIdr4fERp19oGSVyRZau4O4hj1
mUSODj7hbgOlBut/1NP7WjGQj+gMX5gf/VVGX+pFKDcTRhTep2cM0+U3RDDiuc6l
lrby6PyYf6CLDI6UuAOGTxJyxxfQ1DVISB0L+ZZn07u1vpgL2toGDHyYXRJgf6gC
0hxhP32mDKeBmuNjUp5FFaNteoC0hT6tQloczPXmwx9LEBkWkUfqUR66GmSfKkWY
zU+4YByq5Kh5EjnO4vfPh3q7UB/77Fi2mlgYvLup1VZKa3GPtpLbtZ2X9NzJgV2e
Ddcb7A72cWZ1uwq4NcnujXWN4e7IY/+7W8KrqCoWYRaMQwV+l0tkF/PAf/uXsxHp
UOVby+l5wkYcNat+yOIf4XoFqX4T2IV0TcpQyCV22z/OsXKPx5YduzGWSGBgV3dl
E/U/l5XrZMaVMz6KpPO6aLSsBhHP6mVjsyDlmVtg93ZGGWp/v+9r8CiFEaakx+7E
8p+pEx1MI6ovBMIP+4O9z+X10g/z6kLQAQK9SPwBEbXBcQcrwyNXENd4qD1zZTkm
akM27TmxN5pJqOVxVd9LtZGp6TxB5p6YKXsRCLt9n0b61yXgChtwKIgzoI9zFsmE
MKCXDiADVid4xQ7LJolAznFBUxXgaDvMCD0XPvmxRHrWQKcHccw/2gAjTYq5fT8q
WC3maIKph0zd1IwmF+PJClAXSdCSsMj4QYu+ZSjNlI1CoM7rJ+jqL8IXDUV6QcRe
WKNplDyPxwi3nrqHiKUiF+wPWmI9T+8kRQ7F8uJm47j7JCfF9jp7k+zcBNq0PT+1
4bSGVfYmYrgLKwYn8BuNgM7r9CVzyyl+G53HK9QZBpqg1gv2BhsLZuWN1m3sGPpF
4gVoQxr6wtxbxIxvoFSU1FvJK5OooLauitTCCWZME7j0JaUqcdEPYXBfuRC7ZFEk
lnBVGcWC/oiqNqmxWD7GKyN+Gx1nzCEa6ppv+IbqIXWdeG27FTrCtKH+cSiV6tYb
As9ve9tmJKK4vznv2/LYLjwayNvXmUug8N7ScG2U1V1vc3uzt1BnJ1OJGQk0EAlP
PH8TmXMfvLvwYgYi7LfgeM5c+D1MpfBkJ78fm09mVF3p6CSR+YvjjJYe572v11Jw
N8vrfDzwvZlBMZkaPYZkhFPBxfXCv8fNbWAuOmPJW0c83tpvTRHP8yHXYene82jP
3oo1Su3rxCMmMP8LgaU1VWwvBCcbxwCHzo6jrQHCyeLFe2q0vyhBuRQAy2XIQ+5Z
bAND6SCGwHM4bbxxJvFB5SdRrjCYiFJhf3rkYnsZAtuEE99cd8/PVDh1RwFKy3ts
vojYr4XuAmYJvMFQAZqveXvmAPiWrHViaL/dXgQL+j1vQlglutBkDAjiKVaguag5
mS86m1Nuwuiv5jyMaUNzRVjnxSImIeiaiZ8NOo8+MyS7RpIJKQ+6MZbPm4UWTmzo
RNkMPO8sb5usJFRBoDIyen4278T9pbcXSQm1AW2TBbffxEbEhQI9ZxdNGEWwlAgt
Z0Jhray56c7SIrFMakbJR75vPJmGzOnUaZz7WtIC3m304o5L4k9+XvxtQEqHF52D
SFXohsjHcGLptjqsqjpR88YKo84+xoA1EEno0NExK3iXZKwxbItMdSso+30HA1U6
//bpOaDIHIVsqfkBxjeNuroSnC1NMYftFXr6xjTztaUsdM8R3Kwa8CQBH45Qjban
LB43kcf4Tts1A1h7xzAHKCviuznu7Zs1aFFojHs/e+82wN1EHrywcVqeoN58OtY1
Z/0cbn1lpVujnJe39hRv/+iL4VipS/Fzt++AkRAPuEg5u3/GVCvb5rSasN77gBGy
2sRZiswIxhTw7t53/1ohuuZwedhFZosmlWsBpnH65jn2wLf4KxNe+n2ISd0/oPcw
OqzfWdEnH9DVZ7EiJnUntmNWCbTw+uPWcqtJ/MZf3cDYqCWIuu7dtvRJJmy3a3cx
ZXlixcdYh5TUzAr0BvYqi/6/u1A2aIdjhbPNnFan4FIG5XhR6D7Ob65OyGBF9N8s
6MZ5QKOIyfL0CvHjd1rG7pXQVrQqje7fM7FlO2K0p4FypWh97G1SU4Q4NuhNVhp4
Symk+isJdvsXkfmCVHIIN/K2RoIY30M6uPX969wQ0/dprZsoEEUhlqSSK2jTnUkM
p4xyeStihsNql1j+CoJkppa48JY5iFk4XnIuCaD/Tnqlp9zjHg5nUvADADhfX112
mkrKYNCAmeSwJwAlvE87ePpi5BN8r8FJFSC2Id8/En1jkzqigzZ+rExtArV+pljX
KKbVtDczaTcll68mGKnRmZRO4K3YNTTEIvBP9kQqmf8zsCvF2fBqz25a9aeLJW9x
6om+1aP6BWom7agCLEcvqn6Eoi2q03bzG3f3Eb7e6/avLrZgVvSp0p4YlLH7Twr3
DY8cjwZtq7xxwuQx6dlaoSPDU1UlTnFI1YWVl9XUOqwj0hQPP600KkZSIWhFVR7R
bDayBzTSGXNkzRVAP8D+kJOE/7YUDlfUPvfsWgtS5eFveE4TsRvXDcKxLY4l+keN
oBAoYDiZLT13+sz9vb4jejsC+CNXmL6yXsFsVdPP0g/hhJEW7QEHQiUz2G9PqcmF
EXKWTIvhtgzX3IzT4wAxP4061j+83peb88+Dhe5mZPhHyAQJOk61DJw6IlVhcD00
0PJMnVwJu7rBPLY+qXeEkuOnvlfeefv2zBaQ9r93MZ5lyR77IStgJ7Ml5mCJg/KD
v6FK4dpLP4J5KOt9oiDrUZzCjQzJrtcaLawk3Z3UNm0fqvIMb24kuLqo7WUap+gp
cNu4hJ0Fe4sZOhUyx+w2W/Y36PiCHEUR+fo8X18gOIrDSS7ocksNOIIlUNfA3erE
C0RGdOXci7mLZwknnPpbIv8TJJ9G9VJUwEHJeX2+1U0wYRtG+ZlfahDB3WSVl3b7
hiFIroYSOCNtp+ejm44Gun8JA/XtGqAa/c/B5rDJazeMEySbu7+JYyMcodXoQy7m
AMNMt5yai2+55qjpvya0TlFiV2FQkvt1zk6MaWuxuNyvNT7GHYSRHpkxWfrisR5t
e3p73ntI/J/S7x24iu8ifbTA5NaQCBzzNc8XUaWN4QzqTf6dZGXoBa9lo1Cd8KUE
kBkSWNsTu1eTw+vJnQMa/DY/pKHgEgv40sQGR6d3qC7UBsU5NSrLa9wwAvwBguAK
ZYeXOszZjBtJhdtzz2A/q8qyPx1iduA8JoSlr83E3yl831OrFX0YM0w1lWtncy5i
McnQ7W+JHmyKB2Zbj+EAcH0rZ2BpoKqNcWokx5Y1rWWqC4uOu9jQamXyHDGNWIwG
XBQvyD2klb7G7cfOeNDuSWR6+wZntu+/CLiTG1N3ESFs6S88SEIat1+9ajpnXGmb
8U0obaCoYeOabs79v+et+kF6YZsjQggfnj8/Xml6+pRhU2ZMrzsUIdYv9Cp0Efoi
gMziB5ZlWi3OS0thwZIkIjp61flkjRm1DPiPsIZfmdZ7e41o8NmWrAPx1xZGj6nP
gqyz/Jj5I8fNUFxK+VWFhtHUPjFREKFZa260d7LH11GzQ0h11YwSonEjQPor5lE0
4e5/ak0Irg6MG8q+sSkKUxcDr/AdisH4/B0VaiM7kbwHE9C/u7awrAKuhpNvAN3s
hSA2casFzOCfs0jHtgTikP9FYL3iZ2QLktSw6U9d5LIaYhHMkm48tLiBF4xnm1Rm
64Wq8om6KumwL+XDoTbT7ouDYX7/bZlXn9xPS+T+cu61Xmzy3gjYyLFbA/U1F/4q
R4f832EgarxI5pGDcOr9D+aUqmXlWrmmfNsiPLDWG+WrFVn2GgxYhecYp2MVlSiQ
xkJ0pW5Sz53ZLO1OZX5ZRZD4tT/iQoyaGJyjS+usajcVQEEbcUd9w/iqZKuq3dn7
GWXkNSSA/HtZP5RUkVNsh+512R/XJZGv+ixxj5rPL7r5nNm/yhncuBccrJO/u6zk
Hb1S8StaMRnGVw5VRxN0DWKa1RX7P3DOxiq09z0AMlMppJlrVgpeablduP5y/bgF
Reb3YuejF+abkQgCHteUL3b/xQUR8onqmCDgbe8fZF6GZB3pnyYWcLQETKMcER5N
RYpe9lB4y1ON71g0IsZcu+zIuotsEzWotCTRfx2oE30sEKsj3YlCkEaXKS4NQ/fj
rENTn0kGoC3+4bwenHnmInvKzLbR6E8RqxNeNFcXT6E6TgULM20Zc59Ihv1ZxtUV
De4IctkadVsTRAOCytQV5COOo6uQ+E40tV9fe8g7pgFR1atBZp6Gs2V6MRbSU4kw
tTw24SXwSXs7SiVOvwiAyuoON/mzw8qZO6Kr1L6M+XR7xcHQ60wrS635nnSnH7Am
j0oVOs7vT1rdYhK037rAE6Gl1rqWP8KbAgNSdG+01DfG/B4tvUS4+1ReqXAGD2JQ
9OwAhBPpJbVfV5ovq8vd9jYfeNo6M/P3DbMVMbb7XQ3/MWBUoG/ZjUmZX1iVTTkI
SbOZaRzmgGwQbgSSiqn1rWSjDyfSaaC0Om6Dt/2/V2DejOkGVw8Cd9oXjkl4/4kb
7P9HU+NjVi4yOS58ua5J/9Cp8j2B37d8ZGfbr1Dr0sAB8tdWg/fqteZKRBYTUod/
dAC+Ske0EHq0J9UDFoE1p2K9QIJYEDQvGT2281QZFKVp0ahx6mVxnu+CkydG6Iu9
Bf9dPN1aiabIhVU9xx358qILAYfwd4bqSEv6YSFfRDTqXcN9bUD/vyvxCzLrsKwh
0yRsph3FPCFUWwuxKLZkzGdeTza5pfPse5C+cxIoDhiNzWi1tDyWq92oUkO6KL5k
wSShHRLzKkVEAFKcBPyTe1p09UUYg4azJZv4QCTOK3U9n2buJiLFNlLv7WaDXXtt
+1A164sAqBjebpGiPsdqvwxL3RmhcSD4Ec5aqA1/opSD+1Vf6U7TpgdXAFmzM+Jq
8WWiTR85JLy7KFzzteP0T/jwBNzKhyTogbLH3ATxEbsvQprHxbz8Rk32rL0uYaB9
GVOv4F0PyigZvbEWTXofRnd0LHGDIEZ1ViC6OnNPodeICJQcNzV9cckpuKSvG0Ek
2q03FHs2sWlr5KY2uiJvNAVoNjCTSEK7eB9RCJMvVakXeZuCOh8LZiRNrdNMTmjs
mWnU5MjkzEE1M+QTJQVWugJ2bBjlblSATB/j4Bg/TvDQjCBm6GSGeJsql4IMrYIg
2v/6YI5ATBUNIvOCzAJp1yd56MbEYEn42v3/1Ci1M9aqPsRV7j+gud0ERqO4uQhE
rBsJvtGOu2AvVt605ozvnx/0DZOc10u4a/XDrZB5SyKemi35sOXOBxgxU6g1SE64
OkBpuFKRt4pP04Jp47UGd44sqNY6OEBn1HsSYEmgG2xP8I4q5jnVhzA8yH6yPqnp
MaVSSX7zMXBuxo7JAs31k0xRqqeW8zbEG5PvNEDoApcozviAuveFDPsKHlm+P13G
89hq/zTwgNrpp5kymrCdHhFKpnV8qzhFTwNZi7kD2vA2W6kAP/Eo+hWGLvmSgqzG
r3LQQQ7m0Oa4lY09cxHKeP2qIafRDb5nC0c6lC6GgXcJm7XwcCiYlXJlAGOgGNdU
ebeK8OqfqIpPxv2z+xemMh7BopVTycaJu2Et2M3ddjDcPgboLgZ4EIyLUNS6Ahjj
m5+JuUBFrsd6SjqP3RQJvdQrFCpjMkPFmFmUc+2GY+8eje0ABeh8+sz4OaZ6m6EA
E2bD8TfoeqEdPkDg9uKaSAfDVsOBQDrA9sct41WrcVOYdSTHzbel42bk03LFBHF7
tNCrYTTbiquKQrkaGnDGqeMH1fwbClUxYs5gQRU/I6YoltA758OlQdQgZC+yafgK
H3EcDsjOyEZqXNG1C9XjyVcyRhhTYppEHMnwbUpKu0Y2Jv4rpGnRZtbqjGIyyaik
9kUak1qkx5efkesYc5MgmKsyjAjHGBFbx+B+lAsv6tBPkF8DrN4DdvOZ6ZVPLgFj
j5ViW3lNetwTD6Iexm7kVJ7NQgaAtrNw70QCM8tBERRxAL3HCPtlxxynArv06mC5
Be1FWjav4bGiHUNQ8cDN41qYeQ+WspukQBHcksnfak4HLaDp1WgS8fEu2TilxJvq
aqsj1X6iRCy+mbw82F/yAbwiHRp7PrgobbG5AKhf79rPj3njROaV5Od4pg7gZsJH
xLUK8fck77YJMEB1u5eu01U2m9+bYntsQjHMbwqp0U8mgk8yc1hy79bxQY4BjUPh
2f82CUD7a8CbYj+dVO20LvSV1EA2RpCxIjIZVkn8YAxBYIgI2Ro31YObrz5hQGj1
B4iMi2aCCB5j0svn9+I1+mQRq7XkfGn3g89mCWvNBbv+2Y9zgmaQ/RqDKJXrvrJN
WC6hGe6VB+NW/P1dIlqGSW5ypBSWs+3Bxpogs3mcHeFsqWnkykqC+8zXnlbGff3Y
y6+KhuCsmgs5BtNPquFzSpCAC64KwfDN1B7UIXsCwj496ZYm2yxwL6T44VuYtAod
GVRzJTZDzvUmXaPwTTd8Ok2NFl8XJBzBBUnYEzVyOqTRECtk8AnhU8o2LdCMhOva
DAW96Ef0q8/lk1ueOcnEJC8ktHqRLGnA/Tzl2kDwTtx0xFJl/REM827WJpCfVoND
UTEzoinoLVnX3X176VnTN6e8KeXoDIaBAZJvgmohYUyjRjFTMfpZj3zJrvCBi2dg
pHWOZvy0jPSRUF/ratXunJP/hi1Y3SZKRrwHMK5QLJ/FPxjZUyjoiCcSKmx5ARZK
e5rlzekn9dUFAlNcU2FJlGrKqGdfluyis1isP9IFdlKnel8KWCjjRR7KEuVPpUUH
1ZZc8wvzskxdhtJQCKYsQWxUG88RUIbDHBNPP/q9YeA0+/pYdtzsJBmwDh0Ldgil
OqnymkAcKxq3t+W8qdMJ8HMxb9ydypLDp5vklZ8uyowSTfgQbH8CV/OZm5dzPyqH
PKddcGlfP3yFK/O8qF/L86G8+MhyNL6B0FQykeF+0r6QSjRhYGwtGX1G7eM0hmyI
dvifIZ5tNqxCimmIIGkOnpcndNLcSNn38nJR9D2nwXTb++Lwx1pRYt5GG7mfhZ99
NDDVZXEllM+aQaiK6Qj7MwhY5zjkiHmyHPpyCmaHcaz/Bj1TtcuOZ0Jg0RCEcX9I
KnzNV8tB7Qheym+kQA2S/LEkJema9cR07h5lmacmTVO7CabpavkkWE89WadX4Gta
SpVyWOk6arCr+CWip3mGSX6VK7G7kV9oupZgZkuaEaDe8jBdEu8iVcu3OKP3obre
HJAw9TXogTU2VZyBsldyrE0zm89DomCb+iHyeFBMj0bgmTujW0cFZFBhaVzKK/jl
sAvM0jqAwm+e6sOWH50/sGzwGTsoR9G9EBDHZroiWaYzC7/dbE3rmW3vwBgx5fHc
KG9xDJK6syn9qyG8e8tEYM5BeyVtV2nsiMJUKWoOUpqaFTyiBOLet6k7Snb43C6p
RzndJAsqpniz1OiUJhH1AreEQ4KbDZ/p9uFHrk4TGmFe7N6rYkr9gSKy3E3NX6iV
tkflilDd0YxFg6+uhEzj/aI1iLwBlnXxShzusoyRUwHbLEh6WIulq2q8JeRHht3K
MLTRJPBmolP+jStE+sock7ipPYJqxKYISSNlSvM5JOA5rZmD5XOpoi/G9m7JfEPP
utgbi7vpqnsyFnJGNIoEMAvEE9QlpkV12Yf2H0mKMKTl55M1+10KopOTil5qYE2j
5tJ274ME0b4VRjHZ4A3Udu+215DgX5OGXI67YQbJ2dKRins83FP7urd22mMgWRiw
guxzSD5AeWrc90jX02mH7CtkyzKWpsMaKZ2ahJRGXz5I2d6Dbtrfy4jyuLv8rUZt
Dzs8VjlRfI+R0gleLEUTGa64QOgdIL0463AB14PnvO5wOExqc6/pWkvf+Dhw1JAM
xXWNsxVbA1EWLC0rOFLXhD45JZV+/cYC3nsbGfad0QH3VepmvAG2Jxc8FkKIsiO/
7jwXoxrU76J9ItNiAtB2oYbzZaHrEkZI9A1Ha/mP1pxbw/nU0V8AYt5DNMuw+/ub
6MJ0bhmeB8h8L8wCWms8zqj24HInUpGCAwzAUFPqN7rVTyHBUYosgwOuI3hfQJL7
tp/IyCVgJLnqeDWZSl3tXxJLpl3VDyYsl4r3Ws2DYZ9BheWOb/MrKXd1sWXM8psY
rQqK1n2VClTI5RAwryE0oZCZStcjhLgHMPlN1griIty2nZgSENwt+ReiriVUi+k7
r9WNyrkpQmEHyGXKVv3D7ToB58NHUKtSihcehih3KJWdLlqzRAoSxFFue4vW2VIC
RhOT84AE2nIa3PQQKbJGamuPVoQ3gsHooD29NIKkS/nh20IJqWlloQdjdTOkPUSY
NbVCW5SdqBsPzqNsgLiCbtXhlDY2ZIQWYm/akusbh79kNbNmxAJzDYkfCCAyCN79
PqE81pj085l59tdYgvn+7HkQEuMAk61LeW9ypXHNukl8nnJZhJTPKNbED5tMnVZu
xgfleYrih/W4yhSlc96woDTLXMSS6wqm3IlB/DUsZEptgkB4+J6bEHDJRPmwE7s1
k7z8YTSDKEKKMUYnZHgk1VOMiSItWWe4OoHt5qocD5HDLHrk+qSXqILHyHJ7Jeha
/WmHv6pEu/xMqn6q1CO6+zNx/+M4NLJqthhV1NJkPdAu5nCBgEG9nX+tknpaBIFL
6MO1EUPQGZR7yolf0k/ghm+I4dx4Nx3woW3LgnXk+YoxIvjhl8bscc9rEltvLt6/
cqK3izjjlC/102ZUaEFv3srpU5CkfvL+gnIehTzCfR1YAlYb9uqC0Zj2Nbjjkzj2
r51R+b40G0QfD33dFcBVUMPP6sSrnVX72CCaPp8x7yErQMFE2hoefD0BN0SHIwUV
hKvyGoqVfzXfe23sAzN8Ulk1VbfrRnhsbavjy41rRLNlD3dBZO5zRADZzhzKIlHF
sar3yTnbLGBFmyJBojFUj1W/Lalb+rHAI6/r5eu7l3nvUaGULM7AJeJGq0ohYS+l
lv1di/Z9KDlLzhG90N+MR6H/to6Mbf0ovj6uMuHGsWZRi+gkq4XHwYPxdK2Y4zhR
nREbq5jUGjo9dXwa/k3j5rjeX6iOCeq0QuyCYvfgqTbAdtrVA4RNw5WfpWpgVBnC
npbbvTzzLhPTLNlaQGxSfTkkRuDnZRyQBaPytYvBStolCrMFI5fBEgtgH0N1Gtv6
EBbJVI9FAo7Zr+CBq++dydb0grMlLIGNZp15QmVCZAzm0hRMvkCBx39ykoyMJ6Yh
yIZRhhWfc3el9T0tHf92WLrIN+rnKOf889ChZX6iMlKO8RI2CaQ/Qo0DzZii2FuG
QaJbiTbfpXBMxef3cxQTniMSCY4JVJ7sa7BXtXbumv8jE7kfsi9osqxkQt4IiuUO
xLBc4YlkThFbGK6Z/1aNmLJVgcp2JL3b4Yt/6EZ/G9pOwpau0d6caHkdqzAvVMIO
ojaI3rzGcO9bCJulfgvDUdH+t9e198OYF5bR4h0dJn0GPbq04mncU9vqtBxGRRpP
+nc36ma3VueIjJqrHEQ6bKgd0xUOoWGI/LUQMrWYTKpfmqQ8eSoRZQYb2RTLdn+I
pNN/hRP2KXs3wIW65Ukhbat8n0tYf8nLYskceEDNX0WnFyz4LRlcb4hWqZb4YXFn
62trN1bFZPVUUe4hWlHVzO0/eXCbzB9GUCJ1pIgVaeeDGUeGOvWKlkTJxiXhenBD
Ca9Bl4PGkwsWgYvjUz9Dhgd1hAeePs7ks8uJWQCT/0xl+vm97dS1YtLWCWJoo6Vs
AavkR2v71/qUAnAcSXM32qASWmn6BaXZ3s8+9Lq1kc0Bms+btGTOpZbZdecaABg+
3xPZEtO7L3X/Vv4DqgK1A33nd6LoM3It7IjSiiDlzP+AvFEz9xmsAwHaPpSSOcOT
VkD8+whevIzjqP5LdDC0iOc8zrqzw1yxQ/GbEH9eUhFvCP2W5hBgOLuIqV4uWJfJ
dmqaiC0DhQlMdj2/GTZsjk04Gbhc2qC/7ditGUd0EQMpQo6vaYyCyaAjbOA7SqzB
MkSZdNfuBazEms3EHY3Mo6mMj0joLR1mxGgzBfmfqQj11sjoE2bb/sDsZ07jtU36
HqJy/62fG6FHCeZBed+4TwChT05ebcKczMLXR4PVe53CJNL1MbnOwpeC2iA4/Cew
JGVImDLmWSpM18xwpWeLUjQPXuypybHUwo8wOJYyfIoShvvG9i5uu/4oLE9akk7S
Tojsdnc+3nq5e37HdGwoUvxKw/CpXtsKW+hf0ggJqZH10WqB6hiCgPB0bwHxjdLI
KXS4JCMGt8xcSiz4utOCSKlawJOtOZFjdIgNAyRxXvkgmRRyuJd5rmiK4sBGYi6u
xOtYx+6uypfbDkrrcn6WBwFTRif4WWxYDve4hnMeZtg/g+tJoi+MuNnG0lGjhaWK
6hSaykM1m8MiWfnjs7J4v17x4jLWFk1FPv2kMM8KzfFz72p7e2HzFLs9AdsUxuL7
eNsrwfV7Tod5roVy5LLj8BMCj+7cRqnUOgn7vvxBIZiSMmesHLK3fUQidRJtiOCY
aqEUhCYLbub6Qge46p74WCRJOi1xEr807g8o/4JfjkcGbv4keUBw745ifP34gVUD
dkEsHHI2kULt7OGgLvk5T6FaaT33WP02Zqlrr0mV4/uh4QxNgk15Xq+HdsJ9pn19
mcUhSrRXc8AFkyN756Sbo8rem0MtADdyqasIio4c5ztXKIJMrDGcf8KCqgmlZ+s/
gbI3Amz6D7YtubK6pJjtEvju5DHVlJmaCETniIYuWuHntDjW8KmdbBO7tdZlJeg4
qZ7mUN8WVfRC95kIB931A9xCo2lny9pWzKruZjre2Prf+bwk72kEkTANhwobs+68
AhQ95FsxM2Q6V/Zfbj5p1DFhu3z0sNvEM3N4ZULjZM9zHdFv3YytnOpKKqG4BNne
6P3psHtUKjTpFLXql2UbVAlGY4gErFx9mH5yFPJGyqBwDC5dFt7W0PdDaG9JxN3v
hfyI+coPDeWRoXuz6LKWPwOQjFz4hpz9b5p1A5/01041BZPE8xRjm0c4Zo5qbgt6
YXs9HrF3mIYBxObtfCaPbsCntTrqyEXT+QPjPWeDdWWGZp63vFyj/bpgv+/OAt7Y
pCgQp0cELLCIYt+nELDe/1XMVpwXTiADtmDXcGEtbtbmeeCI5jbKHjuEfuaglvj0
LYpbwl/Ki7vCTHuqqjxqAkQNaGluX46GtDSmb0082JCRff0WK2Nl5Mg0PxQ6CWJs
Z8JS05seX6dAxuiuoETN9kJIvWdzymdhL18puDkQrPme+sk/le3lask6ENCFfZbM
x7MU3HFZ0WLYr09Plb3Jf9LEJ1O6PoVS81LBqGZ7NZHyZpemkakvG+RP35SjYvjl
GG6AWI9LvaMtvJyGEqQGtxP1tbav1mIJkkc9VyZBLZtTGihgoax2qYxgAgNGWVso
2BT4LzmiJxAd6QB5ONwRYTq7k3l2gGzwCvGhJijKgxNiceXLjloAw7l7qGykg2Rx
POw/BNCMGOC/e2QFnZF/9UxrT/4D8E35W4Hqbz/abWCINihej41gx9ZP/3Gv+7Ku
r6pqiNopTG25ON4cNVSTQmPcoyaFar+hQUSOUR72nJedCSWQDth9nzBf0TDyRoJ3
wXyVwyAgZ6Xwi7sP+kjM+5Gd+PmMw0gYcc1jSwFY2ldyySQUBFw8t12mH2a1+RXj
63F9pPaomZn4+Ae7VB8RE8qWXm+N4Aa+mwj1h6uiwrO8041WNbnTKJkeQAbRvFWL
zpr1uEA9C5vdU0X7IGa3+5ZQBhiryYMj56p3g/jlxamueEwbhOIr3tX5J5Tv716b
1vZGc3Auit+eJJ4wlW5HFQ03Y6FMmdWHw80doHvj+63f5KrwvLAx9xO9eWHVLP+G
6hx9eHJTcyn2lp94E3iv/FPZFb7EkwnTVieprcHJdLZPJkks4JKpjYASrHR1j4Eu
7YOirV2d8/thfs8CxnlYQt5M91X1h07KuBlgyZaHeNyAxKbnp+T3AWeHTwZZQbaq
KAu3f8uuF34rfuw6g4SwbAvRDR0+71uEcJuEYfJ8F4m+w3QF8xvfaLdmJfzhnXnK
By5M4SkZ3cHNQ2BERZ8Wx2RjICvVUjtWCHJyBkVNdgzJ3RX3qlYABSYwzKggUQ79
qYyaBvu5t0gZ2TZwrqW5yRC8UszNAfmVSy/EfTa8R+3TMhH0VHmTDVeRBZrTzYvq
0nhbE0D7x1q3TClD6tL9ew91yWV+MDnYHzRj9mWvjn0swAgpITlUGj8IlsNkP7rf
ydCzFEqBOzKjaTh9XiZgGYteJclO/icQIBklbcqfioZErsTI2ZZBg7zopRnigd2m
FtyoADQS9+3uhAsjXbJlMyelZttsh/1jfPLkJgtv5KfWt+xACWB3BAC+KIJtvYP8
+octWyjY1oSfTnK1nZYd+AGqxGy2JAVUFhgId4Tt6k7C90n8Kojh27PLr0gaxUGV
+AeNYi1N/ktoMEIr2mHGZcE6bqR8XZ+a+8pXtYv8iPlaWiLCba0i8HYN6TU/B2ms
wWZmj9P5ubJu5DAxBj60GySNvUbGnNOi7MbtWDRsTPn67CUip/fBC9kNqZOnJqyW
9gG1CXDN7NdWd59WfsyqTJV3pWbahCBs1HP/iriald9nhPilBYFjtg2bbrLKmU2N
+8wWNXqahpH7gOwTXDFCJjR9ztS4MfwajCxa9tFZOi4Y+jHUMjS1lCmahXbgr+lO
mKXd6a61PEDnV+PryeDM/5kCr5McM+5ii00JfEnSKyiEH2/UrfLk9lluQR5wcwUG
TiWxMh6HmJYfOsRoEcy/cGNfkKYWy4R2OMvClDhayUK0nphZ/Ey670nQ3qoBaDoE
uwhnVlB5LfLZe4DYBj5bwXXAqJmPosllaw/Hf7d2X7xrPFJt49h0tifaJUQ9JQ+i
UZyZIwfLOiO8u6+JWQQtxbrdLuyXEFqs6YiFCiACxPSMTjyqL5vqsJnf4BZGsupF
C6kb/CafxnLqzizP9sK2AEy0Qgq7UMbOxImMVyHAvj+wCpN3solKBKpUxtTuRBAk
LIW8zU6P2TkcojGL+86s0lIMHXoxmRcnOvlcCcghmLxqCewFVRnuAt3+SG/2VSJe
fLsJgYi5axAVSwHxv2Li/lXiYMECEXGWdu7txPFg51PXfMaW4HHfl8GvZwObgftj
IulrRlHo5V/yFlUV9YbySV2jmZnEcbMgZEBVFZxH3Q1uBluo2ZV6JonPyWi1YJVH
AaqhPojnFbKbTTpfE/nqLiEQBYWPa5vZJMrSV1aEdSK8dITrXxoky/mjecvTh9s3
MX/kVDIubUtuPCZTD0H14m1uBzGfi3C64NZJ2G2fc8bFfXlD8KlGoT+dIu6auWVI
Hmb86QFwbxXjKAkEgXr46UQJ8JkIdeoQXvKUZmBKCXv7woRyJc2vzXw8s54uiMwL
OA3fd5v7PxiFR8yn84OQ5b//Vb1Lbz6v27lZLLJBKz3t+6LrlHEi2ZP9ZdcQdt+M
MOoK8vftRTQsQmJUtSJCyY6SBWxuLIjEFylPPOgcedZhEC60UBoGv/lZaWzK8Aik
eFLr0fsIA/gZZKMSPgonzjTl0Q2heobJJm+EEHZGXy+N3/XpBkZopPCYMR64pW+p
o6Czj1HcdviiKzpJxxEidO8LBnBx8AXCstBc2YrXxjPu/gUbJQusfD2t9rOwPa3h
GDLY2wsBM4TX7TM8L7bIF9lh+vr2JuE9q0fSW5ZdnFuZp9Te6VHGb9d4zGLeatES
kZpSjGxsFaKnUyxBTqeeejbq+EpgvMcsYIe8wSKK68hgt9iK1l54XQFjxt1Pu+ET
q0TqXtT3g0shRgbHb8f5CqTO7Ds/Ff92pgU0soN37fWGknWYtFsUjEtx4wGRMwDg
OpClmI3E6L5CbuvG7KGed0glf1EbJ4kN+o35u2OZxJ3sCr+PUKCgNAAEwEnJNmZK
afsjMszaRUDeIfIKJhwVf5FtWnHyMCQxMivh2Mrg6RzvTb9SNZW3vtI6V4WOyoih
dIwXo8ve7Sthx2SeGHJ02iv3ls7kZ8Z6ojJk37mdxQlQYicPsfpTEHxtdSGA4MSp
4JeSA8IhxrssEQQm1f0eXh34ADaKnct3UMX9qjLjAW6qF2d6VMQ3uBXxnIQlcLZ6
nx9IkCg8VhTtbTiXIx+7rPonS30vs65qtfwFjytgDdyTnbR13reO1oMXFI/8eBt0
2qqrfSCAxu1pkmRbyBM/OvDl66c0kCPUaPRVyDAQDu38LryN0RZREY0J5nCHfbdt
0tyPnxrG0zUuZ66Rx1YlCkel/mJAeUhXrin9chmOSKQsTWG9enf0FPVY6FiW7K0Y
GQWuOkn8aTr1JkI/pLMBzGja66Elm/9elHsKd+CIraH49ZXWp/0bXvHpd18nqvy4
kXaK3HrajvYhWySLiQRGxOcp9gsb7Ip2Oq7JODn32mTFxQFePNgkP/80wuPXDQZS
5i0FiVh9B2SjFRucWd3tli7bqLRRfP7u/niVSVXqJ2MSjhB9NK/ppRnjjKjrh7it
R4DW8MTmqHF9s4ieckXx8KdCujD9bd0VxY2EQ3iB+nMyokkPkMnLXw/9g0yorTHK
Y6m8ejFcGnRaDJSnDeUj0VnMIaDzHYfJzzkrDS5lZ0PXb3oTleESoKSzFyQacG1H
ENhIhy1l5tIhfqBmYrZipXS/oJ0TeEtrnAwYK+mGDbWMCYufvAG8FiWXiwfmIXcQ
D+/fVfacC1ZHqIk++aV36nYwsPHWNrIrY9FLqaNqwpINtHBVDY18fnPNmNq6+Z8K
ULY/zr+i+yfQXxbcwDCOXwhK9jpmJDRAE8gGN5f4LFKPWWlcuKvthnRdJ1nQBHwy
VIGWmHeEI2l3HTFW1QalolFZTrQH5uKfQcekFILoELt6hAYKMQXF/MtG+o1Rp5iz
A8HfJ1jgslC7n+vh1Es0jx1Que2maCT7cIo3iMyL5XzP6cd2kR/Np7lS9OxUiH1h
38jxrGqjpN7KYNbAS9SVwbZK+tsYLDHDvdoH89CDYR2DPb4ZKerfWQ3IDh7Q2WFp
TcYz2gGyh1VKYlrDS6vbC42dYIXF0cefABQAU7IJaHADeG9jsDkqgQk1gcirUXy/
jehzsXiO0ljTWV8RpQMZRiKUuiRoYLW+3iWs33t6muLVYQv1yQqwsS5IdnwVim2W
Joo7j6RDxiER7a8MvmBCUPvzkzWV23HW2UsOwuFQRBTEDaiR16eY5Oj86J7vscYw
TviHzB7yURIU1qWSTwGZZ5fprmz3QzP9ePmlhdoEjea8UDRHFCimZmKb/3gbnJ6W
bXhD/CK/voK0nsmHkUL99DTG2IDTUqwW1faV2zOZ81pR2Ng5nF9zLG+44lZD/XhF
mXHpQ22NI0qe3kepUOiOJsHCnjNQHsx3NFhqC6T1xZPLJfgDjVn3M/1mI+7l8HLj
cAcbeCPNp47t6ZSUO+JzK14HqV4/dhHFDnY/Mu/Nl3ycBTijN5u5LNPXcLb0NW3p
XywDdsb8AiGCL7dzF8hNAKkHWBUTx2ndmRqLyRrGAApIyRCL+STBk1e4gbJjNoUa
c257QXaPsfauqK/m9nfuf+YIlLvAAfHoId/u6gNcVyxPP9qoiJDuKxWUzNTIED2E
4qLPwXxC5u+gBsW2I+nlAPA0SjjRud/hVq3JqqrDdCMLsj53XS3yklT78zOky84U
R/aXUnspsXOwFrz6sqiZKY/0n/yffDaot2ztnPofpRPTiICMoPh4EHuSBLnNANeQ
fbS1r/Cb9eu6kXjp9IKKBt07aAVnPnDGEo3mcJ81TWwptALmH3Glk9nGMZne2q/3
xXwELSRzrxXOmf3+zGY/KEkw7RrisB0ue5mxNIaEEZB5v52lR4jkSIq+tvEvt5JD
brf8l8Uomt7ow3DG+FEm3vpPdUFG9WJ65CqjyTmxWdqzvRemAfsWijQLbGLtKqcs
paGyUVlM+h1ER0tmLsRTNq85XzbahUsS+jUYdjw9Wk4yOSnNwfuczU5CowAIYK5c
6oU83+4n26MXG+L7zYzl15RDLDUbz6k0A6L++LuBzWRTFEKzLAxLyqFah/Q3LxsX
M+Tup7cYprSKN5o7nOiLFhvBosrQ7gppCXWWIrYizTcMVvWggHisoMXH/iRP5wsR
O0Eu/WbvZitHG9rQ+ETJtpfutSThdpNs5S0fSeNiWzJ6mq5NN3U7qTvgwaz0nbtC
fI6fA1Gwy7w+ikVeVbDoehmz2QhJit5BApYkgX/eryNzn8XFMnTnZFpU8yfOM3J7
5oYJUWDTMlCgML7auj/8+C3q7va0/AcRUjGaxpcvx9uiVXNbd1yRFBOjcI60K6Hi
CP6e/mnMd7/L/0jZxDU0pWRANet0MKiGiuK5/vlVXlXSXmE52AvrTfsl8kzswTTR
OVDboj/q2WoZzpK6QZIdyKLIkl/toQG209dD+PadCgv19PbXC4KPmIyPnjgMOdOq
bmrRMbttlY6oaKin1TemgrHTX99Z8BIrfuDqHlibdf6ezMvpm3/X+F0l5GXDiF/k
8GhxU3yc3LT3vIPZucGMFKsQPITBtFfNZpMYoNVQkaARXNyDdlizfykaSBW37tVb
h38+OvozGs5WeKXJQsuB4janRqyiKK4cjrUWbvC9NbV7PeM1UmKGWsCHmnhJq5ER
Gq7P3dxQbhM43dv05V0CmdsMMV6Rqp9v03G3BRllPfuJHR/L885UsFFAxLsi5KkA
Gqu/UtRfVO5JrZEv4O3ITnRDM+CGeEdIjQPEesYo1YvcpRrj9SmjKGCIpzCJd51f
9bWtjw7FQtOZqmsxgiSm7HvKW2Krs/3x6Y5nEMvSFaEbSKn3WSh5axIotNY+g8XO
Q1Yon3SMSXX5XiiepMBixesrdRes/WikuwCLgrTcijKG2IuPfZmZ3rZFjuiT1to9
LHPHqAkB5Xxwn7ErOFe3S3N7o65mjfNdzDv3LVg7Nwsu+3WVKtEWs4nL5LzaPXbP
jX5dAG4rgOagO3u36G1w+4qwt7W/BPejdvCzOqbYPK+Czp0eymI/PS4KhxGCcw2r
4rtl8rqjixgGMoEp/Ys0U42QNdXI9GNwQqXMyws47pFZoAyDbLDfnXPW9CNhVBMC
K5Z/L8nJbMq3JXTinsxEQgB1CJ5OqaaGdD1sl/Xr6ngowRWgn3RpwwSMlmA3b9Mh
Db8ewARL2aoOqiz2jXpNkHme9WxcwrrgwoETlNVzbvmOhTXU8781uAQdZhGFrV8N
7vQi289GI/ZjhpM6xNXyd1XBW6OnpP+F8ytfdTjJt3cCsYf3o82WsTgHvVAY70b9
H8J/Qi6x2MUAbvsFQulIRvredbKEpE2yH43S5EMILf2kBrXl3PGVoMntr5lU9dHi
PHH7PDoCJzsLWGyEfbFL+gK8l4ZzZuBX0TZXyQbUp6Zr5eDXlMjAuceO5lpqtXod
Tvhi5PAP15237o7WY2iAtjsb1A0rt8jmO6MzjoPPdl7MFfqGCi6BDONVEzXYzorm
15pmqhaajZmDtlpKZ6C0EY2jnQXJnN5AKMU9bHWWurJFWVkzoSW9nYglb36JaZAY
f5JSMWPyE3XTPCvVu48mE3laZEuxIHNba3EyBNpz3IrrCMTOGpiWDJFX3M5YWd4K
m0nV8wPQ0EJq4o4rrSkpJuExR+Rjuxk7WweSocxVNG6rd6W+M/2ca0w5TnV7TNlY
krvrNe/jbK3GA/qcejBDyQRbPrTJQ5bVDE72TrgO4XgiZiRd0SYbqf5ncLrz8OVw
8s8CxM2IU0EVbPyo3LeObGqHpRYIv5mH++TPy08kZmC932JwX1S3BuUspARGFCX2
fZue/EmIdOY2XFpCpnD5k0ML2PxfSgOtREeEfIVku7NzHaZuCLK9/OG7LgxyUpJy
3sTln8Xnbc/4SQjaWkOg4MicEGYPo2Jo4ZahEPAzFS2ez6Rdqo5RaosiWvXehlJj
fYRhm9PTqn2RAdxAPfQzT/7ApbGpUj0m2R7W/y8FHi3l6PuIbr8GnPQPe5QgNqaY
tSTEVUlrHpAyeYdQgsZ+n8BJ0fzyunObBCvh3CJxGrkTN9kW0B3wpFVYRPGlCA/B
mYXV7YFYFJm3+DzaF2lrvYTbNHGhXtmkNIn3sZiZaoBUQvYU7Py+t0JaMggXyajF
s6WqNKO4Zjy8bd7XpPvbuAX68cHp8tq5PJAHJ6BkG05zq8SHbF3dNuhUA59gCdHB
ZBb5eoR7Ol1AGZ6msmCvUpbWKHR2YYs1vJ2G6ZsMmmcytaTn2lhyDmgmivsuzF+2
OvGv3XsVKZRNMAtWkfxnWI5hFcpTe8/xpsLW9+v8a0P5LjVQL3oceDByUwtLhAOO
lzZiXtptAtFb3fl9fbbC0XEas7VECMjOH5XO1jggWFeq1yHdnEDVNH47r6CqM/LV
6aqM2423ZBAo1iRas23HyeeKUADPte3OMj2wBTCFTr65LaGuoKp7aCqDqj9qGdqa
NHNtIH3eN6hrWu6kb2AAH5EHQZUSWtcPe6tl+yeYJ6npHNngvuFjFMZj5nrhCDm+
kyoqDRb+nZmZnKQkD3qpYortSLw27J44SjEdgemeI7m+ipSz6EdX+yrQ4/3OL2CA
uKGF8Dthn7QaCqpbhN3XvQUTAv17u4hGb27982iRFhT16HMQlq+tOxhstNTG6F7v
JTjbgJlCnVyd16vGTqlYaiwp5vkzwesVXHZTshZGJbErH9V/knWaI0no6MiWhT9o
5h3JluXwMHtnoRuBTfRXiyAt11A5xgaJJTDla6bmmIM7FH7Qd5TfkdD2QW824fCJ
FggQTsTJfaJpb2Y4n3HTbKPz29psm2m6aM1CSwSXpe/qjLv0aJwLQs+r0tj7m7qn
zNON6y4fwiY73g1uoXXEHwGezagFwvY/tSQJrM2PcXwcN3/7dGWu3qvNAmUbo4qU
qcfVUwCcaCt9cYnu22uaw8i0q7S7wt6fTP8LfBvVx82dSND65lOB6ISkhixo3u8G
lW9aYXFdBZjVMTw7hOpaUO7lG2KlX0nb+cD1i2zDbeSiY/zRWo1AQvL+ddWuxi5W
GUEwpGGvVUvYrEJm/0GreEsYAc3KhKcoCoe9myuFvXzKBVEwNWM5FbiZBrQpUn7B
6Krxv2LD9afFXTWuzQA+f6KV4oMnhSNNJ4uUJT3ahL4QCWb/CrEnSkbZ2pNA6yri
9DwTrMcC5dK/JlS7atBb9NbHVsE/3fqRTaPnchJkUH2sQI8iOy6IyF74Za9Zbh56
p0VDnDc0OMXruN/gsTVm9zrrw/UYsZpWzqoNjPGjtRcjuu/mnqxUz/VvuyBUdVXk
TTHYoGz4DwQcMjJmkrg88Es8NHMj37F8EcJxUAH5zdI3wTlO6yGclEIx4HWn/x53
D3WtTAxBUCr+kUqDxhsgCeDvLzdB79IVo7ENOEgxt0Pxz/qK3wNYGYDI0PWRTx2D
6UUkvBijw1jDGJVaHHByQj0ATGgIgOesWIA0D7Oht2Pnst38ph1Ztr9B/UD/gtUt
PqlKarDZGzmKqS31ENEFS8e74rN28H8PEDZNumO1GDlv0U0YFvAWrEH7SMyHLHhZ
ylBxYG5yASQvhqdQbH4AMa7dTfsKbG1AWyav0gGt0dFHYoI+Bq/Cy6vMOVYE3+Ev
tu0Lw+ZjR8rpEPpzyA5xldNPVhEv3v6qrWq949pxPst8wtcG/Lzbc8Nqaase/Kxx
ZFQjoD//0Y3PZn8Ux3zr+IO/w0nyTZEy2jd0XpfYMWSxkq39m6p4s9fZQ95oZcMQ
lujBlm7JorE+KP5um3/FQlsLkH+7JXPjOoHrY+iijwyRB+BXz8po5tVpX1OR7vn+
ErS4manm6YZdg0yf6KV3Nx0Q+WsdHkCeIdy6fdICcT1mx4A55vTVrWjvoyeSAeUC
KsDBe6wEglovpAciyyKS/rSS0LT+Q6EIRrPd1pPybBDi/ZDHDrNIgXWSUTtKckZ4
gPwYkrxp/w1V+VXaqWUTyqDnZVxh0tU/o5AXIqwOGwO19iUoqIwPaZPqya817JzI
UvvdyirQzUW5Ouq8NsadeLqZpf84tzi7js6ncLZYvOjOxQGn/wSMzBzdBBTXL0Pt
xURhcq3HQDvHu+Vla/9y2lrClc+BIVlo3LLiExrfj8Kk6WPm/uGsBfdL50DfBDvh
YwBSvxw7WtOXBZK1UKc9Vyt97+NVFGeDIFS2CponSiTclfOyqskh1UKoBhXzEpXp
uPeXtdBi6y1foKDNQ58a+q/P5AAAMlgcrx8gfmePPAT5HlRf++/+QGJUBEDjQaa/
FbvNhU874KNiE5kz5BH2wbKws5WEBbKJ3Jsa10F/8tcpmxijJyHWaz2MiSV8Uvk7
bs7kcAofGbKP/k1mx334NbGxUOfeBmpC5w/23p0Lnr4HpVpGfDTVmcUP8DbILpOK
k7qsfZEAhrS3zbasjD40RB14wD7vGZVr0Rig97nj2uHeAt7ZcqG6RAntKNOjEfZU
1nngj07UwlS6USXIRp0nMQ4gGb/vvYrOV3PQwQFav1BqDev8Qd7CTOmuutpder5M
nyKW+iYe2lp9hUKRbL07yAVm1+iJWOMy+7xA/OueSntGQDSUMVBFUC5Ppohpe8al
/p54vLqVonIBlEz2zYgBR60qWjdzZr3mqGDJdWL9NzapSb95O6zq3YY9qHCwkpe0
i+Zm3dQP//xqTMaGDU2HcuEqiqZtoaM00c3EJBKJftr91hGoUblKnPRrqyPqT/sI
DPBglfJTSop1lKxMOIMpziGQYHM4k3As6UXr+pF2auvX5oLU4rUNsbB+w1VviAQw
uFH01tt3PxfmabWxlhw3SZNzBLwy6sgt6qHupA+RPh4soEMBCvDZNunfF12nE3UI
Q9bIDwlba3acC8p7TGAlE1BWrhFVHCWaAK4We1tI5sI0hI4sCEUicMV2z9hQMOJ1
bAGa+enlf4t+ufFqqaPsW5es9+Kv8j2C/D8RnTNDqsA6mCgYfIbE1TZ5rWbciBsd
YtyH64VgFdr3epfTUfhPQmLCGJztsQyh0KgeN03nq29ZfMgJVCYQkMUOoVOEPZsh
0yw/uK9cQqaT0RpLMgyewj92WL1uUI/CDeMGddjDGAhcHBOK8ifDjiRAw3tERzxt
euj11Gi+G+Yf90rB6bH3gDSpTHB648izz0NSlaaYKKmdCZxejsit38VZOyJ4G/Kp
WBnT2EgVmNPJP5AQ62buEg3OD0IFE8P1I0ga6zuhxG3q9C4aX4yb4s8YvOkRd21R
oz1lO0xdonaCD82opblTOUzhN3KMgXuJuQV68eiD1xJSU/7XgUmdZXrd3IBDtEwN
7zFCiXQqdQ9Tcn4YVognCTIvz8OF1vgsRJTpudL6biqVHxXN8hwhm6R/qs0ty6q8
MKXrs5dP+Ly0D3EDXrWLWAGHRNpF/uSip6PpV9qWYKqIuYf9IzVNzW3x0celxHTI
wkDZ0HOhDJVDfYVTSHVerqL+4S/69qSPl1P1jwZbupNkZO1xYZiim04rJuHYiglV
63kV27XDsxKPGbPoBs0jYnOxkfzlJGgx7wFkGmZqrnTp179Dez4PgyehmpH4eY9g
VRtT51bN7m5kd5VTdoJhLSCPF320juyRKquiI/UwWTqvp8z+XaT1m2NQWZTiFE7F
dH2JcixEbH5JpTWKaIC/wKTas1+DVDTcTbJspz5DomRw+A7+x0vE7QkeU6HzWiSU
FqPlC0/Lv9fG0JritBrsqK1tSRySVoCIoEE2ez8y+0FzDkAuLLYK3U55pqub2TbW
W6DNxbwEwFScIQVnDAKelWr9baRQqwze9dfuNIYnHw3lk2yleuejoeSgdQ/zNg9/
Q/dFFVRgMvc7Z2k7hPak2Pl99mru/u1eursoyNsYza9EeHWbepdvN/7ifIr7S1XF
0zOZHcmUw4XaMUlCtKJ8XiNByQM4GYgszr+EhD+SSaW/U+3nbzfdz3wyzgf9iPx3
pEDiBHRtIVYPc+w+Rx32K5AR2nrLqKPxAe9fZiEtZAjTVYpsnCvBfTAG66gkDFN0
eqOXvgHft5YfZZSCjd1TjA==
`pragma protect end_protected
