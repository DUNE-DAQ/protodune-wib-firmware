// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
akuqUFq/mCIY3bpOGF2+uMegOfxKE+ELQc/X3WSzed13OeaSOwFhXJCx7ObZyvkG
I2T7fufww91x24LfnjmRloYIrRbioonKGDIyMVFQm9NOocmJcRsI8c3SQVyDKUZ+
eilaW7YlttvcPNvGtQt0jBjjNWIXRQ4LyOAXDz28ebI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18000)
ae0am3mRv9VgzeEUEJBXdpiSQBQd+CSEvksPKaAczpoOqGGeG745sVu7TVvqqGq5
HICRmV543jB9FmKtjetSGoTq0sGeHeL/1pIXOJAzdGRvPtbk/REmT75DfLuTjDVN
FPB2KeMMP8qHcBVJdrpt2B3dsPcD8FjrO35rsznUbGQP4bi2zAC2GRok0f5y8Caj
VMEpWoMkeol2V/+KucLI3NJGAbbpB4YmOYqK8ADtLopntw9JHBBY44Hk8ZXunNqS
cgakYe38vy9qVrp/a4vjGLUVieomEzobfKxDPxmtQsRkGcC+ZPnk6A1M5sOGblXq
b4W2Svjum/1hcmznP5MppEbql8RpX/y8bxHD4zsuZwiqmeF3ingmCkg9EQy5/HFw
koZNN5BeGWd1/TXuRo3xt0RqP7XYJz1Juoh37GqLba+yYy27xIv8QzQ8sm2oZlu+
0E2TtyidXvmAJSSx3LSZWBKL33OjomMmNbW7gBM3QUQqp9w7QFj7W5CstGgQGo2k
CAKwbmyQkMapJtkGGjgrlkRvTOc06TAtC53u6Pt7wpNkZMWMavTXYqZXwgwKWS99
5K8C735YBO1V0WYjxlcGeeVyhaBg3ZQtKpQ18DvbkmqpGJS1t1gJITQdeChi96ck
XDs0NyGrXmGVvZoAIQQfXM46KZwYpmY/h8YPAD1HEGy3T17/PhCr6WoFkJivXN1B
q08+R6HwAtLoU39G38fovC7L2Yn7FwGp9lpPLU6t0YC2dxRnd87Bnv2hTwWSFbR+
+/GPH8nN6lBtWdIfoJG/1dFO86bi6MkUno8T9s+gitb7QekleH81nukl4aF3SFQz
A1hs7CXMolQHrp+ZtoGLUYxKVsiRy1DpYaUqIrGjIuI7U2IZ8Iky7ofYaW7fTKPk
cKNTZESHQyiDovgBFvRfmhHwJM834eR89fyR3S64XXi1hYxbz3eWgwsVGrG936VO
FBRVCLuJm4FGMsTOPBIon1SuJlDUZohuUeJvTPlMKOe72DwpOH/5d0WDTI8djxV2
Rz83bnsK0BUZt6yinbBYfWH7NX2qrDdkzIhcMRnRdObtLdXF4b0C4daS3aGk299R
2H7RisLjt1JhLBvIq4zZ8HtvAUogld4KIQaAAgrz1DvD3nUtwBH0fdD2V8/XFV3J
guIUtyBGlJReqTDYd/QU5LgXcTbOvCuWI/PwBBruscJ1MUopaiHeymUPO66B6HBV
X6ShoDKsuVCOJDJ1vpgyithECe5KeO7rTEDudCeFDfdKEcgh80lCMirX45OjSUUT
nACTpRkyl1297Xm8tEnIIZ5gavCAI6r4iHC6tIwH53JqnWPc4Qn9f4oxMgScZEKz
mhPOmlX8YqKzAp80cAhPdSnOSn5kEIAHexiLghjGHIV9HoKQzAKq15QX+qPXlPX/
tTw1oF1Pim8LmR2Pok8ps1lzwqOmo8WfCnsuhPtZQctSK7KkTBQhch+uUeLUERB/
XkSMxdRFW7N3J6JzeiOxIU8gFtnHdHkXkcojOrhXzmZ2FCVjLWj+JwH9WPEXYNmf
kHDrXOTOLrAscCd7gwwTOFAWCWO/xFpNJyIK3U6olWbgWbzMqMEuc8jfZNhfhDBd
RCrmnEMghW2jihNav49/LZRX4FBLLvqtJQauWTyugrASDF7ncPGktdXhVBB3hIdv
knE2sCNNJHinVWOi26VtN4pZUjSmWGJRSVpJeyWZAUqRH4TysISAvH/xRDA1j702
hFKbjghIXP5QtSS7BexrX3oiWDZAT8zj7vDC7qrM5WDSlmPARaqCsf7sHX7s3ZFt
Kzp7RzGa2Ae/TccYcVrOATgA3GsLGXulUim4PE6gLhGXKKkClDRHFZ4SpUvKea0J
KrVFNGVZuQ5siz92iVVl5QO8aZgohQlpngyRtL4nD3b8ywH0roCV9N+Hl4oP04PC
mnXqGTOkTUKox8tbarWiIHPh5F05qZfulCb+Pz1PYdz06BFm0iFt8jm2XSFA8x6r
CDl6LEOtnqZnDs6KVjVo9TjNcBHpfjJHhKIKi483zcJ6Zsvk8OPfirqVpu01qbha
WIS7M0drfgFNmHAMjp5pMfTa9O91mk0wX33lQCi6q05S88QwZpJQdQHIzjBSv0ro
xYCnPuKNyaO+Esu1fyN09V+4PZ7luQqZYdsteNCPu9Z6TxePa0KvesZMxiIk9xJZ
LQkAfvrrBLHbVs6rH4hoA+mmKvJ8zetShSgSi1u9GbgRvOdIVTSygmBIUjUO8oFg
6MQgXomcYw1XYGIx6E4jBMaenH1wVD9o3IFCReTPfK1lj5DqvmMimy0ZFS5XBCKc
b62FdcjYq52lBwoXVBVvwALu2c23oce0YUkI0ahviFomtC0cbmDPzJUHoqzyRTHT
UhphjQ0z5QogOfQe0XI1nvYvOljL5Vgk/ycY5dgg3Fd8l5zJ2D/YIzZ3hvBD4vFA
vMy1SKe/iFoxviZL11cVIkTa0+3SXN8MQUZahLXDxV/uijTKgjHCwWyKXmhWwnUU
3CCQcq9Zv/0lEbcP3qMCZieStYHYqXg16LorgrWSkM2waXVzxJ/7woz3XSE4sJ5g
J4S8kZxRpbh7SkIuJZd4qq4ke0mEgR+UlQ7MjtDVFUYmPJYhVy0TMOd6SucfiJ8z
8aEj9lgGO/0wtQpyF2X0uTYu1KIKHEevm870GPudAW9Z77FMx+rvdemCCCY2FsYd
nnnvOml8um8gRkirBYfrJ26i8vuzmlJe+qJK7FJ2j/AtMSgl/KqHFrwUzkB43Bzn
61hZnSOXBF/3AVGomKBPHftNTljiYRxL0SpEydNSHpX4lxJ64NjYB5YyYt1C7tpW
nnBMglQ+GSXgbXS8z4w6YssVgO/t4sELNgU+lHeHtG0lcipvZxtdXwXlXOMmsGlM
UBwkPjAEGnXno8JzHwA5jpvuFNNSjQzobrcgATSMGLYi/xBGUodtvrmJPFIY9q8u
ypNGoj3EjIqkQ3xSAJ52fHTU7Wzrsam1IOgqeImnAySRvfM9kS0crQL22fdwNxzI
XcUhZS3R530oUjANd4ki94/4LHi6PIHiZmCEIIrWFe1x6eJaddzHu7wffXLDBeLn
0mGf5t3LqSWUBqzakEay9Z1qyZx8HFcE/0ucXinJ05K7CIB6K6Juvs1QuwuX3al6
HLYwZf18Iq34zyKNYRzO9Q5mz+w4uxZKtEriDhHgjCyBpUX4kqMPy4GM5VEFFeFz
9my3mu6/kg4qPwmvCetoYm9ID/P0IN3WMu0bu29WdoOBNh1EGG1JAtrFTYMa8wdT
wuEiVizYtr1g7r/VL6/y1rRU5ooLjCT19HyBRWIWxVuQIzn1nWhhhqXfMoh8LqTm
mbLcU8ibh49wp7b5zqtPo3H2mSjibn0sSIA1U0WCNx1PCy6AfaU4/SMEm0ns++Tk
AC1lT2CdOeL0znXB3QJxisDGkuEsWET+4bOsbXk2XE4UYvM0ezvz3YN+diQ1jPYX
AE+dEvWFroDEjPJe9rVWFgB7LHzv3yOwHzUArAzK4aLSZ9aUvW0Cf3Xf+MuXryQB
CIKWm0krOpLHTCNUP3Dcq4cD09xfkNI25qZydniwDRqkg6cgkQSlROt5XxeaioFk
DgECAeO5B3PDzrEogkNU7LrHzkNm2Mb+5aIyQ9kyiywfI61A+kI0WbDBE8Fkud7K
RpgkVYNi5R+SuCv8bWZ++hxHd6RlVel34eJ9KzWGtDtLMBwp0fKMYQmeJS+2QHFa
cMyzAQlq8ZxzKhsCPoKdpD6ayr2oNq2c5wnToVlVlXNDuUXTCpF/bw66ako38Fwj
QnL9NOvRYKCt+dVLaeqw3gxyMkyW9Y6fyIcbX5tSV6lNpsgejXexRJAiSaMOR7Ip
61z2s/L+nfdP8RUGG1sRqKzw9CZpZFyaOqK2jTm6rcysOE9wLMIWwh/xOdES4A/C
liMBcYs0DtUmk5AuOeEtJ/wsPQdTUvXiZRnZIVRh7qIS8+9RWvYFh00OEqk89VKV
ZMGB2uHOgXloxSg0EmublESu6FmSbIo4ujpXZUUs/WcZlhmivTSbHgkT87oi9kUs
5EisJbiPmhWDao9P7fNcBvxJ/lmtTOQhT09uI6f2cOUkqOZDejcjXAVCALq95YEi
9SIjuFecoYCWfw8TiViWemj71vAxA5gdz75AeRigMIGK54QCGQq+sscxVzlo3hvo
3NkmitcYGQzk8frQeKbF0JqcVAuYTbGuIPQNrp5huKFUs1aLWEJd7NZrK8fcJRYx
V69ywckvCBlGdtplfmijc8vTW9kv8JD86chCLMW5jpYR3ZfNYVemCeLNl4NMng82
bvzKD6jjyycwoIizruCFnMgDzedhUm5IbK7ep13NpCFk+vpiG3eiQIMO5uAX2y5x
h/VuxwmAxZBsveCppnhJT+5ri1vfDGNcCntUGp0OGXbqg7JbR27Dg03RDEa6F3OQ
XuSus6aH6ZoL2kWFimkcrjkpPH1SlrFn+VPWnYOQT60G+ADbZ+OjU4dbUl+P3yam
TpB4DAKbILlOw0PqKHTE7L1p9liTCySnyOtaNAf7BHPRfaPaXFbQUhTo+qcY5sIy
kgsofQS/vzVBspaL1+F7qJCM4fFxI+m91/xUB7SjOfibH/k2LziIzp3R5/BjU9CC
a/6zUq2QHCOg/Tqc2svR2PpT0RzGOzVPr6gwpGodbrxL12Fn1ngoqkJ2mnF5wY4d
6MVFddX6E1dtJjYiKqg3hBioLUeqgFri7WL1VBsHjKTtCpVEy4eM2UzP23jEDCfI
Z/LBqyoHF1cNwJTg9p8SUjfuCHlLmYNqHRjwLJ5hNZ52ZBfnirinwLZk+GaDpaJI
byesywK2FpDlGhdMsY5s1Mut7QRnbPA4aDMFCNsiaxswt1op8t1WTY+5e7yzwVI5
P2E+frRxKhyzITG1q3Qme5Cu1NftDy+1WqXLi/eDP7RRtdD5lEwaJoCYWi6XMETu
NZ1KKd1xVYF9gV5TlbggPY0siVNAnlIqLv1u/Q6FRprmXYtr3JjftqzkdmtIYRk2
0qSJmQubfPJc2VEQTQja5JpgS/ymCJQojjei1g5ZxizEETr7teSzuA1VCvhcbWA4
3Zze95oDt9Uiyv+rvlA3sZoWk2fJ6qbOJXP7AgREvgMlgWWvTSkeyvs8/zPfu31K
m/D9J11qJAJdbEOHWsKtCwxoBLLc+Jc2nbvHA0yCaIPTf6GpMtoI59lUuIcnJtEs
flN6yuW3AW94KT2gooDqr4QhZHVR2RS7PlOozl7F91fEOV+YB9lxrD3RwT3x5ZWi
DcRnEXM0q5BrGRNoCBOjfvGCCHOJMAjmIuzh9rAyRVLTqpInJ1JBhBy5oJE098H5
RugnrX6WiUOeW0ZhBQUZfExqzQaEkMG4H4HcjbC0rEOQy35dPhvQwdBqVWii+XVe
YL3IRHAuyPOv8E+9wNdXkCZpUKibuRdcANmnsgN8XhDycAgNxWnQsKtG3neGaXqH
2N5wru6fUjbmSIXPGbadIBcjlOwk7FOpyOnPoyYuKfuCt1eTPIFUawFQT6cfk1lO
fgILYN5cVz3XsTj3T8rH+iQer37Ye5rIlKmv+8DxX2N5+5qrpjgL3thw4myNAJrV
9LJGvqa17yL5xRNK/at/5cBthHcuptio8sHxz48UCzquVsU2amd4uofghF93whs9
qwYA7b/D80fW0wZolMPVTUgi7Kc7Q2vZu2+ghtwmNeT4+n7RcDD7s/JUWSTtKpq2
BClhxMJ3EdCqmYwXbnFieyFISfjLqWXlxqAhJHjUYgMtpGaqjmToQ0tKNR4cM9Hc
8/8VR3JaDQVpUFDu5pH0bQXM9NSfbv6RUwWGOzCylA+7VkZWNjqFKSbqy1OpmAGW
89zPuIRf7mryxYGrXiPmhw3KYzM+n4CKB0bPtl31SDWVeN0NSrb5Gpp6IdqIXCLD
Xp2A7cDBTvLs9o6yP1fKmDchvDFjYcge1dHYBrQQaiWgDkWPhrRAo0NFyQcD2v3d
Vt6EouF8Vnve0dYxKW0yHAHGfBunq3NMrKT4M2209LoOuxg78dQrTqZOl8t1Ymgi
vagx/dVwk2SZGLf8bxejcvfpTXGdAxdAwpAa825uj7TMYobMLuqdyxxHu4cOpaKP
ekOuokN1uousArnKqCxKITGRMAL0SaLCcDLx1hfvLHFgLvOgYLZN6ZI84r7d+0DN
Tbx3Ie+jBKgURhcBHyrF8pTxy8D8P1SuvUvMNtstg0rUZ2g/k1s1on/+epQ0OsgG
Hvg3d0+63xCRb6OJdmxXEtPR7AfLfEhwcRl9uoIEmcPu6w7TsY9QNwiHUbPNrUWy
rdz5ItqXQ8cp9YuGzE8Kr+QIFKFbDl8fe5W9Djkszl9n/2xqcbj/swKiIC+bVElQ
uE73nT0nlw4ye08XmHkwM+m5Z+m/EBWsLPYkP7yNhkjCg79x2He7pzlWsb+fstGl
JaZSDTHaWLx6nQyGNITD1vzkTng3wBKOa8IHssd+FFuU25F461/I/OONBlAN09IL
yy4o3LJYLvBRSuTg0Szs27Egn7PE6/JNmMK1uNEhWibP82B03rUm88Ueq/Fc5eQQ
izm6p+t4iQEwnQEAkFx6+5/LC6CHffwJoD0iC4pest2NQyRokGPAypeNYovfWAlC
jWzsLnXQ22Ws0ieVNNJgF9E/9Bku7jAW5zL2Cpp4DhrsETeiAh3rd9FcpLXOvSDt
mABaWIc074vgwu30rouGjleW/jpUq2alOqncwVHdp70cGVw9we8CZc0K0ap3hxsA
KTvFGiPgKDwtXh4NN9cRAFqKQA1L37kmuR+cYElUGUsjmUQhDs03casoMpj0UEpG
xgSF75eqz8QOvYSjj9yrHc/cfK1tFU0bDm7x+XS1eGwLIhQ7Ln8DJeDR2iXEfZgG
kB3f+38bUDe9a+zJNl+Iwco2IPyo7rKqAPh4hMjQ/rGS2z+2eC5WnQVUPvpfXUfd
aW1DndCQuj1MwjWEC0iE+PdK12ByhqIBsUJ7kdvFeTvuKnXwIs0SFKXCwaF4OeBy
x87qESwKae5uS02yjdWS2l66zWLmqoQoBtiIb1wfQa1oPOtInwXqRnGcg0Hi223z
zClkRoWbtjloboobU27OfGhvjZIoiqz5oShKlqgjHO9UFMwSEv6yluB4YOhZSWZB
FjxJq42iB3bHRhLLRMQESWmy9nfmrZgYwVCiUnwx9qoUnSL+wpTMOk9WVUnIS8mx
MWobWHixNmLWmKYqla4IZFEqwB8d1zv0sKA47uKwGeXnuxkSIDCSerP77AoPl35v
MgPDlrUXhC4qDrePKkVldH0QcOJOYgrSIo/YodXZcaoFyHuBvHkDs5QAOfMpcTOQ
yLYrt0FN2M8HWh0D66dNWkdJKfZKys52U4l7zuNg/4HF6TlPrpFlH7oPg7Jdhhrr
7/InxCUurYS50NioEMZLmmDjMKFCJ6RmDcQ6zc8WSBJ3pZtLqcHDBgochXKVOJCo
q2M4ccQNhZqmEx50Hh4g51k5vAgTNvXzPvtnee105mAWFotST6va2v4J/8dlO1aK
a20P7tzlkpYYT2tzlwOiHCAidqhJrzj4zo2KM3Byh4IT0MoicqoXDy8x4ijiayuV
dDlrPg4KsT3Wpw2ORQ8o9MBs57SfGzf+5NKAVHzxjZ7Vf/76tmK4jg2YwoyjKVub
2Elmav7Nf35VeSUX6d98ckp1HE1VFSk8B9WOTm1KuV4J7+GEL04wyCVElOrzGakS
0KbrO7PetWDRrZJQoBDM0K9zkhGM0lJo4VIAxtJC9128uhK3VS1h5rcOqd68oCsX
G8/6c2hKJDVDT3yUqZJ/OOQhRgZZCihtpBoxoOoAzsAjIh3rsVx0Ah8KqjJwmPh3
k0XVihlnz8PtP7AOH9eTwJM64vDttEB93pz0K6NBLVL6NTHfXkQRmzwsBMR4e/hm
Y5OYQDdbIEFY8FTxJpaFsxMT75rMmgvXVj40Zf73xk/V/6EoacTsd9PV7JALwbLE
3b1U+y+3jCp04Oy0teP+VmiA/fsq5khXKWANiMCWuECscsvWd+P3vAzvYYA8islH
xRCDoXbvrDSoTvGz0sVhXAyrOl5Tp2i5wucDlEl0ibMRA6VrhMyVsTHRGVd4N1vf
r2ahEik/yDC9PTIaxL/t7Nlkb7LM2xVz97hKI7uxtotyzYPhycdu1CPJhY/peb/m
RP4EUCWZt6rK+EUz518VxTA/ijkrGtX6HYG1BUSKHuDc6LCuT1VfJv3eJRYEI8YY
8ID8b/exxXZz4a7q9jIYVIA58r1qoI68VHFzrGEvvAcOOseC4pY4OLEB6X3mkxa6
iwDnp+CkRAaIrFC67Q8nYzKStiyJASbVxndFYIQDo+EgOYe2QKRa2fqpEET/MPIi
MUeDqQVdwdI/Y2Vr3LnUi3Ny5/ZVRvlgJNlU9Vp6JZx5eW845W8p59G8pCAciN++
+5QT7ljGr3Sq6N11VKIrQ688UojzpMb2qmJocEk/cSw2G9R6x++jSbhV3wl8QXrj
CFmloHcY7Dn9A2zmFrxsquKAfUUx8YXmJNH4Fi7MqXLrHMqh9/C0Wm5MbnSkvXOr
+5yLnBYwQCHTL9wjs0VQEOxQctJUgRS9VlDpRHzmgqWt1jpKnfRGdrjwVjGCEIA9
noTdGc6VSddlTEJMlWGus/olMywrXHnCkVitxb9v2Ml8QbstgLG9WK2Ws9JMvpX8
trXpihFOhQ5SgnC66kRhMPaxlYapmfEqROgaTdYDD1od/smXdEWAbbsP+YxWqBHg
85VTWTsRowNN0Azil31+mcsoTY/nac+bV1j3GPN/DZdzvPNc+dGMw41kc1jPUQSt
cPw0G3qJcIn9/6eeGawu9x3Nf0tYBmTIt+k6E8kn8CsyNDFjNVJx19AtSUlBCHl0
h629mm0xv6+GPWel3wWqjiNbNEZKpkS8tXC6L4H0qjL/VtdbLq/IDYcE7rzJp5DS
1DCxd25imV+5G7JxmNBLJNPldzitNnizpvkL1VOE8V8r25KP/Pmk0+a6r5w6UWfI
KoD6h7hQNSO9vUDEYaee3wRZY6QQJ4yiUeMb1VRLu8pN2cb9QNjEiBAOCXWiRDXo
iaSRtBP6CgcMgUFAMIh79P0wInIWfSFbjCFlDX87dTv6JXjeKKGeAowu3H8QPppr
p2ypsFqQD+tpyshDQ1wLVE9zkuF9UEUhua+OnjEoJYlJNhclzSW2PhHkkLO1MDrl
s0vPQdgJRKOD0qhMkQTvJbRvQDYwDF5lbOTHgDrHeGP8tkiifHov/K1bDLS6FYlu
uBqfkY+A7uXDgj7we0Q3ddV8osSCG4Ls/qdCoXYrgJyoq3xKkeqdZJDpuxQSHx0M
DLGOWaSZGmXwjbvFQlIaesAdgngtU3L7s/nYVmUB30Jz+8au7KWwcbswWfufVbIl
/zN5CeU6OJcTyjyFeO22ILp9AuEjRyMyXnaORlYVPLJjm7PygFeQhCI6mpJ8rtci
OIGO9/71bqTqjmEanX0uZG322sS7zYV6aqOt3fjSeD0PRoNAB5+/kMPbm9WKFh+J
HJGjyP2o13xEx7YGx07G2r9/lbQNfuQkq0bGLgBCsCFZIpcx86P8Q5YuRCNhu9K6
hIy6zJZcK+DpVoSZWJZEcMEPsYamN/l9NDa1y/lS6ZA8pEGnARXeOd9X3ZpGFKg3
k50cOelQW/o1K5hTof/lmW1mIYXxJqlKNfxfyZ4Zn+UJTQ9L/wqpoQANaxYbJAV+
xzNB8ZRijQ2vli8Xvxuh0ZJs5Xrhz5//hYLNUf+bXgDd2G5co+6hjsEeh2UZqqCc
6PW/3YyX6D44Fy8WbBsbFotwbttKVjfl+nTb3/6Won9OS+WiwJ3mIpW0soei1gL2
u8mC+osVls51ft0ohwnMuXMDsZbdgpJnyjZ5WYYP+p82FjKHi9L5GZ6AyKOc+YqK
wgP0sx0oxfLnfxDvecmZ77qm98BiF3n897xJmbqgErusJjNHASwhB/XhLc3TR5iJ
C8sU9uTRb7YPjXOP8plGcUbVXhwpnvkki3G/TDsAsc1nrnXoZ3B41lAQ4fZTwdkh
P+v99eqUEU0tfwjcPrfd2YhdtloVAqIBBOvBSwPggfqu831hoj6k6TeSQU5/77Ag
8dOMvGE669NN3d9hpE28uTChYzx9Ju7lRF/pM6N8emPXSurYBndKUzPh7lAOdfHF
jLtb+q9J2/A8+FyiYeNo8TfUaqzPi6d1MmuCWWfQp2D2CCbEPzwpAokbrximHcps
TJHrioKzSMrYjTaqq1RUF1GM2zFYxzsmBkY/hTyZvraOwRTSm4HtHC50uq170S3d
UEUlAIB+wNXA9FuruAznWF4mAtAraDOKgBxAO1lQP44pjpH0cBRUXoYu53jQcNki
h0fo+4tnknV2wFONYu5Vh/cc5kgj6qdtk3G55OWJB1mtp4lducxonZY4YFqxujcm
mbl4n0D8aA7ANdAvYTSvAvu1BviLMliiHrzEHoft3++FxeobmI6swe4iXCVr6L6/
n+vcRHw6Qjh6q5z/kahMEKS3dB75RqpYAG7ujrSzsGfhXPoxPYZLCytoWdvjMdha
cER6o9U7/KhrHM0VlkxBtBcVjE8tjIwJ3xVnmJjEKfTHXqTFTgAJLPrBpv7mB5AB
R58B/9ppt+siXxy138TACzYuS9p8pK2zHfvufAAYhd8shFPsODoHwx3rMmIzlEVC
sx5nmfDu3LsxIBDzkpEoxx1R2hAYLIq8gLVM9x/6OuUruRzXXLrSqARf07M1olAp
VWM8CfU0SbBqAeK5yNGxlig21vfYs6FYi+FbZSxbhhQW1jrr85b7TYoU5A1tarNV
b2JY+3II5xUyPqKetfp+3QoQ2pdo02ZB+IX19JO7t4IsaNo3AzxsTUkqLvo0Gc1l
jNgfxVVKvZK3bFwJX9C5zRm8PQu973wHTewpznmBBC9XbHuBlHKEzestNDY/OxSQ
XlEIUxr4LhnTuOQLHkgX8bJYSjiVprvZEi42SVVw/2OoTCXgPivvepEor75cxR5M
CXbAT9NyVj3Qxv3Vjv/enibUh66sHJ7rrZBRT5Dktu27frbR/MOhAMghnWL3cuTc
i1nu4+CDf3wSPNuLaqH6GKHzA62zIzqXz2q+r6Z5rP4f9XOFrfgbQlbvameSaGsC
1O56miM9ZeXl7t5EhE5jCPCjFqBqLw/yVP4ZcSsM6wc7S2NzO8YTEvBZfc5noFLI
1jZ39HTADASHwYBPf2KS6I8bXNFW0vVtCl16t0sXX++l+aTnyJXteEKCXv66OAmJ
fmk1Yd8bIllzBnix7IBMe4rzaLTjWo7cx8p338eKWfnlJzjAIFvCFjdJxyfYnt+n
IulnpbCHxhkvM/cgu5ATPbfF9uyTqZE2kYFf/t5USVZIKHeGWHjGWq7xW/hWTGeY
+82CvNZasgYKZp5QSFcLI8+uDHZTp8LAfZ5Pe8OaYxDAFkwHOfDrL05UywXwfoOy
kF7kqJHTKtnIujMY6w82tXH6aFWQeMpcUjaiG5W1xaq0EuKBZ4KP7QnGy7BaTUqx
GxfFdpzw5v7ahdJDYbJtgdFQSPObCm/oPsp0aJtftwa1sVp5+cQw5uXbpwX9C7ks
P6ie1VPSdO5+1HjZUNoJzwsvt4JvFqK10A6ONK2dhCv6qFtKPNnL91dBpsWVuk+t
QjKiw6qKmrz0CQFYkDUq6w0p9xAHlttgnyy+qc7KmrGHH30R6GqHIHDUV2HB3M08
8knlDFD8hFTB5SdEC+p6grg+rap6P/Zhn5LqXAdAV35ghN72ta0Sd6A6+u3MVqFb
Sbh8sQpZnD4HIDFQCgp7ktLbcRjn9ZBVijozcP5RO+GRbTaAMtcnunqQOTRYZmqg
vZ6D6DHFK0kjrP8lazr++8jVWKSxHkjMfRkSR3kzMQeS3T1lRzT167XJX3c4+je6
IOl/kqiz/ESeKxbTnwoP2G7dtc8sPFqWBUDKAgH2JgeQlVHOb5a3BLSs9Us5PJTj
5I4KskGkJ/pdYeIrxNpBgVqguGx7rb/iL1Mg0OTiY6wfacCDCiKYnn64YUYDVTQq
sXW4AbfezzSXBvDR2hX5X1/gVLjm1ozi0V6ZGs0Mh0x6S9kxWldA1UmxdjYmrZXM
poXuoa1uKgiMaHqlZKcfTmU+Lj5VRknZ/gf5REE2xR6akp1aa46HSWZkrE2a3eUs
rqBBv+U146eVTaAzQ5AX6vT97P+SazS2KnVWim4+k7/kazxSHIxYrVHv12eApUjK
ii5My2du7cmbQMhE354RxBTivoEM2c3thzUG2qCNR/ROdGNB9Snr1dBWdBzfuZJZ
NejJfhhF8CEHrGBrKtH9vpxOVlRqMA+DbVdWVDjTLbrUy8MODzeazL3n57d7dIY9
q3ylJEe23B0pAr9DyxWuPk8XfKiAUGB+XZFlS+VSdSMxtZFA6lbEJe15BuGgsT4h
Njg/wa1gRxesaj6tp6OUSXAEqMQgMFjnrX7HCjLtEDqOja1KwSDs0AO5hf6GID0L
tii6YFIsZkjenLkUXpXRXwfd1HTVVt17v7crLzWNFLtbEZioq7NRcWkTv+gtarXV
mjv1BQs/2lTsgnX80DZMTrHrwYImvqA84IInrXqiOemQ92w0m26bwNsdMTKzXhyf
wK4UFFkhkMZZllSFVNulVrXrj/z2gxllOwDw0P5DonLXKhu0jl5EgX9FNd/uVjQi
S/OV4v6DXeXjoRe6OuqcFbnIWtm82ZpYDc9X1C4phjP7QgFih/6DWND5LQA3/5ZB
474oyrWJrfRsfgH46i5PPlup1n3ZZS42q0DrlHJ7G500rKrcfj+3Y4ZZAY41Z9Ba
mBTjF+DKZycQ48X4dTYHA+Tlm9KhK9S7AJJngxvg0nSqPPJt69jf2UoXSmMBjFqH
YldIdxHr3GQEDHYcozWlLBY0bjqqNd8UEfnirPvIAHJZSSpZHkuIL2fBsakVtLf/
K3oBFnxq+zvReavfE93DADMpDgJRo3eNqoaKYQm1xfkDly0D1hSouibHHmf7jMHE
mkiAYmbcEiGA5kjla+0vl66llSb80um7idV+QQYk/F5rzLF5OyV71mHAj2BxFIDt
CF/x0XXSQTvizyPzLkKuMtsHZ5JYL9qIt3HaAIC3c2W4wTLs4p8W/qZgEG5FfUuG
k4zRAS53gEwdiHxpFPaZwyS1kPYeWfEk2l1OqoOz0a5cvHrRw/WqbLdb9EFGKkWa
/DPMkCWGYH+rV+hh8M6a7Wts4JLAG2BEidtucRmal5tDGOOfqgyDBdDJzSmbIxC5
s1bVYrCHTh29YN2yg90eO5ljEC2XteSp+taqsUeQuUeuyFIGunldY3Sx1Arr2gux
zfujQn8fiXxkSGfTOpjQYjhBuIQOwSynnM+lE0oD7pHafZhhNI2+RDrmc9zhENUh
bfaymvbUDF5vMwrh/BGUhTdXgOlaM1ZyzQDM0e4PInEYIvx0zPExn1TqIfYCT+/t
GL+GkCabklhvWLE/BjIuLdD1eYkVgB+XBVzo8mxKLStz0qsJr7EB3ErRqj24oI3b
AWyj+x9eiUOp6AJ2nAlaKWuaYNhkNhHTmR8XHnoj0hTuHxFdVSZgJZJcAZheITb9
gVE8jm50FB50lNo1Clf/eLzcM1LhF84J/Rotx97KxEsrNhoWquOimwtWJRVW3I3a
rS/cIsdk30js4rOq3iz0O9WOJCPzZXUTylyKHoFYW/yNR5DnP3nWNoDi5IGwFAXI
0fVSIoFr+1G1KJpOekY/eSu0azdyZ2hruRJ2zyv5mCUc0ijvNL6RgoNFtoIIFtU0
nYdLDU0IOTQ5usI31vAPL1M7JVD3NAQ/G2mVFRFbRlL6iQumfygPw2tgoe9aeU+2
Xi5wt1qclEcNGzgOoSjP5m2bjWHszK03cxPmd1iDxw3YwI24Ot24w8zCer+t5uT2
tKK67gAljVqRQqrD8WKoOPnOBWcqE86tuvJGdV/tHPqYBfzSWowWnzZeVwdniZZ5
jUFO3kCLP+I1cdVP5BxtDKXjArcrGPJGqRscv4bpYmGXV8yA8rilDWoKkdNJUiFJ
5dzDNKV7r1fMxKXZA2O6uen7QLv+zUrtqFlno25ZBCvnm3LpQ6DZN9SZXpWXX275
5la+kAC6IPPbVpy3csgz7uHkQNDoneOY+jlxA/oZ4ggukI9tjboknztMC9sEZE/M
lPqknPiQyrzMLoPMOHSrAhy/+cjPOS6enS91rUocQMzbHDgYjwq0lWw7jSilLfas
a+pCfgPE/KqbpaR54hsimjbaLk+8oqPx3dHtZdnZIOrLosxnim07gwbxsfYf3gsw
ghqq9BWwEG2b/dCFpzAFYcdTz+Q+cMGUi/abnMJkGsnJO32BSH7X4nGTNIZ5dmWg
ii9jNOE9GaN22IjZGmzRdPShaPGoNnmIghUbUr1yGNQdOmbbwmsPNhN5s0Mx29yv
y0N9fCNLWMSEA5kh1GYzpG5dGwsqz5ecVMpeIlIhI5BCTrvQ/jgK+yrDuwWsJFUM
UeH9HH7wbfYbvQFpA88mhb9Efcc1eMfuNoy3cAjHcrQDFH5aZa3UHTWUEuFpvtao
2XGUZ6PMxKM0elrKFNElPi0RAk1t6QA2mPXw2JPFHBHDkO4+jc2svFeZEoN/gaHQ
6VmT3qeu8c1ND5heI4Cf78Ql53XL7wgnoKbJ2SYqq6bR+y5fJZquFKM7QP25162X
xbD2ZPrINwxNLQVmRNqwS1Rj6N17Y4gsrP4mZSEADwdw052ZK7C1JDZ7MScRvkiD
/U/wOL1wPkN6pVWXbNtaINQ529Wh8bV3m+eyy/lW7f7yvaCJWsOoTAmlCveuGnxf
tMWUtz3so7sCekLUJMlQQ/cnXLuttzQAdmG11RtIBfQqdznAIeSS6TwWUHy2sf9x
binbWAUyDfokflLRf0UFzqyNTybhVE8SnkgSLqo+8FrPH33b1TDaMCuF7heEF/Lr
V9zDG5sxhQPd8238u9JGyrBHDr3o4EFMQFaZS4GMbGlNbXYyj7NJrUJQD8O8tqG0
XeOW8wZCcZ2zHEZaI3MfzAVFq9wGUL0kDMeFgra07ShQVso9BPqZyzffqDwk82nb
ydF9ZMcd73v19tIzQ2gIMOVQZQxi1wNQVOZ0C5zt8Ohct7e6rqFPNgeYzDBPqQeQ
IbA6+vDiN4XCD5lXnxkgSFeXiN3hzRDPY9Gvqm4+DxKGpyq1AiInp9nfKN08HlW2
THc4Exn2b0Ciuqf3qknRMmNp/evrUxgEdm2/4s4AK+YB9HfA29fOIp2/mNuyQ3Pk
GZsWrIY+6DKNEPMgSAlm8lJloZLxkC2XOZK+bwkjeLKmi7FFOpzNHyICoQ4UHWRF
fc+NdjDzxm/4m3KNdwqmZ+lKq3GA7L5P7hDh6O4Z7C3fksQ6lrWQ8sxris9ubadh
19hOiD70wpKkPrLgfilaA4NyjStg+9PTtmZTLd5PRqhjTd/CpHNgfRuA3uJvNTiN
p65vKdlSame1NzgrL3F9EfZEyuEh26xgKkoz8e23+NzIQs71EvO1Ny3lHVZRbr3b
4b1TTeL3oTf2NRwCVEANukH/9U2vYHy1+q+sdgb5vXLjwLPwJR6VsByQjVa/p9zj
OGejZxL4oJlHj1YLy5k3DV/u2xFRfXqfSBsE0InX4Ap7NDAsDmeHsmJhBYN6wgiM
HBPwv5oWd1lh/A0CQTdQnpAe+3RbH6cmQfCC9FjDge2Qjzt7/ZZ351lfVzXDwLAU
RPe4EzsuTVeA6lf73++nX9e9QiwOoCQJaRjPF4vZS1DID4MUEYkUj4diUXpaAVLB
sIue+NL9gRfPjCYJ+EcWFB01KBZ8cHlXYmsRoTJEJgXdWvHe2WKd6E1CLG8g18Sn
HsuoQW4gx7FSxNQMaxtOLTOQn8oqu8RFFENUsUx6MXQw4/2vwRQE90ivzR1FkGMS
LBa5r1mZ7gsTpuk6aMjA0XMQ+BrNOPmoNCgmouCiVfpGTEHB9k7uCy5S7IbylWND
TE9jcNv4P0wVSaPxpX1/CSPSg2FX4hzWlTjQKDDhuVUs6EPT8rh3cmzuBpxQlPj/
kRDhhBVCrtIZ59MLTt6px/VRyqzqkDwhVtiQ+mHvIPJfprud6NoL0+30+TNcvQkb
uQpMwb9/c6cqjYAN6b+7sGAPZN/TBxieb6nM6w2VSh8kz5j5QV2gVP6YteQP3X7B
DTaiZKoFh5Eh4A6EEjZkb/aD/iriAkWLm84Y62nCkLfGPYUQNbhcL17q6N7UoOal
ssgHo4jwzo8H33uscuj4GLZ7z+t4Gcypyad0iDRFJVp6ZDPcjjpyDlsIJb9raKon
+C8iAc37Upzg67LLlACiGpu0GdF3P4WXnOXihowEmtLR23XmD1/E4a8ta9Oh28KW
bRMSR4cg0lbBezz100I8DQNe0PDSqC2C63WMU4l0N16oDEGnj7Vejlb9uH8idP8T
72AnQ1T24LvIZA6sd+6268k8NFvyqISJHmKpoUxEzNbogefLsQWdtUzalmUUzFjg
VlOLfQ3d1AIcGOxsZ7j2tzCzfLaVlAqszjoU2HrqNv6m0KbQxfol9nliKnb/fkUx
pQr/NPUOnmUs/vFYCZv431LrJfSLrfQQWZe9VKm4aPnROM5UZnGQWV6modi+hu2t
Dul4GKSjvr/RGZlkUz/RKiVKz+9RZK2rKmfCV/CWwHK0k+I7BKLEg4/imyB+i6LZ
bETcr1mI8CloWRNqLhpG/504O56rK10L9xgDOfnHYUv0BF6469qv/Ja2dq60OYIN
wQXAbuSA9RurCCBAn1N3zuf1ACuPnW1dDJb8R9S8A7J2G9KTOOpgF+vcn4wDur8U
FLK3o7sdL5rU4pZt0jD0JcbFv0RcNLIyIXMBmwqcCmD/AJK2ZgHM6WsFBn7VKZ+Q
Frf1anyR7V68Kwh+F0zbqYFaB8vIasi4tjfnzgotCeZMI9mGJuQfQQc1HlUQVVZm
eAhwNKWhivqkhzHcRSuxeNprGszU6XIYCzYCDrl5TqA/PDDAQH7ZC6oZZR7HOvm3
JLEfpLH9BuZrBykSAZzutK+TXCaMdFkryrEqDn1Yd1jEIKoSIkC4JIHu3SkEWH0m
Lvo6owNsEfzQFh+Afe/4Vi/QRkRSDoOuPJvXvN4EKJjlVCEb+6gzDch/YkQ/GF69
R4gLCXeZpEav+aG/X8VhN4RDrVWTVY32nE9nU2vhgEGc3SdtvsagZoKaWMWDksnG
YK2L0ndijkPDRxHTz6HVX9mpxq2Nx5DdpUEOAA+qvNIInuff7dXwdu46B/tL843y
+CVO7dsHT34Zf7gcUk3Ms9nMguvL7As7UEQIdXl+xJeUSUCHZqQvExX3h9y6p5LY
fjSdY4TGJUf1rcjtiYxLdeCYLEoZ1+E7AogHZSFCcLkxT4KQEhAqzUvZXDjUjyok
ZPdTlTviDYBUjv2Fd2+y8Lz6rP4Xe5a1oTmlWThMLYL7JaXnCnIJqykQf2HtfIxe
p6PvImIiA1qZ5OaFjYgawDtTxORBqDqX0d3uUrsgH3eP3595lQE9VM7JjdWhDiTy
CuxBpCQrMFBnVf8Es5iOjP89wiOi0LHSIaeMJJVc7vNXi8FauOiOmrM6biH21kGY
uVCmy7brqOTylmUNvUyJj2FiNwaLHQqzqzxcfsq1erkyalf+RX/oRKyUxeIJtlZa
vRtzBehPMG2DQZBs0WnjCKzXQXtZaIfEuAJdYDJ/DiX7KSBja8AZVmHnd3jUAZzZ
2sdsDmavyqWelO9TDtj0PxnF83/8d38wINZNuA/Tc+m3FfKDISYUarZKuFdEJE7J
h9ZyCP7hNjXHZhqIavkKPc5CyD2WEBW49vGaEjgm2U99zS4WwkJRpbgRNkDClXa7
ioORzirnt+FFoD2y1DAtpGsEV97M4OROOyEN8o4B8kXMASjJ9PNlLqQxECUmPEYg
+E1kfHIsiyBUjVYitM6OGHWqyFsbWnFBloOLCoUqNKu9HjhBR539t0VJztsv50+0
urS5Dd4yURJlXw1A2JbEf0mqQoWVsonO5k3BQqHhDJ3dhQZNomVY2uZNItbxEKg2
+YUuROX1oWm2lOl+u4tUhAZnYaU1g2jMy+TzxsLgUjzO0ONS6v7w9v+LpLsn9naL
MsN64uBUchaaspgFfw0Pf6a+dF6UYdDOhpMlCs7ITIqHXHzvM1oG+Zs1U09U1bw4
uy5IX6Qz4kmUhlEdXSI9196NLjRgclbile2Lfq6vh4D4VKJD90ibEQtICebn0Cqe
FFrxs17fUDcz2W1lJtRAvugN0ec7gwVVGHi0XMmEIr2naMfDCheHxYXweaL9Elx+
7Ma+jw/e671pd0F4vGtAo2r3mFaWCRLBEJAfZVXxhD59lFyMH8UgbVVW6iGRBNr9
TUO2Z6QGHTSon/OAq1sQzX0YD2C6/xlu/hx723PnmiYhqTRkAKTzMoiNLl1OtE9f
o3csomMr30Ilbi4r65wZOF6BTPIZ7BNcsz6xxKBpT+cowdkiPlIG5pZqSFryYDGj
jSoiPENj3qw77zn7SfK4Bd0YWUdLt4bS6Es8oxsBdForgxkzkWf76eBtA55eO/A3
3B9A0Le2SUDGpe1L8cmzoz2+drfcsVRnQhtZjWtOMK+AQWyQhbOAv+mVMrPVQFcV
LLrGtQsEY2NzUs5mI23Z0EoXQ8XrGy/HNZLWIBc3WXZVqzTCCKw+msrE/+9u8lj0
PQfvH1oAzy2k9F6GNo6ox2zm6z63UXISoO4Pw+etDgycN55PUAhfL9V90Bs6nKlJ
6wlbK3NqYSk752GGNx8Drn9kvzEPixrBn1EcwZ+WkN4UipaOBYBQo46mmg/f6oYC
3mzVmp2k94NBiDmSHx+g1iR5C2DjL+ta39DdDdMf8tG7RohsGR957P7911KpbhwM
7yzuLwt/rtthXgaJWAEFZrXyzIqgPhpdN4tFnIjEc2ywcIoAuK62Nfv8/ctMj48Y
aKAwdSyulO80Z/kNfUw/jW7rHTtNupjw7qv7KbXA0hWt2wVis2Gt8NFFh/BIvDDp
R0CoOIzUlsJFDYWwUK73juxZHtpsjdaHUtyPusAaifzBVOaS/VsPUKhY4kCjT+vM
SJdaYMVWZ/RGoMlAhcMZCoq2L+0v1h0Vee1nJVuij32CLSXAJmWM/Q8pWekZT1Wp
Q8BcCFJb7lxQdbBCtL2AB19C0T/QRQRFJtddW6/XuhCqZ3iA+5GqgZ9zw5sO8DUu
jDZf4c2Ds4/PeTUtCAM2Lx/IID7sUc+nF+N0JtUy7j+W/xH5sj73c3XzCdFVYZtB
dreYckn8FuGobC9F4yFlr/bqbSJ2u9AaQrIPnmOqGvWnruyfOYBXQl72UaQYx14a
HiF4FF+O1sCHLi0Q0RYb7rHxEdx4Qgmkhi78CLNMlVz8lWjYoEKwIJyq3Oisp9V6
oJLSZSSGreWmMXy048Q2OVu5uTmS/qFe783OY5DQUk/rQTdzJYwTlMtGDJZw9Kai
qzHKZOcjjUVH5SHJWVCxixLyp3EcUG4FWblaU9Gdzj734V9Nvqi5v4LNy6TOb6nq
v8L4F13VUJeFJyZoAuxjXZj1eQ5aq0CChjYM+5jeZ1hE1P1sa8GIZmfZdSm6hjuD
NvzAdvjJROwapR/7VRrkWclUMEQCOGcXUyGxaT7d0oooIzRbWSsFxH44l+h7gAxZ
iLWt9tXJ+0717I25977crtjmRY/Zj1WP3CuZFlm+qcukvQjsfpfaZMQ1T31Me5DD
FGCncqHJLFT/70ApRuXZcvCdS9H4KWalsLb1w6Zpw616x08J7wwpKNnwQPNq/PQF
c5pPte0oKOsY+s8DgeOnTOdE0Uf5C848DH9yFCwTZhTGmUpgHJTSXdTIw78yJvho
iKmiDNVya7Y0bQKUAECiTKXvqFmH7cAx0mH+ASwJmD23zaGqTuCLjLHfUo6wWK8R
Nq8ZEwZ2+k8+M28JzYSWG1oS+nqLRiZJZKjsW82YK3jeQqUGNRFaUDzIDxXnzupj
hPGmvNSFf6feIphp8C1Jjw41BaqWEwz0ydoPtzGYooRrAH8ZweseFnEMT5bLmbR8
WIvlTixdHJ2UI8+upNFiHG60sm2meEbm/BuUpV4BRfpKk0Xg4iMC7EilOMxkYzLd
Ssj7bWjWwDRj0i3hNn6aQ7YzHLSuZsN/98AgR6TvabDdBdHSti3D/Hmq3K47Cqm+
Y+JD1UlAv6rOZvaHN5EJzQdgIHLSZTX89UkTZPZ/l/czkGK1x84RuY6fp+H6Sr8+
MMm3AupuurqFmA7EWucFAWn4rA2XGwOJQ5amX64eVlsCLjqEOIB0dCLNoS3CX+9w
NaHTa6YLlMALzJXh/48mkQc4+xTM2ItK2247dFx1DU6XSpXjZcHZZgMk8C4dEHui
0rZ+Y7j/hCNyeXvQHuTnPPKu5orNVk8lc1lRgesLtS8ujBZZNHFYpUvbN6sJUVup
Y0OKtNGF2yKalW5VxBUBL/CGP0xXtKQmv4ZoGU81uDuP+FM/Yglxcdpuy0Xn5qlj
YxQ1Q5Q19Ve1TEriwl9OZmgNRXANJYXE9uIwq/qzamrNQsETZOagaIEF6m2nvAgI
4dq/nOGVNQnVoGlB7EMq0qlwu1pqk+OipGwMkhZ20TFyKFH/kvBenpy5YyNssi31
T9IpmYHulO5QD7AmPpGMfpR1U9loY21H5fgPkyFEmrkBxE9RIZzPzWVTtywpuAWV
Xu1SPE3iWjoMQH+2YIvQwh8n49/5Yu8X3rjgKWCa1uPfI2x8M4Xdr+9aia0IHgB/
HfQJ2GKxYQao0ZpK4RqCTd30rAt12p2TCI6grlEYWrVgwyUNdiJuV1kKBZAeyRyr
WUvbYd2K5z5eFzIb87gPgUlG7HZL3R0b7WHQ0kYQ9YAEKtZe6ltsdbCYZS/p5vM1
slyViaJL6Z/Al/B6DOQqvxOlnIFQUoeUOjaoCejuP1ptCVK9KdQUIpC0aSIkl69e
piPDl2JmNwhGST6UDxQFPnfLhLJG9xBI11oBV/8UY8Xo0Gt6pYGldPAKDXJyDemS
men6Ik7xVewE84DLTgI7aVnW7mWZZctivg83SJuVu9iAVKdIpPhp+sVRPyQpsZ35
IFrNqHGIxsEvqG//LygpePy0D5+dSWLVWe6kRttg8tBPKEbclfX8iu7YfIRooFnr
P6rPVGU/yDtuhN79+BJwDZlsWdtfkCq9wnjvJT4VS40zECXMr4le7a5WyqaTbX2H
y1nrSTWnV8aAxo+pFmnHS+jp9HBH3mUjTb1bjMFoZwUOAWXFCKVzwb8AZTBBXgnT
Wfcd7wqNeagsFTTWFMnhdpEWZs8DECgXzzJ/aRqFj1mpIO6dKjvi7JfEF245CiTN
1oPl9NnXXYUUZ0usUDqWPKzfrdYNYi8UEQGCMLs1MQ8sDUfgmq2id1MThn1EBVTY
eANCfkWwTWgj6CHW8RSql16UCtswQ4up2FsC1QvuAdfXTAsVoNjvf+g0n6czPALe
nlQoyUeK6vohAXZr+Zmdww5eG1XolKIEytN+CUOGL1Mxif+VJ17YeZQRiz0eHvd6
ZZYAnEuxJet4bhWjyWwb04pMnVaPNsGWYhMSBofQLJbT6a25sYvmL2lMSnKb6ad5
WD7FLAUYIzd48lYPTRQYnei7wV4N/70H+tlqsACSsDhJJRLs7++vAdYPKLSFg1L/
d7/2cgihDNFOmI/i/xcwttbXsPFma6cckPgw5bs0tuhVf/APZfqLauyh/6DhCJbD
a3vva/Iuj0YNaD8LRakOabR9+6/BHXQIg900YBhDzQh3gQDFLcECBh+PSCVnoCji
0Vd4zJ30lxfMEaPigszmU/x76O9oXPJ1ALYax7azKpfDKeEoqG+TQQt36ec0ihMh
+C7/hDEm+LcMZaEZ5sMYHwAtca620qnBZPaA16fam9b8F9o9bDDX77iZypVSMvmS
5eScl1XKKn35+2jO7l/pCW9gEU5jRn6etlH87Y9GYAEj0BlxNg/zQJi61kHwKpEd
JKXBAY5+f24GspImA+XKVPdV7PxphaM6T/gkvFjEeSeIJTTly9K2fwFQsLObQYg1
bwl86SLrNTvsgBH+adAOuYH4XMK4ge3saUC/+LyfqnK46YW9ObhtDiDxfSEDziWL
gOjpiWpioV38FaUoRGDAHEnNN+5Ch3Polesic/znALCr3TXAE3HE2QWEeOXUdVoy
Fz2wp8OtXuL0+k/Se38FRKeBAahXcfPcdojA6KzhjskSWtDppRK/f58TInITAQVA
A5NavVUqpB8dHAnsc8mq69vJQ0xFRdTbvUItBfn64M03lcxlE/dPkuaFqoxywhTa
sqGQa2ePcIP+uJ1EtSnrHE1b8DqiyzvdVJo7IreLz2Cog3xL3IXv4TbE27mY641x
De5x2riCqjJK+JZmG3S9XZlgL4QWqo+4gHs94NwmpPfa1/ApuCCkW54FAnAA7hvi
6opKOpvED4M7Musp3se5PU1W2s30+3y9eTP3a8Vy5jsWzZEVsyXQJlP4ZvKc1s7y
j+0Ua9IMUlPU+Jmc9xp0KO8278lvyoqRMkItSLODyzNXaCGiXfVBoOi80Ajwv+/f
B0TLBKovUlGBsz1pNAF1us0nn2Z49HS6fGgUpOKd0gU3L0T52t5cdWlga8OebcnI
HZsIZr5ALjYixhxmRcBdYCdhO8ZteTnX7fFv3GPLekg9OtbfL5bFAiKaKhDzTqpq
GAMhrECDLpgsPBmKl2c39VuUX/Vy+7FpO/8R1/Q7avo6V9oxSvcN9Mx8Hs3N18ml
Hbz7YnLIlpRwv/Cu2Ah6PHK1SIxtM161Voud6Zaua6NZaoQgu7MLXBU57GszLWyf
f/wPBPz8alje+HOTAGG2DNge/YqkpSRq/Jff3dVHifkpAncTtBjmH2YKhYYmD3bC
AvBaPixSSXcshrfDpwS3Gn/bOGVjujCjfpBHv4lMnggu9y1r5wB4TBIQHv0ldbVr
WdS6FRoNjIVMAD5nCar+pEsof3BD4A/Qtv6337HzsuOp7V0p9WDbNuvkJKTQdzJc
Fx2s09R9Kzlaufx9zuLkgQTDnGPKgtHRzzHyp9Jwprbk+wlAboO6wPLpt/F4glyp
adq9VgAuflV8I1ba8FL0qZ3PC9BqkUWZQO/ey2qVppc0SRJZDvw0Zqlb3OQ7InBF
yMcktpdEfRv6ZsQfF1D+xHgvk+3vv1CzZrX4HNm22qEVuI1PjoH9q4uliYsbn5AM
BP0juRS56e/v7kOS7PSn7PfthQSo+18HOP+gFlo3TwH0ag5aaY187M/5FMImYRhM
NgGPP+EJBhT3HW0MxV6FP9LfEiTOy2oYNZvU5R+eBbTnu4emVzOQQp9r3bRlfzj4
hu+zKmCW/edjADp5rbqD3RBx9qjZ6WC57QfgYs9ggn5B6Kv/C5AdfzLhfGPrxVuI
ix4iLoqoPUWsRUMOBo+SiiSd0zn+WTzd5LRgaM3cFC8jBjdD16mK/vSWEN141ge3
uJbLE5rPevcDaMWLxdWOvOpLRLtRBFhwg/OCNyJfp7Q91KKem5r6Yn9gN+TICXSW
dKGgXtL5OJxLVd4u7xVaZOHyAJvHFHDcijlG2/v0RDNNB6wUxkCTH1pAj+59cRF8
p2YxuZUP31ch5qMnfmH70KnDMbW9Eo7e0n7B4qnVx793L2LzYLYLcQ8/Im0j2k4P
BKjWLkkiewpEi3c1vxGbVtHQVyzL0QJ8qNC6+Y1Yz9C2lPPm7ra7eEPNlddDkLxT
useFU2Qv0evgUhJpYGcOlF0BAKFHmNYZxareZHVzxPt/Xtw0nt+9ghSUtwlvOngX
XRSmcczLsRDDPXVFmymSaDrCS1kSHIPREjl5k6+r7YCVuRlo78YdFBcKpqFwHHRK
heJf/rU/jgvAwvS4Knea2BcYjTykh9xppZMdfxyrBC0zTG81thht/IT4d+WhvH9e
F9o1rnNshzzT73RI3qRzXmB8jtfm3K4Y79bE3sGrGI9yp8eByZ2bFU26FStqOz/K
Y7JXu025RcPbOKGKFu/QVtnVfL6GAKehGU3TRrlNF++Ibv8oQBSmG5Vi7HVZtsZI
7bUHhfbefN3gIfxWzUO+O5Ozrqk5TcfYcXhw+lnteBa/qfD9ZNVuq1hPRxc2Vs4Z
M/A8n9WoVYqhNcEYcheLdftkQjRU5Pz1rVWCEBPrqnHQjmLuFZ0W4ikv2AOO2l7W
`pragma protect end_protected
