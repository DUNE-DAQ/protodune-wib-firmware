// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DWiTB483p22QFDWFvHs9SRMEFzziDLMEClrDS9m6UA4OWYqQ74KauW90GkBVYd6D
6ZrG5EdnK4AfXkxBLYmbykpGuMJUUNtNOoSSh7pw2tFjSL77u86htDGd+SKeNx/6
ar87f6D3wckNUP0weYlXG+4HPNa15dQZ8nnmtXh/Sh4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9984)
ZY2+87D0gpLO/nCoNz8NFtLXY30nMH3jtlld86uce7J3RSk5RKakKIzMZqf4x7Wh
HZJFhJc+KfJhHUNhuu8PsevmYX+W4cpJ9sudiQ1JD8O3hd5034Er7dmCdMaS999I
XJ20FJUcF78Ho2lL384ot64TPOVfxw1NP75ypV921o/Hs2gbD5BPLcSK22m4yTOZ
SqMDOJmJaVmpkgWPsnJTmiTASfh7Ly26SWD6LHHTnYRz6i0nII9Kv//y+U8MNyA0
5oTvqK/62uCFcqBGLCutMmgxPtBUUIlp0TolUGrfxmPunFufJwTJ9LzTniB23bIP
FI4kkjLYYlvMnOI+t4IjHEagqvQRAXCVPJ3FauRAptebFKsJynWB8moJ1Bc1qHu6
kpQZ43UTW18ZOlJo4gPrCa8gfzJsrDp+hdGK/Bm22bNUgyrJjSFWFY2BxdlvHnft
TYyefTuH57cC3YlYh99uw8NzJQsjzELYzX3yXJ3Y31kOav+TqCFUMfx8nTP8Vdt0
/VBxTRtJR587B+XqxE9qpjwsVy2KJaHYYECvdSEmUeS0IKAVFDmYAB/tYzQxXCIy
OzdvUVEaWpc6LYGjMBkAsfww5ipf8JtgFJTrA3EZKG6DDFq0Wrspcrq8YoiUa4Go
ylZkaqWsKFD/KGFtuDG2wOZ3Z28dn6nZlQxWlE12bVUM1MMjlw00fSw/a5vb2sEM
6B+027alKEyMTqQKvp6D5GPscbpo7QW6l0OtTGR9/XmqThkHVDdjVqEd+1uyDqUQ
R1/D0aOQl86H28Gm+8qK9ze08eLAcLlM7okoPXU9NbIDplONJkHsaHhX8eoFwNhR
6nCDXRqnCG7RL/bKo7TIBvqM3FsabQl91f3fWvSYOet10txQfAZkeB9MXg7bILCS
Bp2oP0P4XCRIUxOMBrGiOK8NmUL9G/QNQrfWP3mMVx3+TYj/4wUus9MelLozH8TS
yv7hQyXBGDj5JjAs3nGAc6SIjBOqovp9T3CZPZ4i6eQ3hBq2uBlBOe5K7UTRnUZd
Ymz4gtbwUV56Bu+n4JTAcyW+YUxWa83+/yPnFL53Zzy6NzfxmNPRg3d8GxOhIfqX
AySMkdA40Edql8BwZOfV6JiPqnW6Ud3HG58hlsyL7oAolgyeU5ZzFya0519dh9cL
uzmYzmTuEkArXCtmmbbaYS3wGDdHZdlK4ld+6SgU1C1Dd0M4pBa1husB2JTEOtot
QguK09f0FAANhiDVPFx7zsLkbxydmQH6ZpQRvKy9keUP6EGpD23+BhH07lFz/GpX
xJ4Q9nUYdDvBG1wOxCGUZLvAZZv+kEdvRqMgixs6ce3uZgPRaDr6gKkmxWWI7qqM
KxrS7WnKCwrjBu5Bj2q3K0jgmS2YITINuns80+Xx3fRvS5yneS5ImXJgs5bKQlcs
Nr17XZq77u0nnz4I4IZnjYQ/DVsqTYnj6zBV+BfYU/Qz1pY0O1jDN8OoyyL2RX2y
GcPPRiNiKD8SlRiFUlZLZhBMah4XA8ZxLZlSs4+uAiyaYxD40X/RRpSqJPovYYp3
vpqESapphFX5BnzvI1bJn2WzJQgc2hhq8fBL9mMIlJUcHLY2hmJoH6DKY4FDhS6L
gLei7BOzfVrZKxhaOWLTDlhl5f0Nx3NiUG9aY8KCCXA4hG6VvU6WdY/NQeciag8Z
MXUumrole0Bns0oIkkD3VLiUAhqddsIVu/Xqi7JF5/kYCAmW+Fflzc/wDMYyRDUi
mJ5hcszU1jFts+24MCbT7dRiYZwV6d4Kf6IwbIaX0Z62Pa5d0TqXbJ1x5mNiZLFe
3JJ2zoKwfw+50OPiPnpEkZzVl2enuLhM2Xb893v0mArBHv3dnW6Dt2JdO7GIJYk/
rc9K7MRYsBPDYSs8tum3DjERxKVFRmBoo611n/oAvzifOZQ29qipzRFN/KAr6j+V
M61l5ONkHJYiCrbRZ9Gyxf0uY3kgV6MU9OmDfpcne/Zs7Li0sVNYrKQuZwZRPRn4
/TIUTjii+zURmo1SuagXX5yhrr0QI0g2FwRsdDwKI3hph9k+olLZzWohlW4vvY1m
wBStS+RWcz/kOCmKyhrB0SEC2KsMlJW5b93RLH8PJAmxcv3TVyPwDTdFarUXPXdi
VbEIhfquuuFYfvvjfrBRbmej7kvN4xXnn1oq/bTmXUcgMacSWB+m3FV2YVMVGI+Q
bYG863LrQAXCwXKg2/km1pFoBVOEjtuXZPa1U+5whQLJM+cKt+uAX+M5scMSRtP5
jD/n0M0MXRdIAPYe/kljbzSTIHlVEg7XCD0QCPxzNldwT4p5EWsmq8ZNfzmd0sSr
/s2u1OmVBHcFFTWp/Boe0IoHvlUzejNLDCrSVAAdBHNqZB1ZJUDYN091Aml/+sDj
zsjekaAtGLxtxb6v1WDOMWCP+dnaO+a3x27gShZj3ejUT4RzY2G8VC5b39/2RZRf
5lpbgwbb8cbfobS+g7EvCafqELPUV8txvSI3kZhoTa7SxoapoMKd6xJomOWOqvI0
vwyFGk+EBq6CICMz2/3lVOFjr8DOdThmzhGEfqluxLKdeHQ/YU/XOrdL6Ju3dpbt
eksDZF1lcPU3zXqnyGA/lvthZ4w7iTRonK8DhFl/hZkXawRAwAnZ5d8Irpsz1Yqj
5YQm8c+m1u2G/IqOUJHoro1yW4dDaUfusmiKuUFWwSCZ396pgiFrs9YCm7JwpEXd
4MEyQY7bnuasc4Zkliv9h/w8iOgUO60lRsShEyhamwmi4pderpI1LVs2atoocKIv
wtJfmbhWX90GhbBOo81PYd9fkpLe9jZI+Rkf3tP86PN9IVkT0qmugPqLS25MxDgA
f4jYrjv6WNDHtZDzi4tS6aRtg/Xs2eHlzxSLqYeUENcBA2LeXTqYefX8S+LpcrQX
6EC6afAEc6i1wEca8MKhn1y3E9OSaSoeI1qEzFvGFoh9htBuHHWvHd9FxwRdaY1A
wvzg/WJa65yfd1rNN7QZGHvhQ5ZmzeJC+FMDYM8NuAQ3+rqDvZuFqIcubOr/C2t3
YJxWLCKf66uQmaXAfV+CyWhrNoam4q6DrBhTY6YzozC83cCCZQJYbgb3KJWPdt1h
/80/5AQ1LEi2XDapWzsBecsGFeKqZDR9eFTJRWbwVgSIH3aoXz991ghNjBhktKR8
TAv4nDeiCJNw/GVI8VjpCvN7GlTbRVeDbaCB3zfXtS84DYmSBwqKRodZKoIfcrUz
sUxvEqHO95NpZRCVuy6CLdZQ/USxBr7ImDfTNdSSgeLM7ay21kii/QDHza9o4hes
mBA+2Ez8kGJYo4ZcuQmbGLHkp6RO8KU8Hzq2xfKtkkaO5en05F4Po3zmrV/eTnXh
pJnQMv8H7K9r4ZUFXtntFzIZ2EKQX1p8TSS4AKfux3Mj3Gk7DvVxv3mIyWUW5pva
3DNEpn596uuorv5P4Yk5GIMUJ4/hI7hfVjSMx4B2zPXPw5ZhR/th4uXC2YbVnqlv
IJHGj9bXo7QPxHgbkVIsTRsocxu3OA4NQaiOvV+TSGT7+TywJuenvOBweayldcD3
RVUqF/aA0shD2cmZf6rI3rsy580NZ9UZFQ9Fgl4qDlTWWZnyL5dAsGnj5rqrY0HZ
BFioXvctl5SR4gmrT1P2BjPJ314lasRyLPdeexHno16oQ/Krnn4g4/40sBN3mad8
Jj7srWSVAuOA8c3UpfIDtLOaZqaYgmCjPQy7DoLvV4IAYM/O18wabOm2dPMgQMi/
hAOq3ii+tpKltix0Dzfro8PSKY0eNeyW2Yldw6SAS3CaGunvqF5lqdwWd9zZEDO9
LFVJaduqzKn0f0IkOjg4xtC8Yqs5rSvUyIwBeZ/HkCHQ6SdOJ1I5MxPYWSrbi5q9
rhii+zqeoN9DqwjIvRWntuY2rY9K5mXD74V090uUX99TOdJGu+WCvhaxxaBDmcxv
uFQF0Fm1hreE4TSA4zYovfQxca/5vt4IyH9hmF23KtAhLYdRjj1lWy9ADIa6Xkts
pQXOL6pQPi9dutQIoWFZGwB/lNpBtMoV0y8nWfFC6yvt9VC8bDx4f98XrSAOhC5i
5zxTHb3ibO0hwWO6PxQIdqiXHv0LXy6tlPrxISvDR648oBbgJDGcvfZu1alVBX/O
YfjrfsZzdRoxBb/oF0DF1f+9QKSHxf1HMYxIOzrNqzFvr47YBI5Jvs051/7sB5Fq
++Dq2gmmb53fJYxx31wSSAbStI/2MBTmlw0ipLFeOj4pa4KU1n5TCTI/BuYccu+O
SJtwXiy7fa76laH8IOUv0MyT+p2ZFES9VuY4W6ZfkBnIlDlr64SFeluYrWfcIbDE
bSnvufDcsnrxZRBjpdzvMaivFJHW70UtWz3FXor1YpZNyVW7KaDmCV84zxrQPAQX
SsKaCoJb7t7yfSoAdUsjVbTL0HSZCTUVdICtBYGWkfvmBcClYDM6gSb2OsSfb4Pw
NGppPSiXdtMsr6b93mTALwIWwK6WIQ6ayiFivo0rSVWZXHwMTbjXl+cO/Fz86iyf
nYgC4wkfqdFUYks1d7/c9CaM8mmqZ9XGO2gUXUaTwRCaN4PSs2qY2cwTqa8TSM1/
dYuM4ft0g8uvpwD/5N09FzyEbGqAMZ227OHgHskMH24ppMffGK+9fOQ9q4tb5liI
ZrQsgvnkpmhMSnX9/Z8TAuGlx+w0LuQu/MCUiyulnh19iGmakxahzSE6Qz2NKkwf
NPwMIf94ppxS/+cOv8D1bay99VAWblwQXvJaBM8L+FeAwqOQnskLz2dVgBM4T+gh
17oVt+WcZBvIpih5cxh1YZm/5kXS9fMjJ8x04eCv3d5eGGKfejR7MqFASVQz5ESY
Yu2hKdKNho5Jm1nzBKeRrS7y7KYZu/UBy65DalQRvzrQ2bl1t+oYH+dX3yeWUvXe
B0f1jdyNsL19rlHD9mBPFF8WHn4J2M3mXfvMR/UT3jPk8Xjoh+nRG+IujAbTwQj8
c9bD1YNUpP23dfq/uikvKIitUBGTTdAbtHTvNuCmjVaoUuC1wD1LFwboieBoNJxF
LddJh5KvJXJLf5VCtI58pPPEfiNo/BGcJ/3qpK6dPyN2TVg8NIIt9YjaIK7/Wch/
lYnCf0hm5QfRBN9fjRpEKEELgAONWE5I1xmwzZZhUE2gYQXuZ1mifA2fp0UEaS8o
dqDq1i3bIhCy/dy1FRqJS+XH/ymB62/D84PPL7QqAZ2TDTYpktb1pzwHlz8Roe4b
Ym86zmqYDr8bSn9V85ZAVBcaUwMEceVSvOhOIY5dS/6+wv8E1OmK08ImkwwqKGH6
n4pYyvHG7KJU0eFXYx0cLXmp0I9544/zW4sjv1/Y8YjKbJ+PGDJbKGVLU+cixafv
iOWGoN6B2Gi899WuAoH4PLr+TtA8n071xmqjq2C4fpV0VNYtw5E6knRw/IctLG+o
6edYAfRUKuLvlNf/+nlbZTyNGGSuinrfct1asDoUjfWcGY88Ze66Tr0tA7Tlc4Mu
JF2RKRS2c8GzPwjq1Mbr56iiZ88JD1FRQDTCw8BB/m7/P06GFK3ISvZgZu+TMydM
pzTnsl5GLhjnIRd9iVMCBLE3Kp8l2vMdiimSuIB7xvSBcvSqc+ew5S0/KgizLtMw
Gm/DWhPO3uv35KsMWBk+uXHJoSy150PMVD2696FIJIhwwWRMw8Z+JmUFcQ51XmKB
vY5QKRDIgL5XjnNXvkeiRG+GZegqPGINhcoWUsVlt2URFAp6H0mt0yj1WF1ZDdgG
Ryn+ElC7IdApBZo6CTHzhqsHGlxqmPVLpz7awXSXyN2b+okb6EPQQDR8ImPf+4fF
sWmaU6cN/af/q8RHbZVBZoK48yf1NvKvR80ZP/QAPW0hdsSguRcLeD/ASpWqAZ81
BL0yG2HGm4roof9AThIsjzGkyn/C16RUAtfSpqowmKo3VHu0Im5J1Se1RxGj1Eh5
/1ftnTqjrwauZXRxPhCQxfbJnI160KVihnXL+MXQSNp1XeTtrlxga02fRjs805ma
ZWTDL7In89gnJcQ44stqbsFGARsXHFVPHHFcrtaCQIvbk3WEiMf5L361IX5j38Zh
4dWyx0wNczIHDzKdQEKaDvR5a9HSHD8DvYgtYTzDBlQ2KdncOKRItR/m+mfi+t1F
VJpoeL93NdbBg/5rvMOQfn89CDxrisZtkQOOwqSgEuBp5JxmzuXCFCdOm41XAvzB
KzQnWfwMGkeZkRv9fo1kG5MWeVueS8WeSi+8bm8LUu59ed0ErF6oXB3w1I25zTpP
Prp5GJM+ryLe+pNI+5mVW6HNZOea5fXYQBmHSJuSAJ9XjOdDeZ/TLqaHb+3ulaeu
mZkxtsdmhUgqrzsJcnGDcok4xZNXm2mGjX+xg7r1wmMkgqwrnrqiOjCjigVUETa4
13XsA1W7wSntl1wlTTUKgfWNisyy5lHM2ImBwVEMl7nTL3ops/ay0gjyxnoNzPYZ
7Gp1ofM4Zy4IaGxSj1grj+QiIeOsATtaNZKZRR3rlKubzDs2uB4tLorxcLD/BmYX
paaJT51WVqXOpaPQJEfLf+e1GfoS4GMV1orXsLWMWI427t9xzNdSyDqTEGtqhhKl
Q/KyuVI/UtxeQpc49LGF7u9tBMXeVGb/igZduzT9OTebkWJT+1eQTBD+vXHX4+us
8kmlE/6Qaexw2oAEJIpFHWXiCge+EwmRYQXwwb+Ysus/uFqT/tWFmuKQRjL750Dx
HQUGbifX+erd040vtsEPOaHnADiwQl2UkRYD/tBJ7TsG2JhD1z24SgpfWXNET0cb
DWY66xUefI+pVy60+j8967KpRX8yr/iae1VETmGCNdNf+FCzNzDhWcRKerYB4owg
jB2jVToH6qUbDUGaRTHXItZl3yCC8oGqZYMX4hxYuntyNz0HAK1mOXe4Lowu8mxR
06E6kUrXoELKK8otKif+Vc2jgFAPBVwjwjywWayHGKuaZzHWB0YkcZlkt1lrMczn
EZH34OnSw8yKWw66xyGrbsyO57SC3cbe3HtmBOXy6TlMn5b7W7I1SO2eJVbgrPi1
gLzPXZ2VKo6pfeLTgLMUH5Y3LMM6gJ6vk1wq3TAbC8Rtkc2K0FGH2W+QjymjoX6M
qf5jOHfjUrpV+00+oNqFCxJ+GTPFCDJDYofAz2evYViWBpcKnlBchr6YjGkPPDnj
zgYjsSmDc7bP+NAxHwCPMzqW3S3msQygDaCovlPy9NdTvD9bvF2iNZk/xz9A+kD3
QH/p79N9JilMyVGguFol/f4lSG7xQbiitra+oF9fIM6j9i1JwNmVOzWxJG49rO28
k5Dkw+wQQT6kh7DRQ/ocNKMn+kMk3XanNuh4jEXeH3VzmVw+cAQf16fYEiI3ltmR
gf6SoMBp85eeC8kMlyvV0I5rPF2WMBHddfX1fr3ekBqtrG5TehEeEfM8ETvD34qK
2gNkL6loTeJHhOgTeBzIfp/8YtuJldHsqY4dWb11dNVRJgY/F1oXVMxPbNWdmoqY
k5OdWjmJZFyDWUT/I9wOJTBe1PLKBtowaYUYuWSZNedP/W/FppoNfIhvu6WzLtYV
Dn4X1O95V9qZiVgP3VbEXTaR8qNLVlg8T3njIosGw5x/UCdYM2ju4vl+8/+8Ba76
n/ojUEIUCNzadvLIidZcDOz23AJrdC0VuRs2zdiWFUjzlp6MkaHHTlwNBlKDUEhz
pbDpHFsXwJY8wkxYcEJP7MVzDtpUaGzz4cFhGrRA44lSQgTLTrQj3EQipN0kqKQw
O3Qc9UUM/X6+tVxwRvXbj9gWvU/lfNzsLvRyJU/6DkBfyjKWGJVt3J8CxnGFdwtL
51i81lH4sQWk1sdvGCIrv6kC+bJuBgtZt4CAPVWMdIwdavydByYlAXPw2Z1EF8FG
cv5E2SVa+Wmv6qPCdWeA628Hmzye/aCEX9/EG0b+aeMVIEL2dNyEl04OltOMrR63
ZjLqBb7rZZQS3FXpV/GK1LlQ5H0e0ujBZRxxcXtyhzebERw5zSwY1EbUcgkUqWDF
A3s9oXjIQiANJBc4RcrQIdUSYcVdCFxdyk7gRr3+kTJrCe74GFidM8tJTOsZhTwB
tgSEt318o9zr3C8ZWX2suRu4aMicGyvhGS0byr5BLsNpDXaY32SnHTXJPTT616AN
SXBPZSLJ3lZGSfj4SuMPCLScKSKM4luJ9WMeza7p6T20M0iODPKcV/2koGep2FZ9
uPDXdZrcL3IRdFMK6mqSTMbNlUDdaHsoTqXS47gKVXUYLTlDKEQfMS0X8njTqjrg
oXlWhnKIU6vwP9IpzJqTSZGQyVNBO2IwadIJdfsgLiSohz6bLFRtmdLH7O+lQiLC
cQh954BYKouDDTwRty8sMRyIN6nvhLhjEaWan9UIx4190s57u0+IrXNEgck3Udbh
8VzZGKUlHWuLinD+DrGeiQbpUkJmLnjITEj2GmOp4dtEPBx2U1SsR4Iju4EZuXsD
8PVKrGinO0KmRCIrTfz3YL69boUsnh4lIks6KFFwpLNtI/CW8jXQJs71QCBs7yFB
rjS7Fz6jE0CvFZA+JFv0F/eod55PdBgZyFRJlmseVV8E93hf1a4HUWWpioOCadfJ
wGyDyGe7r8LD2OCt5+LuV0+as4nnmjeJilA9750zq7tlz0L/RUybIyPIndzVsaru
cTswCuK2OluHnCKTxdk9MKxhXWudS+bOjhNOQyZaaPQvw9NuT1benSpDRODVSoIN
o3XoENSpiL3RL8+gdreiviBziyojEr21oVlLJNPJU/pbIB7bopmy4/tmvqraqri0
wDH3zUTU32SvaS6owkxTxY70oLg45t3XoBQ6Gcd4OPwAMgH8pBe8pMFogDs+7ZJb
RuLIdzxoST3a5nijoTngn/93a0blwlF08A2mnpW9SRiY+tAxeYTR1rAM5JrUWlJv
q2FdNjFgRJZCPcK+ebKoPMklcGiublXEpDydKnIOroB+JoqhrIdGXI84/M3Jgp5z
U7A8/6iagFPgWbcDnzAlJZcQoqknGzV5qrvkygStQJ6cLzLxY4stU1bmqGfvQcD8
Cb6M4RhmiHXYOqGGntJ5Ob39EE21uNAKaa8VtIL6zVqtjyvbLi3aQ7ThJCrKzLQl
7Xw3Iv/Xd4n2QTN/G/K/HZYAusB62ixRfRH+KqOkC35lZsr+wtrW9BZ1RZUE0pZo
0l2+DYYLwJli3vKqSyXAOdNTboMJ9KjlgqzUFxXVbQ35VAQyaNfuDm6+BwgZep4W
cLXHzR/s5CfnXF6dCVx+CJHhnoo032cOyMQS7dyM/0CMICAnyx0shG9JhCRbKnxa
bfNl0z1wsGsSqdVwIeAa67fhJ7nF4mDvGd8ESQDzs2A/clzn5b+mo6IxIjaDK5w1
zFXoCb2u86AZX4xe7/vUgzOpDQeC88Uj+euCj7ZLpjIC52GmAow09JoTgvYxHYW2
BIjXyLqy0DwzYCfRlcNVsD45c9A+Zswz7VKtG3k1XY+ZXzC7WGto8azz8rjo1HMS
UeEi96qVHoNRfrQkbhJV9uuSic4lcJoEqg79lFgFiUUo57UTg8drAG8muweqpZo+
yHKLHG7KNaNcc5Kaqp8L5nEU9nIhzcR9OTMUxvGKTQapbyOV2H7KOd9oPjqrO3cW
1O8TDDMQH88VKqPBmnTeVaVpZnDfH2B1q83jTWCfN+Ati+OGx3swRCu+tiFeoLXo
uTjpqgi/3wWJZD0rH5hbEs0WJ3ELHx7NSXqggiEDKsWwD+Z3K8rcFXJN6IAh1bKT
8SUDLplfnurszZpNAzIH0EERVUcqjmRFmsI1r9qrm8iGxNVtx5hHGSzK3swFrRQR
3fgMRH+OFXyH2hBrpXYdIO6bPP9bBKjGy/XAm7YoI2Y7eU6xLSxsTW7wZf6n9V2t
pRCaVu0UiK+oEfDyjbRymauyjPPh93oc0zJ/aXsquy2HiR22mHM2KcMLWoR58ERt
THboalospgCGH6NaKayLu9806wYoF+PVBzWd74SPJnef7RcnHZoxLywtMtruENub
hkcbukCt/x9fQltluMXCQExT9ACAsD9fQNQhHGnnac+D5EJ+De57mM/6CEGOYurj
eLwmawMc41EnyA1mFGmjHRmKpDfq8IM/VWm5KvHgNO/NfZi/7dSIT9YQxyHE9t0g
fovUZi15uVdxY6OWadXPy1gSAU0NPQjj6Q6Gr3NwrBcMyx5OD4DQYHAC5AUGlOmZ
53TnbNcRXV7XBPNTH7VBoI7eg525bwb+nf7c9QphhTfYfoo4CaanjQdoij4nbZjQ
5KRTfYUQuTxSXWg1k3gMPdGEkgl9Wf2cs8Fy6QqmSahrH1O8CQjc+0JwfWr6A34z
PxN8BXgLAFoMOc2spf6cet1fFaSVtMijixmkE6UxoZ4iIUHPzO0beS7+tOG4uhEb
3gZf+RqV9l8v178ti0tI0XPpyG/9z/hPLXo4MmRLrXheK2bQXJhVw1nLPTnixUk5
brDRLmlxAt6QTjPpYf2jyIxear0AeQxacPCYyZteDXEIQtGUtZEvH6d+k7yBzgd3
F9pZUX10Ep6m8oYUWmeMhgGoKVcCejIVtFVI9xjI0AtTVl0VO+pdC/NqEmbNtE5H
RPyP71nXxLOiZY6ENSl5dIgYK17fqKtcr4Nej8TXHhoRuXsfx9olOFdQLZDJQplx
15juCyxwgwOuCMyoIAqg0qro/45JflNrcOm3A04ilyefOdHDla0hBEJ1lr9vc27c
7G7ldmGo5TjY3hwUp/gq0Hr8uw7w8MdO/mkpQNKDY0ELwomwpzh2slrTnp8ireMh
rhTwo4pwqhNDZuGC8NOPRUfyk4HZ3x6NRIaKhAOi1tAHtAYLNjqLR/agrE5kwP+I
S97fXENT8kblZVKXqHYgyHwfTXTP9wQgvp1JjJWa1YK+yT2WyTj9ZrN4ZyDEe8zX
IunvWk9atTd/QgNtbgy6WzU9EIBuxhgkeI1cC/WHzRRSl2kCdEBrfnqlPbpr6SMl
Dc1VQfRO4Jw/NvZBCyNEs8HWdwHnvqfnoF/23nMvoCrAyMqAc/i7s1VxLKiWn7YX
i9gAqzzLapCjPVY3vQL5MZC3VWvNgtzML0ZtgH4q7f7z5jCyVe2f5kpFm2mShc/O
+doo7CUbaxHDlnIkJF1IXDEeWPrkE5Q1IDN3oQPp729cpBOaQdju/CCZ6e19Z/qz
pslAYqMU5AnGxO0PuQZxhTi8acNyySJNg0oPYAHg7JBTAPkqV0pG4UszL72AV9Ws
5whm0hucACXCncwHEdufvV+sWmUv7Y7WhkKkBbxU+1vyWtHIuwXcY7FSq5/Y1YN4
It0cE1irTpXKNoM03yeaCCGkEnjnvx71yTjnHHDMl39/PS4wnYNHz2VL6HyhJZBS
zi1zxAKRwWPDn20mWiyfrXuoUjVhTq4p7k9SUpQsMDepElPlzHUsk1KyOvuYpEXc
v1/vv+yKRRbfH0xSyOHHKuFxIXXy2ZqMAjWBsr8iHXgn3JETbbUt2p4YxRwD9zzC
PfNtt5s5MgfrctaUId2kLcQ8d1LPLoXb4CTJ5fY3YKJ+hJuuYTbaDk6+ehmz1U50
eIURNHvtdFBQawjQZvBDCXLhdb0oKsnbq6CvGR270foC1tl8Y+qwqBdLYGrgMZJK
imR2FXFQyO0hthCzP1UKvzwE0pRywUwFXW5aHruU+W+FyiLIk1PgZ/hd5P8X9RDz
1NHq1v6NKiDB709IItAPOs/XQrwgnbVH38BVzkWXvoAZjuNwVUHNyNIqmuJ1gnUU
JlHQhueYcRV2e0gJ6Ad9O7/kG9jT+vSRHsjgDggf1AnpMYv8r09qaM1PvXLeqngW
3F80K01GtgquLDAr7efAU+j85kaM6q0ymVQ1VPA4/Zbv8tJ5alp+MBatSMjpGiLh
MvJD49tNTmU0snxMiSE8TbarmuPo9pc0Mb7UUG1gwcqlqc5+jTgs5IBXoZknye5Y
aaysEjGvFm5YB01arCnaiIC7hZCG3mM9aE4gsg5Npun4v+z9imybC3N1sOpvFT+f
w+zzI4/aefkt3TV3gIB60x2yQo1t9Yp+6I1qFbWyYaLfKTcYwZ/EVsaPW6MAH6B9
OsUk09u9URZnPqsdqbYtVsD1tQ5gqY32p6NdSJyQWyfZ2EsjPd6n2Whs4y76vPt0
KAUjK4pdatHLxeUmGVt6Ln/XChnnXcRsrD2g4Z3wWuYLI1tqT24yPm+VJPl5Kjao
7yloMmZSMfpX2VT0/fWRRVdk5dD4gwHd7je/vp6A5cQTRXURzqUWJAje/ueKhLYb
sdcSD4QqVmSGCDPf1ThOSnQbzlXB5b76UrmXgyhjhPW/+ZN1sbmzYd/DPPsSBSCk
/CmcNrBlgO++nB7QXwXUOwazC/vCToGau7FCuMEl+wtgH9DLaAVfTTZ2cWE94vR3
yLiQj9Eg0DhFtUPZhgbk4JLa+02m6vZ6Wz1dmAWgam8kJ+CBWDNPDFYBHGIKB0tG
16tn/s4ow3HvmhXRU+XWm6Rvjf1BRlI9oSQ8FO67nBOe2Y4mAXYM/mMhoclM3Swf
tr9HxNbxSYcLH/DuYXdOclWEDng/QGi2SiejFIhTtuLZeEpkvQt3/v8yxBJgv/MM
bqS82EHDujL7NMvie7/8FlEN2+F1ALiM6rUnbPgBAmOMc6dSSW5JLr+rPDZ54hBn
M8in7ZW3mTpq9yFsHaXyI20aWvzmROdp+xr948JCXVFtwDuiRb/RBaS2VDYNkaey
ge5iXUoL+X/vT1TumkBC24O8v0+rFYSHT1T775sCaCEWDpwwIlvLnH6yyr8uW568
5e6X/2Lwd/u/OqS1eVL9Vn/6nBxzNLRUvO6yEV9jHvrV7Cx3ydHUvUNhRKtMPFJO
917mZo/9XaJNqCLKhaY0M+H0pBfxgG0G7Pahu0zXA4ouax3pbxiF2zRzeMbLu//o
2vdB9MHoFbM9OmlrHMw2zV0Zwm4kAzOmq1IwumQJkgcviHS5BruMjOS+UvFMlnHD
TfrJlQa3qcgg4gSo/p1t18aiqkdAfp0xrXFNj197QuLESjuhEP2mtLnJzR2f2p7i
DW1N5i9AMfRIuvD6/kvBdYoW3wszsKvn8uULW1DJSXtPq6gOKBlMa/6qWgs5HnF4
XJJldnGabGwVs23/xPdgUIINHDVOIMJ4m9btwJCjBiKBx5mr/FZAxYVHVh/nDBOV
vcjsGMRGdtZYuzLvaX4VzcVMTMd4z64G9+E648eE8U3m0JjUgvCRsjwvurUzPc53
Qq4H5+T+oM6zTwqELbNwN4oiCbiRPsu4x0l6Uzew5UP5Ny9fiIsx15wVSN7nuACX
vCwZCBjtIvcOhoxZhvlIq+feS7K+vO4xZK2UbuTLkGibaL4ryaFcM9owRAUf9uO2
acuBBvOsL+Xq7wdF085g6ZwSlwicixRtG2/xIedDtit65VB/W/iohVsW1l0zzyjB
`pragma protect end_protected
