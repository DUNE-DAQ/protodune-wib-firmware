// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
m7Nv0qhKZrEfrUTBByB6Qc4XLkn/B1LG1yVoTAhNYiRuX1yx/b5UrQ7uZvegJGPt
dsU7xckAu67QLe8TT9vNnSfOaRLT+uQ+De2frEZzklDdD40M+tJ221EeDgF9vFlc
/RWB3Wo6fVyQHdHOiErCjjgFCfDeD1FV98tTa67b/GM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1728)
xoTDhNmUChzQA9ghOsjY1+L4+cqRRQx5mxBdOfZNle7u3CC4OvhrfMXIRLgBH6aB
QIfDQlYotgIBqR8U/bCMpHwb83dZCPgsJjZyHs6mmPKuJd9gQqjiZNuZ3gqU5Eep
qz6CZjTzUBctBC6YP/9dc6YOIBN3qCURprClhd8uAC/dFx8ov6xuP5FzwtdTxd9J
sMnvshaHio2ohwj+idc85DAIyzIgGltgX5NKEpoGWiMO+62djj7QpyH8i/N4dWLH
KHXv+GlGga9lH+cr5B6ZF6mCzx3kxDAouw5/tejcIqznUPomVMdVqp0vynD3/zya
v9k0igvLzuwd6Bxtf8x0igLKAmKi269uJspOvCB2ao5D6zzlfYx4GCpMwI95Zn2o
35cOwbO1ajliPz7veiuJCsk0dp4R67TGbf3T7XhiVvHEWweaerXUgcYfRzFmRnQL
AUwnMSNFkZOzsVvm2MLGzrgYiOKt53so0u3rmT/Un6rno5rjvKFfj06QP2OEAI+C
XcmlGZhyQs8ThkeuelYmGHBPGcGP+kPyjcY3C3m4uCtlygLOh9yeOcRWH3GY6tYy
K2hACBSCLpDDZ69xp+0+pOTBHGc23uS5sz3dG1Ye8cIJFSQzjBomHsJkUMm54AfW
nlL28x/GgXVJuFXE9sJjdGhhxyBSpJ5Gc8V2EaPSgvtAmugake7WCD075OkSCvai
kGzBtP8ZG7IcP4tvYmwxIwsfUcpIcHYN2JS7puiOrNatq5ey937Ck+2z6pKHCqty
WTukNt1K4+J8mVROOHS2yFOdfO8ShYC7FkMBycdPtRxfHGduJMaBLYDAHsuKddBW
UulEeumRAf91y3yuBizOSvMxXq8LpRcZV1IlgwJMQz/Zo+5/4bf1aGkqnpe2ELiV
vi24hsxyp08b2uA5XMz3ap4iLA2/6SpkfTWmewpePQSj54n9+VAXhOloDzNwxkWl
IpkEFS/1tR+RSFBjS86L8dH+7QObHJGT0MsQV5uSULFHna15Rib4vhAXTQfiWQ35
6drENEI7o9YYYp5s14rJuC92pSbevw09JNUqYz7uVHZFX7JYsPurZQReTO7ZY+Ya
WCQHGjX1TYDxPbitu35jwaiMvKJVb2XCy8M6UBcBJXE7B5fCzgybYuQYFlAGq/ME
QTSbdFICLgxqdK63XKq8ZWZcJEO8Xcdw58JGi4pPndu+lWFe1x19AIuX6QXy+B2m
+gdKyfSBdIAG6y8G2C1it1FqZIri76EZnK8t0P2q4BydFBjCpjwVnV673fjmG8/y
dd5uKNwfG+oWyTxT4nDhA6z7ePtCk8Tko5C7Bx5E0lfZox6kj1YSNG7K2DsHxfFF
U3C4TfrdKOjzcUWmBDVDQHmqa7YpN0ff2sKX5+wDDWhYaDFD8oYgIM9glgodDtFU
PuOd9awuCsYonZLnra8DqKhsIHpUqj3xD6uIiniLJLV8inx3kwakr8sN3vpFfKMp
RMWtGB20o3g7s/ZBIRlm+r/85mfq/zRh/kzBUQRwaiIpizzNyyUABauC9FNFElfR
GPY5NxIW7ZbtwqLsnMyVMM8LE8BvsO3ZQgDhLP8ny9DtYQBHfUVZdX+Hou9i6cLS
CMf7zdFI3zOsUM4gaNeLboYgeE0PrWY9hJRuLmcWl8QXgoMM2Npg11MSwcSrVsfZ
IVplWmvNAhSsiZn6glZUVg6SPY9zj6t4dM5ebtJiAP9hC3oi+5kVqj/21rLx8ZOo
9JODOcT2twuwVSyyxDm4CLuM979VewlmaFoYJmr7+/y8ydIFLZpW8S4hK69i//B0
aUOu26og86p9o7aECUFt3fa/9s7ltu25l4KX1+NhYTDr2B1/39riOxefT9NdW+iD
I53fs6t9xG86C8ze7a+luSVx20AkYWotAQmySv/hv8ToDHqCyD/B/DWySpMwi8k4
WJ3KYZgRIppu8wXtpWuMqCvL9Qfm5XT1bJQuTIMuYkKvHTeR+Ks1yVS3eSmFDtOI
UhPkbuXXSazBloyc+ubm4j3+fx62VtKPl8A4ud9kjfWlJ5KSrtpcAJJ/fN0KmFsU
HxRE/r797UUtZ2UjiSiCrId0k1ZaSwdC+EkqOUrSZ/aXoa4yEfNQL/fDtU/sweNb
ingqjviPNRJNvWCkyC02pOTW8piwD7m5GuUXUmlgP0rh0umMoM31IhgRJFoiAqCM
sm1klm+8LgtJPdTnMEmOJ34aCJ2x9UwiA1JkgX9u5AsW1JDSyFM2ItGaNrxIsAfO
wMsrPl801B/fDpz/tPne3cyI0Tz3uhl0SrbqkU65jdENsF7xLAeOFY9IB/ZCE0rz
`pragma protect end_protected
