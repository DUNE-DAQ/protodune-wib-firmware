// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Br0NGyPrZ2Xc/EORAgyYelKPhSIa2Glc6+el3rp9NQ293gym3oeFA2M7/t0+fLSF
936ugNvJptt8Endb4x9I54MtEp5FE89D32DDEP3S/YhHNmeKa70N6DX9ve5Es4aM
y8+aMU85mwc8qqLIgRIcwzf+kzyftbTm6mq2K7c1380=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3520)
wjKls88vqX8SujtsAlISRXgX9eMU/sEaQWkwyanxbMpFrt5s2Nl4CXTFyFtNAtV6
jhLhQGmEOZUedOaGxbrBUbvS9I2dYCJGFqj0XBmySPeNrB/UuO5E0aTaSdTIxKt+
OYfAwiwr9GoodoEOV8g0+94Cag9GpfpPPD+aeVdA1audRvCZhDvfG9YLeLfxCfeY
vrukEGOhwCdhdx/1qYClqGZqx6psXuVESSKMZvognOdiMaqjwmnPyvYn7/Do0gNG
PITpPTCksQUWVKDefEfVeS4S2Fok/0yriOJNARzCUKxAnfw5wlvBrpYpUcChFip7
KL6CqEkjrq69YPrWxjOplkBl9jR7TnczVxDNDW7LEbeVzZJ2WZvXjSUGrnp/lSqQ
Wor9fYHe+MtEbmZ3gBdjP0fs+WwzyvcY2YTYPDre4moXpIVGl246Yd9TvrzK84qx
ZYZU1X2hnEYns+1Nn6cz0/QOkgJmASvaG2Gx0O+MoklN4tNrX9LjHYwQGozdy9SU
+zWbUwtEvkeB1rj59Fw9AlMqf14H7GY9IQ8t+3xyF6+KSj+STs/5ceMjiAvJkZuO
qCq7mZs1ZEaINYdCcmMwH5VHf/RDPSEyPyEBgtECHRoORAW7nbCiR8Zu5FaAAYN6
JjogihdyD5P5Hcnx5Y28idJu7om8VOmpqSzpjY1URkhbwuapsZ/rpdjsL11Ccfne
xks95oWTkEbBBQrmj59wd4Ra9fDkoVjBIC8ZTwVCXaVVerXecMPwkuZXYzpSrwy3
qQWlmbdTKrqc59CIyLLgMBB4QYLyEwZOgtZApK96usOZucrPdUmte4c7BGti3bSA
MySqW4K1VIpoF61PKlK0gZPzMs6E2i/97gtH0LcKTf8Wg38xq5FZuBEl8iLV0bFz
pstyshPJdlaA4IXxq+vE8jR6/DilA2PCMvu1lOny1BQ8146KRp5CPwiH0bqGDiyP
3tTSmQ+X6CKxgP50YvbbP/hXDxm521wvf+rNNMw6vv+Hf/zlfBsuWi9Nt5W8aLRA
1+AvshPKa4lz+GJpilp1wtOqqgxmHpDPTOTD0QpzLb02X7ikAny1IewpSrhDqZLy
5MIWya70njO//8bLDWKaL0pEWHXCRY740n+aLPH/Y+Zh7uPQh5I3R5WO/U9D5/+Q
tx/doNiB5POinpdkFdRjvTwFSwJxNQWtWlIG1bfXNHVdt8tf8qIFtvIlnBpeqlGr
x2rRecFWvpjsavwCiqXGtzPk26c9NUVkso+Izhdk69SVoJeZBUCYeX1hkGeYykbJ
/Sxw1VwOCPRx37vC2X28BVsnn7yS1KELVjwt8h7zs5x0I6k7Xjnt35zFTlVg7vow
L7lWO7vZUOKQ5MrZXuJAu1ssU0zw/PskR/NG78LzV7xyRvEnjx7sFPAMs0pJrdA5
InTyOUmti3utWkriy1EDJXlF20+XWf1yw74xuHQK6eyi5yWBvFEgjnTy5Tjk0V/1
cy8JwIQw3v3jsQ2Eei1QrfukDj8MeEG+3p0Dot0vEbF9suZ3AlTypAnvZ29+BO5r
lVcA9w4eBDFNtyZZzbv1KMQ94M04auFrWWNG+IFRoKen3vGrwBMZgl1kxgw30Etc
n3AZqaz+SII4jJOepX1CrLaWOoKMgNi/BUQEDVDbnbjv+suUMeh1WniRGpP6jjPY
jUqFcfkfKiLbXt6FMjdwe4n1ByDaKhIjvDxj4kEIi1d9ascXLIcr3SAxLC7RoHzc
7iHZPYLtP3sfMvm/iM5bJC8LV0NJiXfoqsB7B1f2VAsnC2aSYQYX7AZjRqePV7UR
wX7tnFfwIkTOhMGNlrTQvsxcOgaKJy0W7Pf5wzDoYW32BtPgpT0gmBgmlbYK+YO9
8aCuF3z3N29sYBomHE+aNxK1h6XKIUFFdioK+yn+g8BphXqY1xUj7ky+stKoxtXv
W7eag2Aruy0Lji9aDzp4/nKlKrh6dcjD2qm+wOahjPBnb/KIiXT/vJz0bAWw8zOI
mI+e91d0i8yO8NWSLcGjSH7fZm4ZLw8pbUclOg54EMQJ3W+1uMHxVVf7jzl7wY5G
UmheuCjmzmXIW5zObhp2yKPiH0Vj4Sy43YpMNWaRRV6xPBQP4phK1nJHY+Yu9aHC
+wAT0r+y2OfaSthKFGsphKr6ly0zfGD3G+8FoGZX2jSlTeIqD+D1iWnu77v7yN60
nGlGuyErVYhqpFXwZreqcqfQ37/xk1qCuJCxjkqpTEqxSTZdZB9ocJ4sMCeP+khD
SEMXHoEIMMhTQtXr1iOjL7XavMQ8v7XHBG2uy9DrYyj+n4yIUXYJQIlcc9MDs+av
vBsc6bUgry7RshrZLBmrsJbQD7zHg2mmNi4G+dDVYADrKEL+mEjbiVPQA6hGH3+d
PUCEKBEfK25SrLXeDEUN1l+KBaARMsJbFVebYyrEK+HeIwmMOq550kV8z5cvRAvW
u9Rom54D3+VNgC+RBVvRx5uQR3FuY1CAwpKpYdXt5HVIKMgaj7TceBxZ+HWXdq9l
I1nOpO4ZHUXIQDopbG3Dzj2dctLAiyOv/QqChPRe0fb50GQhnjsxAkf3aLbfqum5
b5YeiLtPa/9RQR4+TN+3B2C+HqpXIh95AVz6Tzr7NSSW7JGP7YM6947ChEh7w5Hi
EHNrIWWSZ5pU0XIsQCM7/5bWVpxegSwpfXZ5Q0kV86DAncs8wBWYls5NBohqTa1E
aNI+2loazJU45uUiU3yFJug7QLKVPqf5P0bZN7/7OCOUIieJ3GJ2sOde+P5Lwa9L
Vk30larkL/Nre4l63eMlpD52cIz5tFVeRt5sM0aI1czBy6K5tYd/wyP7GbJjq5DN
hv/ZQstfckKggkoGiJmFPLD+F0nWi+UHf7R/O+dINAM7j4+0P5fvkZTWBAhG+HHZ
IgihWt6Fw+ygK9GLr56Wkadxdirh5KzQLAb5GdmhnYRgLrj+StPPB5jvvGmtTdDz
P0B/K6p4iOv8VPpivqc8Aa5yGhYUR1g0NOW6tJ9Z8O2a21r4/q8gWALHjHMhr3Z0
LM5NAcAuPtW1M30pNNDFPw6QPvUaFciYT33dgB5Ki0u3VwO/TEVA8Y9gi/KYXbY3
l2RsiEl4boaRReVrkdkHmxk7BMyzh/t2pLxRLNoI3Hu9hJMj+Z9oRebWki+NxHSI
ENLL+9A87oClp3iMn0fe4DPdZ/De/sDMQgprBeyP+Tb2jOmqqTQb7k0nJTRb2pik
t5Bf1HNjLg0bLkAu6ShgJxjM8+4lzENvpnISmA6yiDH+gSOcruyPXh+ywxztW2vB
efqqvQ78EjcGhWCRminCjDTIm6bcZdiBZ5aS1lVBQbDQ9x18I62r8FNQLQrjWfX1
WOV6HJLexzPwCUT29pDsm8THmr1+n7nWdior0FAEugrcz0OpoNg3/W80XDfZMRAI
Aogg1s69OIeKYFe0bai3Jli5jocDVSsGjeXBoa0QcE3eR4vNQITQoyQIU1AS20IV
3Uur9MabqrW9IP+VlL/vi5jvz381xK/bh8o6KMITgctnvQ7sh8Om75Iql/U6dajc
DV+Z8GmoQ6Qgd5gU4ue5LRC2m4OrtO6GfXWWYkmTrOTxCzOPLxGd2jI769yHtwr3
yXGALHQz3ZD99wDO+XNESay6WHJcTilGYYzXzGmfv/LPQr/mBIUDx1TLa8UDeGUt
WjDJVmiJvblHszU+U6Yr7BY389Blwn2JETMnW/rBvW5OjLMUpyu7Z5b7pIBg8RJe
ZUy+67eM+GTOLLSXoY00UKqvNc+ABfvN+qctgLmaLvTUkNE7DBT992nUloIBbRHQ
m4KaQ9yMzDzlGjGD7lyDCa7EEPpR6wP3s3PfVjOYb5/s3RgBrc/Be/v+hAxvwyz/
b2WQ9u0dM5Guk5ciUWPBqK/QL6b1rljvGvZZ9LYhAB4Mg6bR5F3Vu6Etn9hgHozd
5ESo6KJb63G1SL1t06xLXKex/4YTiqKOYtPYHERwbrMJSLDV28iDSF+Xmr3lz9rc
UIxCCfGOZuYt368LMzEWsNPKzhIe5BuiXX/Q/m6g+0eMtWF1JMDSaiP/UWr5qoM6
BlfZT6x/qkd6GYOxuF0No5kM2KO67bHV7Bta0GfvPcoAc7w5onua4zrzh8uqx471
sBgpSV6mPLFCpEF/iyBTpEdTkdimofeqmOhemMi30oPPGMcYRArChQa9ZWf53eLB
d3jp0NnRNLVG0RccWqrH8eOu7Nv9EC/fJzFCpzuO9p7gY4EQLkEjUlbYSTR/Hu/M
o9ObIe/lu+9nsc7+1A8Gj0HOoZxyu2ElIt+970DTRytWPWAPVDB5aYyN1snfk4jg
besNygJsqrxjF9VVa5Xyg+6xRO4rKJ7IARooGTAW2onBUf7Ei8lZttJ58MucivZY
w3Emw0tW31Vtgdo+ixwJN8yDt0CukTaQ9/ocmZva9PPUff0mXbq+xKveVlXyxMgR
xjsy5W9yKXWx+rnWnEm1SqmpDRx14fdlc1SQUE0hcGw+W6OBeuvaOfBoLJPJMoLu
0S7ERT0MC3quQeP1BLTK/0YDBUnPMTGa4NGFg7UcDZeXWb+ZyVfkVIb0C4v2PToU
TI88icJ+g3oyD3xwFt8MrDgN2SQs6wmV1T8yn1ce8CK6CYt8SxJvbnBAji8t5B6x
t8GCFNPc/Qb2s2Apka5yV+07jRD5ICLBv04/uo1kHJBVzts71DMX/LpMghqajQvq
UenApOu43RQtdxdQ+NZslw==
`pragma protect end_protected
