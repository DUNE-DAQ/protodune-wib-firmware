// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:55 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
syi0pYZzjMiuO8eBVnluvxuDWvvUoL2GozjZIO4EKVSRwQVI0LKcjDHr5CzoFaGN
+TnA7BYgyoCf+/8IJVdiecPYezC2U9tQ9z2cWyLaa+qMSlRm8lSVGOwht2mMlCgR
29yZdn5Z5KQGnYPOUDoZJ6Uzc2InwMGQ6US0Tl5VPhc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
euoZCcjJ+Z5IqOslGW3fNTD2yIUJ2nvn+tqM/uGMpCDRGWZJc984B14MZKfJG+Bf
G9ECI6DxdtcjbEy0WZ9knK9gDn1IwAzUKugwf4e67wd3DoQ641BoaMgFOzPAtobr
kDctk9a4OKvFF+ZIgfgIRYw155yRQGyj6med+0SQLB1KT54kHJR1dIwfjC3zdEH8
ADe4NBnlNSqrJILomLmoQViwjMA/XqV+wjwrH7MgYNkB0YaPbsB+ngzRXqvO9bZw
oekj0dd2YM2ThIUVIjYsn8PC13cZzft+ljNUVQiyKk1eNF6VAeMD8XKEQCNAs4do
HY+owtjc82sR1teyJCNFhXGvIAqSwuOEIWd0waZTGdyF+KrzbkgVht33iuGBCNVe
zxGKm4RZdcP9aAf9JyA4W5JQrjKByzBhVEUy4MK4nUv1T9lcDRRNAznzh+saVnQ/
vmJk+RSNZsjxv6KPlEG3lk6CgNy4xqM5QRc064i0ur4G+ZiS6xi0Rt3of7J87Fsj
SoBI4Unl2yJIUK78s1vxvTUcuZihsWk7ygOzt5lc+1kVct1UIvN6BRGZylJ5gnJQ
4OLsviEnabeS+NHBIlsNJ/HEUliZdQAQSg2+ZEhc7v64/njG0pFfobUJsSxwkW0h
fAtCRwVktTAhlB7V/EBMUBKo8BOWTO26jojDDjlS7rqxSF1CZ2M0ouTFRtBf1a9z
C+EQfkzSjUDSZ29z8RG0J3cffA6rsaXdiqgiGO4Mh2De45goLof6tR5ey/OaKuFV
9y3dzyE0/0FS3+AGC4M+6/05NsSB0EzsD5UWi+FAP6cUSZKb4WsqWxQ39d2x5gVv
mKF4LNY/kNMpqJXDDY70XTlMDfXnZnAkwhbsqaLZS9JwH1scwPeRfeM0MRKA84RD
dceAR/bhQooSS3FA99i1TrL2+QhyezaA3utNcOrP8wqHdVU1tjg8UQWc7rnYXulP
d1PQb1HEgxVMMAUCNj+0abkOjSHjAsQM6q9sxrwnjl36sVkUBtcunA/Nn/NtO52P
ndrZF4opjf7LDytfDoCduW2Sh1nK+fjp+++OkDbpXACy/g9SRkk/xnBlDs+9blUt
PJoHBq6RbkADWch4PlwvdqjNpJKsOc6B8tB4CfT2koHLNSOCGovkdZ/AC6+M4VVb
IKOK23lSdKLz1/ZLoL0sOSpvqm2HZbZPoVyhrw3mZHhl/a1Rkp7N+uYk7cyyUfFn
TNyggioyEo8v6AqLhDbBoLWesjJWcT0CQQa3mb2ZOvaRRmgUPYhx/shcZP2OXOzO
5B4bWqIP6iQ2ABhD/ZClK8tOojAP7tJxYiDon7yWkHIwrsZHPVvrpZ2TGhI9T60s
d7WFk+oKjMaD4xGgI0E8YIFTkrhQsRidRKs6M90h7mREtV7KTedr9hOqud0M2oVC
ELKJwugcvRJFyT5CE4bR66N3YXYqCS1c/X0MLN0OQSnVuh0e5RmpYmrebBwPTkXs
3W09RqZ0rJ46svjC/e8OEUqDHNDyFjnFvIb6hBbRnMtv7NDfSCSTxn0PUFmQ3bYy
j9HVeEb2fSkGXr6gVSqs3+RycG8Zu8mDVPzIpl3jqWVGNO6M3KdG2ya9azU4StQ6
YBGAR0A9aUHlpYAARdiW7BVkqiP800HCOuuV1XvGQ6ZGnSsbxmJjsZu7VGZK1hHE
gqkX7TALmn6u4H4gEyYPRuVR9jsHyZhBNfyi0oM5gk+nWAuM7ZQoyElbIiQCwM53
2KFAH/UmZ1NtMvk9KUc0iHdMhRAlb9fwyhy5vauaFu2r9HKPBka53zlARJzl+3YL
OEdCNZBi2wJJWMaWC8gUvN4iLn5XOa1mHx8rQzE3LxwvGfYzRaD6mJuoZOUUyzHL
FJqDOkSod4JcC59kfbIzBdVuqofaJEEsLniWmuYmCExxgpunkZ0DFps1coAMo9Xg
1NHV6EkJYTrdz4Y4jdMnjEptnf5FwuRJRO3u0BNJhghMl96YFFDnGlSzf6t5F8ii
44cmn3uNn0S6+i39Xcm5fDJDJovdxGVua8u0sSHHQzOSJS6GTL1CGMxw+XGfZhGQ
XQrNGVjPTyJguwtRrmkkMmVoiDnImG4QYe1VlbLRH6qK2lUw2bQsxOtMZwfFW3lp
ttIjN0eRxDRgrYmqcj3x5RvJRijLjBMMWKW5lux5wZqOm40+XcBi1byl62pZgO8U
r5UcdtUN9ArMaiiRxhQ3AiAgZb9zUH0vPSgbV5APFwCau/9sdNHdpRvg+2XRI8UH
gCiIREwk2H/as/lRWFK6FBNMUUj0HKgQQC7Fp+vGIZKcp6arXfd6TG32Ow0163e0
bpDqBs55lzIpR1pd2HNsA6XcvP3uspC3/hxf3A06/f6lzTFrTIJFgXJFIkvfl0px
eHZQcbmWo+zxxjMjDm0GyrR08BnZq7KDNs6SgEN1CWlLryzbNreDZfmpIN8NONXJ
6TN3Cjze59Q8P+5imS/e4oHlNfpCeMbydlgAq3ZR5EGw6NtfkQfolSQpKBKA2rLz
AZJGmN0seSvUvv5sTcUmSBwY3ngZtVp5ZodTYMi2zwGvl3r4V5pV7k5aUfy9ohXN
pHM8aEnt+MMD3cViMeiusyke7jiFdTxs9+8bW6aEmQBG0Zqur2avUFC4iAgBOBVZ
he42xQXlhOase/NmqJKnzhTThIvImxxZROWLlj/FdHB20hSlXRzI5fdVXXSihU3v
1NazHTlMK6Lj7k0mviZqtkyGNASdu6ARf7/t7oSnqytFYEtk2a4T9BWO8q1fF7lC
7CCTdbbyvjqMGQr8S8YiA8V9ic/Fsjz/FckxM1mDhd0Bg60IBOJscKyK8lCZpjWz
i9Yjo7tUnxwgOP842zqjXsFZUt6U+xFJrpyL5fNAcOG2MmV87QZqDV0q3qS6mohy
NRfZ4ewtUqlpoSs6STioosZr4uT7Mmw2PWfNXdfqLiui44H7i/zSu9+2XjXS2mAw
A5Uq9Z6DSfeNLl6ZiUv+8dIynbdrwS4FB0J1LLaOB9KrlK3xfHMS3skEjd7eGIJF
0Qih0nViwNL8+ZPZqEiagtdG+cdpMM/ZRZjX13hcghjd8CAwg1TLEfD7EH3SXLyb
bsJGo805ZzLE4+pS142cI1Ii+RtfxQfs5EXxw5TzrI8UpZhisD4TLIHh1HUlLMK5
NS05K9vsR/5rbOwB5T2mHVs07SCQ2Q9ndaD6RO729qJBoHsadn8FmhocxJXay5rQ
jEacg9dRtcqvQoWsKfSB/Y+wMfV+jjEv2hN0ZJhXS3ajnYwKrfoo6ZMIpCSd7oNP
zRYWjytGnRMfLttFW1DGqGeCKIrtaJ4j3GGTLh2zA1lKvos3oGIw/1E4q8/4zUTE
i+YesAKWBA8jwn1eM+bKws1eOFMwh5WqpJcBjXXALpN8acC93tMFPIIZssqBczJ9
812GMyfxkVfat1MJ7kL2VoJuFmrehNRLH5w2sijQ9bUrj6CCHfjWMVymg1MnorTU
ZAzq9t30A0H7MtuIXKn/1BYUJW5fUN2zKJnYk4u7+Gl/CY8gnTuDqxSsZnFfaJgB
oAdaVT4vCZBysy7wKg7ycEOBnovk2AIS49/0HHj9lvmhS0NkxDbfQNCnDyf90lkf
m9Cq7CIP9bqPWyoMgyRfMUMvIAQw6dLov3FsS+ks5BXOJ4BbjXnRL8W0sGOEMLOr
yH9VIj1N52H2f0Uo07BEl7jyCaOszsVDhLM9LXCOZ3zvQaInk1z/MXk0xeLzb0Xk
L5wPm9cG5xOED2dR2twR/k3xV8Soa3jppt7dXLyLww1FyDtUmEDvY9DHLx5F/bOa
d6mVb9a8L8oAUGPjjBQg+kVX5dV00f2BNO6Pl5ZCncwgmiSZpShQIdp0Il3Vj29a
H5ACzZYnDWoTRTIfvxnZ/2Iwzssbljz8dPCJGOxmG7NvZPGsgj5/YCz1bELXf0IV
hamj/0q8rxYcdeAQbBQ9Q/qBPDFOg23A+VK1knrWoftnpfzUpvwksOEP4GeCBuLH
KpgTpDpSvm6daFPxXmFZL9L7VIlgYtrmpmxNy7b+hG97k2YGoBgbD17KI+WUS8e1
adxW2iOWnom944t0nD62lnZh/bGDyPxt+bqt1U9JjPNUuJVkLuaI219HmwMdCbFG
0KCcKaRTOW/HB1q+1l9VE6qoRYv5I25OyeNW+YiaDmzxa2/i8Umqt6GgISIUs6j1
cq6q+Yzyw5Ktz/IA26Y8iFssg0DJ+eKyYPDJhuL2gBYm3d0lCsA5VDi/AZObmebS
51sBq5lcjL00YYrJBRibFcVYWZ+JQpLEOfdNVQWMkVUTTnjN8mWZ7GAXU3CuCVsM
2P/Dmt5XP4GFUNdi/O+8Tb5Vo0Vxx3uqekfG9f8KWjhm/A4aclGagQOajmBG5aZt
4vgxIBgnLHhNbEupnG+VUVhJJ1B+mIfAjSbkNrHjc3cQ13As+zXRel2fJcsV3O2/
vJmMhaoCQ3/Z4RqeXesK4z+bnHug6MDVDL8Nc/WHYUktshpz2ztAM3OVGMBFlpWE
OoLUVVEXO04L30eAsTkl4QDs1kBB90x4mgwKrsrVXTyo1OnWc+p+TcVoYBFtwtSR
ovKCWTaUcywNb0yXdJObgIFUhvZ8vgJVwhCGpE6bXrxVc0WeuaFe1QvkV9A/hOTS
+Z0DiCg2rOmVbGuUYnUokmo0oJjPV/bB79GJeFblN/2oFy/M6mh4rdfd0xJtZMtO
H6lTMiV3AE8yQQn4AAyKo0B62N3t14di7SzdFji6vhuxYQFUxpnkd7TTfZBT+0J3
Xv2dVtEqz2TXqJfym4HXwtBT9pO3jezTUMIqqcv2VqPSDjofPwW9Jw+KdzyUu/gs
muQklhsrctuA4Np4my0uYDs5dWETNhngj4GVGE3bdTfO9IuMXGO7Bh4w+NLkx9Ca
AHH8XKfBMvLo++/LBE2Cvz36tiU5OlJVnJ0d22Of6ZnTZQGBiDvwcItr5wWdztmD
PI91xHr42Aue6DO0EGUxhSVFzHmtEwNKZL7AYJBPcfnYIG1LtLc/kxSLUcUVIcXo
59gjl7p7i+MpQDAyq6BobGqtWqeUbgRqKh0SerWSWw3OYQ/uKGUR/OtsBSskeOK6
TuvtzK3WT7L1CMiYCiIyH5+97OVsm0Jsa8E7E3yO+0rCac1U/0Xp8N0iPjE9JzNF
QETh4/RfgUrFQSba/IuQZnJpHURU/Z3c4owHfSXn7NoCu6vVbBjPx+fIcohsj3L6
h0WMyLLbLzKbiyiuLAGd9RG8ETT6rfMy/1iEoK1o/mBSggpyX2s3pTiLeP1/Ve36
w0jOCGXKquTR+UCIHo7zx9kMPd8djt1+HJRf3V79Yyh1+RTiUjKbYgjCUf9lRJ1w
Yg/2Wtx/w4vP/AbUMcRyVEx/P4CChYWW0f8M0j5gKNoq5j1bOP5C0c3SNnw0FW6w
lHfYhUH15iCdmMD4Zbjv9Tud9S3Vi/4uOhwwvyOab27iyIA3HzQra7eG9gJLIxrk
Ho5igYtDRi3IHTfe5JIqz+c22RUxRWzzSPTp3GkVyBDsN5W0ju2gG7PvkwvMuMp8
7VJssHRpPCeam9QiVOm7T2BYp5RsGCfGNh0C/UeaVcvx30SWt79WH+wU724Pw0um
LEEjySnDhiHXDTbhacqz9uVGTey/XrWhQ/qtYaEX+C8PatNAA15XvZj522VLwy5y
qJHYklYmrzoMIPczC4foWLW012alyP83FWUwE0fBmDgb2cVVHnH6HiMbii0uBP5i
BdN37eKWvmaMwyUa1ArPglf3ZZluI0HOG0JK1TlB5BlAVeuG9xZ2GzSsMN0WiIDD
dZNVKSWW6iFva/Dqispjd/R2grO8+jZ2zKYKj+wjptofr8WEfxrp5XK6NN8CybgV
d/bMQVYlNLN1iF+7dyt/yxzrPpxTx0kodBzQvuDQb12+Oui7CFUxw2JtsISf0y10
nBTy7hqdsi8A6TzgLUVGxq+0RC5sn1G844IsLJQJKfPay8PGYEGzLa2guBBF4Wjm
qedz6yiq9y6IWyjtZEcXn36v0uIH3yLGHe9ya8O+Sg12zehQ9DMtD3QDmyXniJG2
Q3gzV6xaRVe1TuPA4w1poGRsRTb0ASgVW0lbRggrGu7QvDTVDrdrc8Gk37MZnAwg
Wg3B08PSYPEfQ2d0BPBlG+YWuYTi+vlf0CmpMwL4m/l89QtTmvwLSoO4WkmymIab
WCJOmJLeTmxeqRO+ftQTbu7bMF1q2z/AuBeFSzZLF/kME6YAO80bHx4RdvwnbmGi
kR3PD2ym8BE8pgYmEZ75x1VyWLULmL+Rtu2oBLM5NcEPgezcNQx752scZ2QajZnd
pCfYNGOO4dXxF8VHjtykq0rlzoaQhOcScHV6IbpIOIWpiARRHTyUyyILwhQ1HaPG
XaxkUVQrw3KDBuc52imy7AEEpKwsvTcYfYc9uZg5qCLLvZ458bmfr60yVwlYbTHd
ccQiOl/GSa6hWYQ/1PDpIALEnWsr6H7oBt5Ca9sNi/T3g2p13JATdSnRcvv+T79t
mJIMy9vCLtHJv2Q5P+ebjnWnRC+sTrgSoepemapdqCjFObfEZp37tp5whar1cBti
38qe/i1ji5oKPzCL4ENaUBCjkbWW8hAzPQqNW9o9QwScbNmfsVaT5F0QMmbRe3xf
YRQlvB6KQrGemEcUuhdCwSfMD3bMWFY7b/9iS27Lh/HFpserNQfF5mRF39DqC/z7
CnsCjvNO/OsraBuG3ZXUfb618HvsPoZ9Usc2m07HwfvzRoZ+BfpYeq1XtyFTkwhL
btCuPkfJHMwjWRkaWZtZHywSNSXbnYRog9e97m2/gpRUze+7Pgv0Id8QvtrSB+06
6QUE+wS7hvBl9b3diRBxZz722FV1nMWXUv4/ONPCNGxxyNWWJF0EiaDWS13hw4Zd
0dkibYv7bGzVI15A1+a0QMzlgo+FMe2LCFvU1fw7P4AQlq2sIwQg0mXw5GGlvR61
J/lVv6xOmh6RmkvVwX025EJcrUigD5pzMxR9cbYCDQbafMvzW+OpzHmd2TKWQ/On
hjjHl29nnZG3UDnRbAcmKHSnAANHMQhx8w989z2J5R4ZdEGpqvd6VEWIxB7Somu3
l++Ocr1sYorL1+8Oq0GVo5G5Py6alKHTbdYQdzorQDyARalILfKQ+lJqUCEQgPye
Fl5LncT3zZWcLfKF/69kDL2zCnrpt6uPJu80n8smpvuqhP2UibHK1Dks/3ENi8vd
2E/A7dWptXmQ/2spqU6qU3eV3qC4/tML3z5F/2J0qFgi7zuEMabCrGJzZgcRktgS
wh49Fi2Bg8Y8HtjXfNnSJnn3a97DhrWPJ06kF0Jzs+4E581iRBtGIO65EWI7cQkx
Yw/Y8lF9c6BYiQ8ICQnVWjOwPSGa5eW/t+Lj9NBrFq0dJprXYRG1cqr557dXuRai
9JKFU0AX9jtjzmUpzPtA3+nxB5M6wgduGRPh3c22CzhB7+O3hvCEpHflYzMJYQyh
eUPNv0R+/m7bsgOfww8cXmlaX274HpCinnvJJxM3DOPn23xcEJXTzwt8p/B1vuXK
66lgAWfuuPXit+OnkisX+dVXjJk1DO24kpES3al3vL7rXmVEFyzWwRo1hearSard
`pragma protect end_protected
