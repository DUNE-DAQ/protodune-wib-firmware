// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lYW/taVKANa2Bi1pfVvhxkmS0ItNhaENGkjZ5OOS6qiYgvuS8OkNhFXvExtLAHjf
uqmX4O7H8+iMFoyopySSTRgxjB/wJmfGOrvI/Mg6AOxFD2nXIetup/fhi8OXn4mQ
/SZ5dTvXoyhWUZ7R568JFNIgdGdcXJZm/jScF3I32pA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
Fw+6tFOtZR+h/IaZbtlV0JSRLAGXaWxmFoNDFe64sK+hdP/hu37fX4JwM2myhE7M
JNouJvLDIpI/GZTPW6M6RQCgi4+BCI785JkyRpbxZO2NKiPYqcyIX04ftfOn1k1A
BQzIPDAnquTi3V7ISHVPuWsvC7Tz4cl4Ksy6fg+Yl8+RSCaORGrvYiZnd/TP9Px1
jrI4JD9gFnJm8JcKXC/6R6YSIWluM/gxCGJbYjijZ4FsqS0XZBrW2eaoODoOWDSK
kZwS78CqwbcQjM5QhQ4FOm2EwA3/6wu96IWn9KO/PE0RrDCHTZWmKmyjHFVxEkdP
HVYc0Q5B6jzjnANAHdfWSpmtZv/zgdssNVVaD4Sd92Vseyb+bLGB7lnqRoYDVGnt
/qr2ZlrtBs7NG/B/mr31jY3gj4R2EQ7GjZy7qmwIVJK+kURnlEUHRfxFyFbLMwpb
YSFDm0MMuqCHq6xvz5yiWzDPn2rlZ00xf61OorAWWFNmH9aPwCYBCt7z8Ly4uApW
kYSK7hGwmQwnnXKfzilfFuXQzDO0/6nqKGcj/MNpg04uhbIb7lQhwVTGfxkrnfcb
DFEXhYo40Gj9EEviGxCyyzJpSbTPr6QHnn4TEg5aPJzMV0ZbUqpzMc52bOQWNqs+
P+AnKpQGyVSsfSF7h+ki+qqEMOUOwcwOXPUAvQzPNeO4EuXI2S8xPO6R4B0sN993
s8yz+ScyEa5jKeiYhRpNa1UaPISuDpGHHndvjZfLZgU1HGdTJtWjA39orbI6T2iY
fh5XrjpEKJfJ6Jhyb+7YG9lKTg9urnyoPedBvTASW3kkGhDc4Iig1R3kpGpFgbc5
y0OG4juonlBsTdMuQZZRqK6G3xsfYqZ/DTjtXOTOfBIB/2UYMVu+axKDOj/BbA/d
mBxGY+Kz7tpyeiUUskfkw6t5rtBv68t5qpUfCpbLA4BG2OGD+Schfl02NwydVDG9
WiSNqr/J8wJSCSRwZNCx/cGt/Aoo3OiU+vPndHvit+8+C9vSZ7y3fB9qVG3UIhVs
UA0Rq4a8TMb9sdK3QpaRsOIXkiu3boEly5IH8y9qqo6IeFV2JO+9SSTokfNsJpTZ
n/bR3Njd1F9YI5+m5Fyv9z2G4d2Mjycv+FH1fvI41fbJ3y65mVRBjBuIYsUnYdgx
TT/I6rO40jPosNJyimf+SG1w9L+qAaNziofHX/MdYgWxkCffEqs+koGtjkaLYs+z
oahG2OIYss/Y4rM1POMONSFZ3EV/ZQcCIfVwFGwFow5MeH3F1JdkmcrnpGYc3khk
wENaYIZP7XjCSa+LChWaVXXxeS6nTROoUNAzCedQsG2lpl+0r84ncxyu9Tbc0vJo
uMJcYa4bnQj3Z9Y9mTOrSDU8oFnGqJP351m8ufFnRo7QFfJKovuZR41eL3wWs2Vn
k/WoNtaic1wSAmlx+eerI4OwQXIsa0VEO1kxm3h5yOUNoFztIO/lnyyjmHitXcl8
54up7L4dDp0bwOFlPoKHN+qUMOuqbezepkPfdVzLqwExoCN0wcNr5ZtSoUHlPNmr
kVtoMZ0ZOQDZwidHz4USLTKBN+ihuCafUPhmeMKZnMoNMbH1U+neHqULYR54UQ8Z
kwQA9PGie7RyQBaHGjiEcKkQ/mXrkCcF02ccbp8JMmFNL4QWrm5buVjXFyGPkLhl
ipb2j1KZsa/kOn1Yg+anUEYfB5oEmGLspm0n0w7SmiiFob5hQAwA0vGrTEhOas2Z
3UUJJ7VXouLvM6vRMpSSKJBsOCAbca246N5OGS7hWpGeiEicRiQNskcaeIDzOsZQ
QxTV5qvi9LgUJouCvdaIlLupHwh5AxHKXh+YDtdbAq+xXL8dgPY/VS+TNXp0/hL9
Kl4vNyta3oZAcHVls6o057tZNGLYIHo86lVwdEJn+OATWR9UukLfhpiqXSPNPtSv
EnaN0itFHhfn9kMkXuJtjJFMbB+xkDzdKmzYmGW7vOMiuKVet+Rl8T37lzhznOcJ
KmFb7Ds82BkZwTLKaYZ4ghmcPzlQsNgSgZ6/ujUGjwScXo9kf/JAaKrozd1xo3zk
nVIGCjxwYzqMKVD+xxZZn6PtDgsdBXffDTK2HxpvMSl3OOtTTCeWvY4kp0wO8iQH
Ekqc2mhvFc9ZFTGTqLtU/0jRVw1skOZIG/cG6daen1l58yZiwhjn7laCR2GGn7Yp
CfkFkhmiDlMO80b0oZ8/uNvl9o2du2Vrn3fA3pJeqEzn1LfVCM1hNBs1dw1wVpXn
QHsw/QrrcWwmYtvyGoUWw+NNw60bIbEU00ExDyTUYhDTp1Fg6L3bw+6UtIVPtYMx
ERsipgu0ZK/+6BMAbKlcn4lO56P2iuPeabGbcBPkbEXnAAvKjD4hqL6BYmP77XY1
B3u3sqhueZK5NfzlEC5kbUWF6idjeiXCfSDgB7DA3elYvd+C3I2Y/XCFtYA5i8lQ
K3mTgwYxa5QtXxn8QQ20BwHPL+OWK6nsJAIEjjfTZAvtHgJapD7i6aYpwdLKmvgk
NWjX3wmlNrtpw6z/SiidiJWb9RUIkvdTOh+o13KMzJBPq0H3VQVkO8ItFRJXZ+TL
ebtHgtANn283m+lKz0gatkKjPByPs8/3AEnTLOA8iNwaw1e4FP1UautwhXMYYl/l
rqE2M0upRLku2nXy37IkR3S4rabkeJMVkgOqen1iqDenddo5f6thfYuiMtP6WEzz
vWvAArfGWKvrzHXkexAYvsiEfkK4JXeDhNf8Le7pkTmVb6VJJfoOH1/nC4tRO71a
EMlppzW04gZ2BlHTXKBLbg34Xb0uUiOgPxXXGxPYunZaqQG9sAzAoVM+4R2uBrWG
1f/y9ce7IUz9xedAR++xwNqcXHxheuxrTxukxQLh0lRsc7KoTpsEhEZmzlHokdpG
8JMQWdAEj+u81ogYwqalbN0xAirbYs+h7rxaUTYg+4N5rRQCZssNXx8eAdRggqot
affzYmkaLIgkdioc8Xg4XNZ59ne7ZNvj9UU1+Hp2YtBzm4zTdaxIL7qxB1U+TeA5
aRC096l9lWkHU/qqqAyz0wypUZpqQ2KOSfhCQ6wVbifrUY/6FL9LdQRjzSAo//ma
3YlDVeiIFrjHxolpxUujcCNnztxyER/Qn0NBzM/nbwH9d0FGfYuPg2Mg8LmH6+xh
Kf+Avdlf28rrOikWT6FzidHNtGtNw4wYypsZj9ttQAq10hEOa2RFYCnVyFSomP6/
YYd8S/oRWihnJ+CeLG+4avQDSKUUeezbOp55aVA06fxKNpGGwW7aBHY1TAS7b1A+
Jik29h/9wg8jMztBfq2sCnJHTFxWMAzSEj3MqsJY10isg5VDwUtc5npPJSZhwEEG
ncGQ2DarwlFxnBoxy/i6wQiDWntULk0AJNjrgFwwJXhJxpMhu7cmlF02s3IuMqjH
Z3g5NWp3gbR2QKj+YmrP5TJaXd8EXzuflGlU+n3Nmh25B9tRtz9zowOgBZ8zy+O6
lywe5h4b16xAKYESdS7ixEGHWoYz/AoyPyhBfyrAo4N3IieP0wg0JEmiQ3H5BDwT
1IWzAp8o9Bl2CMb+qsH8WE/RfaSySTj30sNla8IIITdvR/QTVweX28j0sjPhkASA
sIcYqMJzJfxYCSEypBiGDSVO2+SVvG+R6W9BC+bxEmmdEr4qCVJPGEBC0fP4otMq
z+T3cGc90dLzcqgUxfWLq/cczWfWxyqiy0UKZKqSSimljj+aQJEMBaHEH06iCIaT
R/RPpYHW/r5M/ooMr/V2sCQ8jQaDOk741Ebb4vEhGdgDRfrvKea0u2K3gHox6+bR
QaEIoKQ3q056Bdp+SWbZWKTVPZCKG8/iG3AtgAcWAVA+47I2Adu/wAAn4cnerGus
Hs0CTiLjnq7aFmSkkBOW3b3qZkh6NwHyzyriWoXyTFmn1lUxxgQrorYv0ex/2Qv/
PJa8FzsdybXDn7Eg0Dmuppb9U8xZRyXXInxsiKRdTlB0dFUH6NUkf9D8Bi7C3LhK
a08e1L4pTsPQPOgT+NOxBIbovJVvmDgb7kVR/6mvro3xmN5bIXyIxlkm0CpfSs3X
FyYnVmWDy6MjvZ8EIow3etEjFlAbVUHfL5VX4ZYjXzOZgxqE3CYU10QdyiHMesk7
yZG7zrcpFJj8Liho1acJoWGTm+WIDlDNkJrd42Anbm0JVtwFLvc2wH+TqCfVS23/
Rgz8dyD03wDhytg0/t9j3MqTShgOdNmwN0EN+TUkuTF0EMerVJkIzkom39b/AQtm
5lrYKP4mF/aRb9h93iP4J+A7a+rEwPb+3axR8B2eYbV6y9l9iMg61HLTWydu+HIV
gcnaksz4Sdv5Ib3GHwzKf8k9kVWrqiKJkFKZgCc1jNWAmG5OVdK0WOcEnrWSXhUQ
+gOJD8UtTT2NnEKXVTZ/IlJ8QMbTVBwWvXLB47Gs/xrqdUoDV95Tyn2I7yARWbod
6706UVwNvIQBahVfsYc9mBuIgV6AkcVsjlClFEy5+ZK6rv4WCSyz0zA89kB3X6mI
dakabrTsVTpkckQtjhf3onFoB5t5q7uW1iAgFO4CekuVKfY4SfOaAda9ULX4J2/o
+a2POzKSx9uhsQn7RcGx+5vmazz12dhoqAdBO0Z5Yhj9hUmMc3B+AAmM9narcFxp
rxKObIQi9yAdeswIOyTx71ZvCxs/908KxhBJFfcqU31eaGIuKCye1yE8Bj4QQ3lk
0zGb66ih8Cayfri68eig3VhVrZKh5Vv1MK5qxcP295/fIc6O7dmHWzbmtV3BnyY9
1rFvVN88+eeAvUSa6hkRfTqZ2QSdiWWPgjq9huYvcpUP91P/8zD4TM7t67bZHPtL
lz35TpOvPAdVAWNF/9XUKCCRvQMKJXCi4MZkWDqPFZ5TTJHtlprk/Ao9V/vgjfQH
tPDVMKODo3mkA9Yas03R+hXiy0nCZ0afZwg0ukYxbqk4HeUfsczgWm9s2a4ZVDIq
cYgpqOybHybtgkLpDzwnYu2mCp/SLU2woHHuT8JXiLn6Wi0+hDINUXvIQX/L5hB8
UEqCX5jYZG2aIKu57duEdEJJNoXwbJl6ILdBuztP60fQlugSAK1nraNfjrnnWDIg
6bf9MjQ7gvbqK7aMn4jftPVjocXTzLE809+PU8H5IAhK6iXcKyOIF7xLL6B1qgYX
AWUn02NjzJUZ8/4EgFGRCv/Lx0PVJH2SWVnTHlL6KP7h3fG2TYJ4CxJC4p407i0D
80ssao8Hr9XWUtih/TzWn91F0n5bm7zRm8Nc5g4RpnzTOx7G/iAGhYypuPeZ7UPI
939Z1vWxKVOqpCW6qgZIigbCM20JUahNswpPqKnZ5xpikoFwYTNe9cMiLblNUVMG
vJp4guhm9WmOHbXZmlhr1pImDM0XHV7e5e7npfqy2yLjy/EazUXUUvB/tAsJgWEk
zY+jw953/UhyFro31NIhu9hMKD70c2vA4TUWN1LVazeTX2YHWZIjHQflyrwuR+IP
h9x/FXCYwf2F0pKRDsmlisxwBxd9gSXl/O5Iig2vSqHcSCNGRGzqeiNJzM0osS9O
c05ryqmohBa+XRJpdO9fCp/RctD2/qyWkmlmmdb4usrbL0p5KSqTNq+7WVV6DT9f
W0GvYDY8ad0cSt3DkRjFAGPYDQYT9ZHYnBznUjPjQcQVBNND6MfM/HrX4y3oNa4t
DbdHqNo3WdbMQWgbAu3Fspps5GcK6aSiqsYeMoKv+RhkR9e2TOTFan8eIrJTTl9k
kLn9iPk9yfF00EcZcbyXI5j4mTxK1FLlPrapw4wt4gKlxd6tK/UlbSlgVn1Xi00e
Pfrb6LoPTiAyIQmrhbjOBn9nbBQ1Tg66NBO+HyYkIyRmaRjTZT68S4qSZsLtWPmp
d1QiRV2Y1TAQxC1cRWzhYjogDHaN4QvJK+9umMvmOIPy/Js3PXSIOI3XQPXSkPT/
InPSjWM/15SsU3Gwlhxdi9VNipFAlADrT79eIg80OejWAHK39k795k6AgTzh2Jxo
5LAskQLhS/vBG2uv34TorL/PBE6scmQONDxswSGz/Fl0s2jgQh1jXgE9cU1+bMFM
iMiceBuygQPfCCkdG09q+HNrScu2oBhUJMcZQWU1w+klneABWuBf70mIC7v5YV8W
E+f4CKr+W7ZnBhbB410gEA0+Dy/GE3EvLnhRssD6+EveE8XjHyGSVjGeovtPlrEv
5Wm+7ol7lLZdMbEQDls8a6SNF04xbGfxScNAW8By4RF4ap4ZwdGjwSxc7kJ2p1t3
5nGT6+BC9Bzwh77ZVcSnR3gIAR9ZxeLiO34Osq0NYQyf9MGyfyZWUvgxaVrNKfdk
UDS5C09bOOlt7NPYGGhDo0qNLLDdhx1xdSe+QpMaW6Lc8YnXAGFvnTAIPnfWI5na
2Av7i/QgmeT3nBT2dXtoIe7oNjSdqs7Un9tjhxzw+ZB3XWIGE9+gQo9TRCFCCnoy
jFZ3ca5M+dbP3rgTgq53hiCuBnpmW/ZFqyjA3DIR9YBcWtVM/8AL/umVT0xrt111
oeshM58xZcfCeGvttaFrPdN4KdSK6tY10wJ2nGqWnkKG+P7BtsOLv7BsxysgNaK5
oJ6wj8pzvKrsmH2urTjFSvQvil9um/8h9iQN9O3NnTSuvQoKyoDA2+3sTZb6ERba
5i86JK3ddNwNSQ3fg5ceNKPuUkvxdSX7yl6ydS9O2DRVVxAjiPRJLrdqW+/XCG7e
ZZzaxCxgKrN8DAk1K3v/HjGe1NNV3hIAGHVadkhPJ8pGrsWjcoA9rW2mubPVEeUW
q3Zeryo81pAhT8HsxCKKlHp5VPUNnxp5eTdB0WtB751EQ0epInx4Ag+tHkoHra/x
ANRTftrHJ1WmC9PMzw3X8PVkwz9W9VuGHuyFZB7et6QNA2T8qpGEbUsNvl06nNv2
dxaNWqFVm05hsVS2jeStSN62oUpO+XJsC6i1kVZ2ATp/T6d0MpfiEiIH526VFBH1
PyqshHWOnKdDWYYT93sa737NxYffebkjGvb+CiFhEVHQvQrS8brURvs1UIQ7eFBA
KEPibomRxUifmkiHq6b42NIdITAdBwJS0zzbPCbFFftE3cGQOshODEoRYxF+AIyO
HJUckMWsPlJZUtKxT/pwzSUyfdJZ+aofmvMuw2peHPgORwVRbrALChUpHbqnEmil
eMOzLMqQDhy6/+ggO8Fo0YZVDQGXoGGukmxYYV/B4GNNRPruQ0ufFaKtkOs02KnZ
74QaE17JRLZ00cT9vIz7g1XdoQx6OmqqO3G3QkzYRO+shKq61hrZte/mSEGhNOry
rlX6uVFaNAAii+dl3vqznV7803TUxYn9eD7Nja6qKCGlV1u9riFgcARuHkJWiQwf
DQrl7aMZwTipHc8w3FCnvTXV4Y3v1GnjhWwYL88DEUJz91GDs8fpkFL09CbCwsmV
TTWmHoULsR+OWB7k5yikaZJgMpyhtA1e+33GI2cp3y0FVZSDwgZmhGUKjHKeutar
S65ZChJjgjfRllKqEE58nttVa94wLffIsxvOThQDaFrZ+2RNsPjFqdA0nppG7zm6
c0Tm6DL0Ll1apc5F32vvgZpppL6LYL2zJ2jOecS/C9MofhBA0E0MWpxo0rWGvkeD
zXeiKSVuXI2SJKH/JahGESU5zm9Uh+mFfjSB9ClWBSpbRmzuYts7AmgVvsyIiQ8X
5NhGdUOVsgLVpzWHk0gZjC/Coerkt4NMaVjozWpZYfBimxskOws+RAlpkUJUQd8k
TJrzA9FmbJQTIATlVVal3I77RNSd360jAR9+2kAcZrNjBbLaLbvscsxyFLS0rhod
BV/aiovx8R9h2LxnyM17zD9OR00daQw2Lww5ILMHiHAklI1mxLAnNsA0ZgkyOhCu
7Db8LIjSBj7jjPixBpZL+bgxX4Tc8QEjDOFlOFSuN9OLjQnLXrMEPro1iOaOcKYX
HN3mEOcPK4/iZM8fiPRp2QEBd4dbqgnJRtB8a0whsO8Vv1jfhofqgZ9M3uoUYmWa
W7km2wqZitmQOsNf9vn5D14qcfg2O4t6okkzQ6OCTGSnZMUxenYj6YXFRrkvbaqY
Yy/zBS6qgc97gkdSDHzCixWG6C49MlAorpH1lz7qI70f3pa1doqQOoof5psFA4vx
z9Nquv7xUfnRHdSEIgfVWjDpFuLWxBtFEtm529q+Z8nJ5iQ61KtGXvFS9qds+1Bp
h9NwTaJzSkmZT6oRMbxVk2fhhQA5zfSnR2GFWZoA6eylFnjBwz8nKKSJmfP5IjWp
4lknB5mzlR872f99vwZdVkcEoOfkEjSXEVL9uQpwvjrcVy0UF9BWbfJhrAsvSEOj
dUJ+Vd21APZRfi8Hu9nZfRXzdRoqwOhgmKTirr9mb48yNJwhD1zaIf0GRlRd+MnU
9+TLL55eEwX7io+GDs0Ohzo2wTUWAsgFjbrTLMq8H+JNF+v9cBmp2sh8169K1fkD
mu74vpJDX7aHIhRd0pQ4uVNvGUH11RzfKTXmRBHkdQFa+su4CR6NwBRpQF/jeL3A
gMLjFYJtFq0kEHO89mKDHYRwhxwB4u388Hphge+J0p25qw1eg0zGid7QhFnjbrFu
tS6YEpk86n7QiWjKMDapiVuLfZDgr+8qCC3cqjAf598Y3pVicOVzM1TPnrAMHtUq
QxFGOm01GfyLaam9jd05A9/4n5lZjX4irmmtTGRlue2uHqgTkJ0/iXHZ3fapT9Dt
up59j8scWdiHWdZdp2PyqnJjOFcofC/jDEwGNO8gsG44jdQ+DEisdV/kk5B27FZ7
ZfLnymiEY3hJfvSCSW3aogvVPr/wFRlFWev0BnhQDew1TtVO7vrZGz0jMpDYZbBr
9B+VpTZ8oSscZ7us6TN7Y43D9qAGXqyqB927jJGauzbCg0VotVbv+Czu3cTgMHly
Pn5XGhgFesqRyP0GlWoFPiyLQKzwmAx3H2an7eXDctk704Me3gF8DA6U7D8oPR4g
XWUTmKYALr7vK217lBOlH9FUYB2jK5OPQSfBZCoERqbiLUJa9wUqeyYDLJ7ufvU3
78Uf+5cua9Wgqvqbuk5rZeEKfmnjzNR9hoA7OnYkZ5hvzcyqmTU9i0ItuDOl521x
nten+RBfsyis+LK4rzUMgH8YsZ48bAzOMgDzoWfgZFYU9UDef5w37hPAYW8mkj78
QI2NvshD8zXUhBVD0xNZloJhNs628zLCfeodygiZZ0JS+ZurZM0UqUCaxXUbAK4E
0pm4p9XKjIBH+ydFBaW8kP2/swTbKU63Ai+qvYGmZNIzPe2Bf/YX89h9DsB59tCd
tSj8chAseAb9locdqi15tHTUF4oTHaqU7BYhuPSbJtSSBYfc0/Hik8L/Ep8u+sqj
HlX3Alk5o/GdUAIemqQVG9tkM8/gTr1BhvqZ2OQoyasHZvi2VLvV74pyl81Lb0ui
9GJwR/qfj45uHWq+iov4MKNco2AlyxEjy007kyKHAtHLvIbzx6ABo180xxPo/7T5
bwMi49MNp8G+I8uFeKXzZlT1tqSeMYSxQPL6ZZIN+uZVawxj9Qf80vs+mFdnM2nr
saMECeqeI1MnuBDnm/XYHY3p9eRwf0G2BuzCbhGXJm3M3aFR3n/sn+ICMb7FRq7t
c3i/OMDvphdDVM2nrvKUPf4UVRUfgndFr51pGlZ/ukpQx29yLm873xflpX0ifNU6
KPfLDs+musA6wAlVBBfqK6KEokACUDnTt5294GU3HMJwHl9SnlN8OSx0yR6V3ZfG
7rVjGTES3fqkFf10lmRT5mo+eDaeP3zJUt8qp92BqjRd4tYHm/pOVj3pcND6OF3y
xmQcPJUCS98ygmMC37J0Z+w1dXl0JOxnZ12tctNH7tEc2Qo+X6hjB0Vrx/lA8ogv
wye6L6iw3YWWiUMrLd+mtY5ceQIMy7tytM2RI7OjUd1iMX8kBX7Nxj4/suYhrbJZ
HmKBEAqwkDjhQuuYMgJmQqlxX2X7MFJ/+s0sbvlhK0/7FrJprjY1Cmcs9YHJWf67
i0jgitFGQg6FpAPhodFD9HFrF5ZwW8sclgPmsHYUunU1zYtv0TLKvRWSAcRhgkEB
8CATtmlAkFPVc0vPOPAhaPn/74LOoLj3KSYMv+J8AuDGirMXKgy7Oa05KC34A6VC
Qb1koONRF++fcdAuY0aHKiz1kfktl64ZGxcirwOljgUbbs62scl7WqcF46WGpwS5
sNb7D20np3ld0nMfqD8LQQ94RP8iiskdyOTi4UyODvG5ZMrnX3JbD/v2W0jtgmZW
1tRQlOieySoeru6eM5NC+O3514nloKfkeYAnSMD4hCoE1jbuY9hUE0qCRLqqenxv
Y0OWmv9+o8OPFjqDZ1SdI7rPwnG/XaxuEK73MTM5HOFDP4hOyn68aukbKeqopEbt
/OirIzkD9ieL83TQQuNSgxmwmxNca/fjPZ8N/GGUVT85e7h1aCBAff3tvRE9H0C4
xY2Tr3MEJ204WJUziAMYD3KJ6qOtNXZm6v6GoNCYNpoXf6Pyfsy+z5mwwuxCPXjK
cZ1wZAYDyE7mhfEpdjQduJ6LPLd8mlIpu+kCWW8yd6pJIH/jZb89cGbyxuzvQBGr
mn7CtNJuEzQmBBil66CLwRWXBtbz4GQ6pLfQofjzdijpCh2W5I/AFQ/dmr2C1Ph+
F/FdCDYFxChKp64SY6vOyKUVXpX8fBYUkM0b1l8nytHepo+ZbxKaAEhyPLFcsErG
579pdqD8M+lwcrI3LoWFd39VYbz3naydVBlcywZh4ufe2oLvMMLcwPlgxrjlkKcJ
kpq4M/lp+5uL9rEGwAdf+2R1y+OqsXeSyI/w31Pk9XwlGx+zUAUFsuzsucONyck0
c+27IuYclSYtB/hw7SstxHiUF63LCpXfUrzHD88zhapAPSUtHciPeC0xbF2VHHyD
RMdbD+4DkgYn0dOcCBOsZXL6oVcISiW6NzZi7525uttlrroposFM55KERu+yIPdj
/it3ZZPjEPEvpU+yhaZEgwY5bsx4HwrbIhQZ2EdhqLhBPNeQmT68ZWtIFg9KCZVm
L3S9+LXT1pKX848RHhMltNbSMDUjZKSnOWl7xjL8HhlmBq/CgkIUls2F5vS1dPPD
fLptOqmVl2IBQHjNRISY9c8V7k2CU9yzqFBjVbxlM6csXPDBgtZygma96R6L8oaq
0Kdi3wedbHF6QcRWhiA0P8cQKq6YssjKB9w6AabYfCn+C5Q+E5JHP+KI97TMiK+X
EPFfx4EUrSI63kMSVVD84888jmeH3NzA3q2briLf5oIrCOuDagbotfodqgkt9V3j
PwCAsXn6bgddC8k4LhSQ5y67MJSxZ8owEzfNp0glxvgbWPVOCpDi3isng+6LQWxt
yrLFjHmOlZqHS6uUtNrXbhXK3wlhqBzMGrTeO9WJX5THn6NtQ0OB5GYjmymYCa0J
u9KBsYq2hdlTSdGzzNwxC0SnvZvYgKVxD3scexIo9r2upGPTZgMShVZIQ73ydaAX
QFpiA1w9lP5Uo/xnU7GtYzCCf1gpCl9WWInoyo7dbbU7nZ1d4gQ4r4dfTH5KC5ae
kQgKdr8aZrnP267KR1VdQ2JvHR0Y2DTpugj5godgS3hWHkWdNx48KiOmGG/h7X1T
92jBOXZ0r/7nVxtBJUGb1UWqtW2CE7cvEHhxJDdEeS2FFcXqASRS4I5ygR3dSzWR
HnM0hQZ7J4sPmyfzWvtr/GP5buvgr7JH7SObtfX3lB3fgAGRP3KUv2GQDg4trKid
YjQIHFKsLh/++4XTsJ6ROMVDsV4/M8R6MaJq+Gh6v0rw1zFqH2SBIbvKgFn4hmjU
9RNi6BsXBXIUopkoxKEsyHoSxgQXpqwRSANp2aZ+iIDqNouK8Wk9eLw5ScXOFe9h
563IE0PY/njDyTbrcEvJD7uuiQRoa/CNRoWVS3a+1VLCWH+W35Qtws5XG+UtOJaD
m7OLDYAgYYyauT3ewVgUM+56pTm9pgDNqiAFBgnsloysQmHqM43qSB8/CUJSe9jq
XarqGcOJ0vb+qF0HgjYvFUBpCqERb9fRoV9VqMqL52KOZN6qe0k+OHUR61qsXTDP
678uCsS5bpwwydq/OJK+tkf9gbziYs0/0WqtO9w3wHtT7x7IaEGWF0W4Qs0aImh5
pqa8E+lPjuhgzCk8d71dC64fxbovwQ/efgTLtuxJg/MSlm8c1otCGxg2847xLS2O
m33IsSV3E1pESY2ONLrYiJa9sC3PAjCfljxYp7Guo4O5IwwvUjcBMvKYROHGSGrF
ARh6OS4qcXlKsxMMqe3B335eGoh50KsErat6MQj7vw8Q5M48PkKXCRf8xtl94ben
4LFabO9tPS0v9x4xwIpkQ4A0o1H1hLacSdT//QkrkevN3wxHEwEGLXDDTZCi5h2f
7nupAWc1lL2aXQEu05JtiJqP78tHdORJmmOPxXm8VFOdVshooSSbdkU7Q67wbMQ7
8BOO3lxQ5C8nhgBrLRxXRfGOCJOWDT7H424xkjyKBy63NYHXyrF3XYeERt548CjR
LQgFehULJN0yDQSJcDqckBGvHizNcFt26F7oidE4evZuZpNqItwfjTVGZOGIvNRp
grM7KaPKas8SKqK+8IdJpx/AngIjR8RxlwecG3uAoRNWfOB6J6KbmIKF0AeB/btS
N/7LDSo7OUNGYStUQ9VvW30pYcAuKJ4kn/cDTT1HVy9WucICjeMVDE47DLL1+DVv
6FOaMnWQZ4MFBE4K5hYr0UBJvqWL7bPT4QJP+Y3yWfeUvL8nlH9rh2bl1sA7WVFF
CnUZ9qZwjBCQv1o4ZC9UA3dD5sNzGmXu8CAxRHQmTZ8TWzn7BgjoSvrxsggbxHRn
S0WdznHr75hN7fo9qvjcwCdaY4NY9UnMCRY1Gbfn9o0OPVnUbTmKtXftVfk65eog
+r63i9RdQN0KCKLw1IDiYPYfKHn3MUYeu57S16xgCWbKuybF1ycRSNgDnwGtS1Up
B4wx+KN0efsEkbIlPeeGLMkXSsYxQYnGAVOyZ7ZL2dWxydwyS+aMtYoFX6gkND2Q
BlghjhSNhx5qX4w9SJ7QGUojhYNTrPdmWaLXtl+Vt3KXEMA2JGy8l1YOgyf5bULO
zSpH9Cr9u4r8YsIfUXEW0UK0jcVwWHid8sB1IToRIaHi7WeDY3zAhEC7rjpmuVWv
m4GCw9tE13cNqlkkIKBvPUuEGf6xp9enTMC9M+ACoShafvEmoGXD4gAMeCZz+ImY
Bn2Bf2FAbvUACf2ImTrw3zfuaMZrEDNf5T1Ed5PHvU+FeI493X6W74tR1rWPEcV2
hlMYlme4xfTeuxJnn6RoD6nOgbboBMHr6srFt+sLpPWGZzGwOmHaEXa7ZwpthfFx
eG/N4kA19BZrKP+nDAsT3APY1Sg53bkkx1+cGLGZvHCVC8+sGBBr9vjhJuDNS0qY
nlMNu2milmUSKgEglDZMW5YiroQwLNFowkSvWOiNSCIBAg43KRhu3N9t6KvfG4HA
8bnxwDjonTi1NxTP+SGNtg6lTIODy81USqPz63SyEVEDT05WoIIl2wxgdSoIMkrH
G9CgzmAyOBnI93MygY1JPy+cFdRcIeeY2YeJlu5IF9HJCQ6xHx5gh3ueqtEfvrDB
yPWes2PezJ2VUMHURfGnS+0pJRGx1HDN6A2EZUEmOJrbzrGVJdDmkD/hNSb26KwZ
Oj7bZYXe6xDvy1Yi8tks7CbO6AZfslpE9DdNO7GYPYwGZzlFp0hsCX7Ls87lcRwh
xrhECZz3GJd7CP/jRXJX73WjcmEurxip4YVtLue9zq9wNPMbeQ66DMCbJpdQx0+U
lXpbc5kGJG16YUQ97MyHPK8pHo+bHE7rB64vsAv/8+qwlDdVKHJsG0I/KhhfLunq
z38dfjwFjK4vqNNaUtkQUWQJA3RB4HHvklcAd8V7IFSbc2rAnfYl5HEVEJTjC4ix
hBdQuK6fVhIZcI9wV/dtNFauhmtt8iKrnJmk/G3wPjqJsXCeOR6wg3Z3cTxxE9ZY
CSbKP1oeoBKUyM8jm2CgU6QWurUadACl1WZnv/y2aZ+AZW248tqp7fV8qDp2iEQd
71d3VtltBi2u5tIfUeV8vzvU3FcYZr3jQ1k1Y3VuuPPIVs0NtPK42Bn9V33FSArv
dF0DGpY2HBN0BVXYFxmXDmBVNoRgGtXrAEwB+nj80sUQTqWOUcqAC3OS+Kpj6oHF
U1LVBMWyckzC/r1AuMmA1Z6eofq9YeZrQYQPtfTQ0ST71yBzQntms3vKDpGLv7mQ
VaHviJ9eDQWpmB+SqKMjbpW5uNd3+AYgxt/r7t4dD7dUxW6lPrnOSrG3asDQ2ME4
z322C4rdbD5opsM+AHsk1j+KogwQA69HdR/0TFHlFAp0OTuLA38kWjTuJ9XXolmT
FOPVh3g418/uR6Jpp0Y3yRHMkDay5VYvGZkdb0GJcKaMU6u99+AyI8pGVwJ7fNRM
O/wtKSaxM4vWmKcqoMSdjKIQh9/yemHTWgRJjjDy7/Yk7Eb05OEFp8MPwyp/9WCg
yjsqth5hs41N3Wfs0rGN+MsbSV5WACBrAKOg3al13gz5OVh1YOQ2SR/4O9lJG8T8
SBboM/NDZyCfP1ZExHh0GO5m60InTibsMzfaP/GRz6gsYqFDx9EeiNhQd2drWvqD
OQU4Oxs2trT+d9K+Qvj1FG8geFe66sNUbWRK3gJ/jaw8RUWrBkeyxhBdplNRy0/I
b2NiBWwlp2r2kuR4nk7ReaQfiTTmXg6PJ8ed54//iSdYfXA+Zs24OjVHse7W/Mp5
+s0K4+0xwLZ6m+B/opRs4Wumv/lM/d2oB/6pw4FwFMDjbrBwosa0msqHUQmJW6/O
qTUVqNKU+D2CH/dSmGS/AC37Qxk6I0Hnir1fKZPL3S8zsjJHby4v7Y/pkYiOXsFd
sInHqWSNnjiiVITOHDtLuD3iJhVWAyP97xjpni/TqB8f92LVd8GRCb80GzeRr84q
LtUYfsTyjyEJC8yiqXeeK5LVpnN3kXv0x9I6xYFEB33aWA/6znJBTxZN10m1GidZ
uRdIiLvZfxojoKTBTdePLuK+VtShD7Xk5iceFPW7TmdigF6nCIG+yf1z1+kZ+quu
48Nxi1ZmXQLF76RIyEbpu2LwBwLUmrTlPzgxqac579MtoRBXiwJ0DWzA7XjIjc2X
qDJ7csQVisPCYPAhYoPH/VpK4v0BjhUc1DTMJUM6oWT6L4h3PtR52uDuXKgNkd+a
K7RVisX46oR57jvYfMfByGwcJ5jKQdc7jd2uWkuACzd7fXuyBNpd75uYJEXMHugu
gwXh1KM81/CHDMPR6enpGIVFMlBUbltCBCZVPjc1a5rEfdn47/PfX456Gk9qQP3g
uISZ7ko/y8eaZTvpTr3Ao7xhp5/DopqzQgHcicFbgN5qh4Qvpg4YQ718xrAlfEvP
oCWRGaUmMYy69raHBXfHWwcZrxjiZeTpdYu7dKKMQxoNZ6PgspBQTu9payJrEUg5
s2X1O84eqtFw8UJGGEHbpd/H2+gYcTCKhFkaN5xxS0kkjAdNSh3egUMBO3i4wVcm
deSUPgMOp35/At02Qj0QBuVwx3hfJ8H4heaOHi5qdb1r3cOv4emBWEvLtYWRzunQ
On+xutVXC3JrC0ZWZUHPX3sqsjloXSKOWB316hS/qLwFqIbFv6rcnhxTEioKA9fB
cKA782VtRlPsZD0lizFl2w7+i3S+17kDZxwWS29ZNi0QkkP1z386TbfLCzbV9v+N
k6HESsPaCoIX4qSNvuqEF6ejdPpoiG57Qza80eWAUdSkJdY0zMMXnQf1okLWHjNz
66YrzuWy1Z5sC0PFHI6zjlVsHYge3HLQF0km9h93gIU1GUFhaK4XMZ/lTnVFbhY/
qN18EbWGLlsAL9Nc8JXlQeS36U6b2RZDJS7oUD+hNcvYuBtVCjNXgOdMQaVukyub
cdFyp0UcdV2ZJR2az5uPXENYz6wlsm2XgvI0VeFjJbUyaja8v2o8MBcgq0wKOeka
2R5Z21pBEHknkQAlHIxIPtMQiEwSwoWWYrBQhqqfoUsAndOM/fOc1yCnlg+I0+5x
KoXr9/+BxgqjMTCNTonBRpvq3BNYT9T6qPmFWqeoMpUMdcJ5TohGD1TmXqDU6XGI
dHWMxalNZ3l2bxKbzvqnFvdEOn4ECwbeDCsHbXdlN1x8ad442aO/wUyivrTQuBnu
pI40s/ZtWaVxTm5gB7OYW9doOfgJd/OLv/Y0CRnHB7CinBjpYRZwbqR/jq+z5uFo
M/RwrIGtvr9hfzvontGFiEos7qsNOJC8NMVsiHKLQS9kWX9s8uA3av+N5lfpsSUu
GQBUUE8O2CbfdesX2S+dvG4SdG2S7JV4dti/NOM3FwabnZTXsB9LJcIkpmF9unRq
yF13dAe6BGjj25mLS7AAy675flkJZ53hyJ9mYxs4I+iCBBef8OtE0Yw32xhci25I
lWgDSYm4i1qMDlf6arQXLPc6vynii1vEL8aJN8LTV5eOep+PkmjIpzttWzaWOxWR
yEnQI77GdpzRrgVGGix7EQMzAlf41/VeYWi5Yst3QSqo97qaPN/Iwk1pHnaXoHRE
k+mXwhamz74Aaus6inIZOuvn5mRzPwWtV0lF7q6/P1HKd8g2kom8czvMwBPexK13
Pz8o5Nmx+nNcs7NrHqqzKJ8HyPZ1/W5Umeg37kTobn8zRKYceW0IOjalY8MFPDHh
4fjhAuHBUbf6ndm3FR9ZqdrniP7WxjYsbtfWDVvUo69aca4fdyZ5Wx9mzsgvkk4j
JQAre29PBmzer14z0u+dER20PwJ5DhDlDGhYp9d0MGf3pdGmNobsdCZicmkQpUqD
bKXcbt/GOcHASrWP+keOdrHkm8XKvF21FFCQH37268EJiN2JHU5Fv0CIfQduQ4Re
THVePIu2eT1kx7u1EagYZJRvwjiQ/Jwbn+HMQWsPRf6/rXkTqf9CZ+Zq3yqPxde4
PloG/wOljBeR7ROUGzfkwHfpBLS8nyjkNk4VK5HD0j/gtcDiUMkzNOo18OYH5zIc
3JU2pYu6xRVXCgTPAH5GFUzkCyYlI0M9iZdyFLxpAMOBuVfQyFbw5+SkW8vXBt9z
h5RNZUun6Kxnx1Giqd8KjHfv5w+YzsMZTt5nRKgbgoYIqojFImiAHJTC1+hk3jy9
9aGmFxLFMgs7zlp0LvZ3KLySVBzt4YOorBasDBtpBiIhyUjiVLujH0p4w6qNn9xA
GCghNS6yGIkuUDmBGdY6AZtiQLl4PFk2C95NS/Ym8BRqAXBzUylOg3V50Vph1doj
yyX+xVxuwwpC2ZIHimixNo+JCtRRiOdxaLwAl4mcyqgj2kji9TAWzxqLdm6W0hsF
8w8lFyaG6GOsU6CLioxSqfNqOiqoK0btOrMFy2DTV/QEj6UC3L7FBU6cmr5OB6TH
u8Nq39QGj/nazWCityfCLZYNi+hH3u9SxvZZ90+YP2bJR9mGa0G2qyz7P+TkU5mX
O0MI6WFsOqng1QQ1Djcnl+E7/kxbcs+XWp7QYBI4cO4X1rStrNL4TVjBoU0ry4cb
RnjDGR9mXfiTtWmfq3dS1eBBnHDDjy8YkEQTfuhKHM9QPveUwTseYxntoFdNKYrw
Gdbyn+arzpc69DFwpEQJY9uxg2tN1NLD5QCPZtA19d61glGGLOzUljCHRmC/ZkrU
blVTHJWVQp13dhtjhaoUIUzgNQFHCpJFMZCShY0uBU06+/pXlS3hfpmmUzQX79C7
mAURXNEMZl6DVWbFBcsTJ/lb7aE/81f2NISFdtFdUVEtIb2DWoSpOLAlERpeWYct
S4Zz6zIG6pvAUgcQhS4K2TMPjJN+k/EPPDrzqKkTR9kFCJqagzARoZKmXEpF5PXF
pbEC9yc++3E68o5SZ4NmSGkKUwa8WJlgHyWyeLuvw0FzeYUj9gpDo0Coiu83uyTX
VJF6YwcEBOufUZMYSpJzQ8Ak5E2QDorByOXVQQ1hDN0+qYgDVJrRKVwY10RWLZ8m
+14edNBTtyr05ILkjxfsaKFa1GtUo/rftrIaFA8PWNOBxneh0IDuxpIVV5fKx5K1
eL7RIjKzLTX5Smvd1KFJtK0IyeeDN42aCStbST/hJTqg6UmOb1Ne5xMTWs+fW4sz
RnntbgywXXSNK2K964iUKRbESEcot2vc9o/mQH0NPNICAbVd4pq6gxAW9rLaxoV9
3Z42GU/NSTykm63jE6pjEjcrb1Cdqbz4i1kN2mYxDZf3itbd3BOi6KnYTSGwmEjT
90sOwHCARIpTcfJ2CnbZRHSf7fRo4TDjY8ljh93Ukk+vD6QGr1+xvhPtYaYavgE9
Ya8DB1BT2/kZZZMfDn0O4ue1+JxK7e1JgsowrT68UJTVzZgZSXz7FSoS+NVITbNt
8x+hyeiK7FXO6Pd1A5n3FAeRRVCnz8GXThtxjPhn0GJBSbNEzzcuECxXLZKr9Vhf
FHlUluYegkZ2ICdutBhX5O0ma8CJQUvm3bJctk4jhamj2VFYCR4CJCtHXyGZoBzT
YjpbgbITPNUIAf32RMkKcq7aUO7DexvGQoL1G5Ycon0/FOeM6ch/pAXOMGU/p6NG
10TaeLSD4oEdlZr4h8A5kM8Hf04sUxEGvB5MHEYKiADHy6aoMOpwq4tRlmt8d2tT
H7K6zp8EuH9H1n4/x2wObYF09jrTDEsXRuqwjOV5BtXDvO8JwA4234a1znqjUwnJ
idmaL2hJhovKvsRAxtnYv9c+8MOwdya1pEmk0jkcnxk86ZAZAFFy49/KiMHYL5bL
kqN7hBDmuKCt3PM6WuxU43x2JuiheaW7rmxfvrGV2sIyoirRb9aTpKcefyphyClK
kFKDfwWgUpljnyHkIg1E5lZu+/gbtnKd4vOleZ08GRmb/FMpkXWK3K0l5WhZ3r64
qrA9LA3AlInuIV5BDM5eDpMK2orVmdDLuvuLbVy2/Uyr3szPCDMD/zwjG4VnWgSh
MOO5b58fy3V+nTBLZ7E9TpxhyX90CF3HbdcYEUYt5HbPmeweZNnuxsIvwV2q6n2s
Qg1dM1EP/EolXAORM6ShFz3ywnTRUFy/xZNeNG005SB8eKtNAcJ1pV4ns70+A4lN
ASz25rtzcrA7YgY0VG6vpmODoroQCsIgVj37zXK9nFt6QGirwxqiro8PcNX4xrJ/
yGMckd4FPxtCVFPvCh85cgBUFdTitZS4otJRqAk+JP0JYqIHLvgLqA6rDrt0AkPg
niTmgFln8594iBZxOEU1DR1G0xEsjPT7k4CAlQ2ua75ay37DtG3ScXL5aRXiT7ep
KTB1ygc5I/bc3MzmmcUyMX7dGefWMHFgtCZg25eDNjLIJTR9ckWpi+89e0Lnr3qQ
2A9ZgjWoX/CaaqFsp99T94fwgV2MPJ6kr+B9IRY6Vi0C7SYxb2KlQTa+YJl2XC6u
Bb5hUe2EC7JCG2qQ8QFJpin061iFbT0sDeqW1+HNvTZNKLh/BUafIWllfsMHBBbh
pHLC0V+2RmJMwWqztQpWXa5ztiCLYvmI+AKac++YP5Nz0NUjfOwtZ/8XwSYV7g6/
vYLXi32VNxsTTaE/tNicutiWh2qojdFpTjNCFnWMTy0l+5QQtMXwrTJXB9hr71bq
Db3m+47t4k8goXc/cI+rzbUgpm19W+7OSJctroKCiJu4d3FqjgW3xpByX7StiM23
h0awi28wVvtrq8x2aVdkaCZ4HU7QuJEpIjWl2g+vXXHyvV/YM5cfWwcrQwTEsmgf
R0GXSUgMiL5LpNuCWcfsEdfGYqgjimjTvQyinOi+IM7nsf1iolgeQla/GTilA6Om
n72oEoG6saM9GvGZfgg/bp7ySEK01lNbP4T6/LfvvZtD+GhZYKA7b73ekj+O+eSN
4NAWHm6QKs8Obm3oztMT4F8yxdhzS2M3V+zQDsgYImn2LQY0ZBE7uz+2vvIYjAFk
gseWlEraRp1xDBypc+b0WBdk2RMauLrFOFp8FAlcteaRp1pA04Mr0OXncPlsoytQ
rzLq9v15kIE+/ob04+4V7j1O/YwWhgXpyXhI/BgxJKB9tsvAVke13FRjq2PO8Tpo
L4zdTfQ7sr+EieLJlgDhfGRQVXlqL3kIzst8FBJKpaZiBTup7PaSLhWbslhlrquV
RiK5qcelKIOw8w0QZDN/+xi1J1AjU8/gBNyM830WPZd7ESKqwVOjy8d8ngGf+C9n
7WcUpUvL93dJ6Z4TguugErKAVSn2D7i/zMm4Cdh5+wQwQaVpiD9c0yettNj2rEFA
XQnaI1j6C4aoU6SmYCzKcPt0jKeneLJGexWe7vUlm5FlRB7SGC2ihSfqfOCQ5uKL
gGyhEjbcXKzPEliWfAlqPfKiTNqdSIP0c985JJDPpdMPFlJYQGSgPvPS//bSbAj9
XXhy+aXq7gHT9NA8hW9gTCEQByNLxDpC2pk78sdNMv1uVaCbcQqgAJ+u4dP659Lr
WXbTvSnuM5YcOw0Hw9JAPpNPld/s8sP/1hm/bgUJlruj4PCI+No+seiUq1lq/B0i
KMyoWsX4c4bQon4qB0EjqZ96OXZc73ry63fPJm5p2+9TSI7gjxd+61z9SyvCNmm2
Gy5zobXMdWKvc2IOwNjxdANKSv7CtVo07f0ASq1qoFTe8/wO5pAhVIPsn+x+P8ED
FdZwxjwrV4m0l28UnabqdPHdOgDOr0hz5VkBjIjtUa3E0QQk97TZKxiIy4HLawTf
s9xm64VqCHxM8n3SdTJauqPh6Odt3XzTRJ6ox0DRvpSw7ugFkatOHcE8ZF5Ad0r9
srSXCetqRDYySSvWsdC8FYZlwJdEBy5AkaS5Q/GTmo9VVSWpCRWTTAZtmMYlaIqp
xXbi3RPqBN7cnN5QqCtiSc0KLM1f2VHHHzQ8oWhi2t0PurUHJXjOcb/Og410FaJ5
HP1r01g1H56WiLdxdD2Pg8PdddcKpn7pmFDUeY7M7Z0YZOQY5cnemNJPuJzkIdRG
rDGqn9XkT05602uqyOPpNhjKxP1jrg7oLR98uZIi0dfJa4CV+870vyd3hlF0dLxh
BIMaG+yw6WIO+NtznpESxVPGFPTtyXo85n9ABH5746GPI5k6RzSUYxoq7qMksswr
maWBraBYAo/06z/Y0RVoMgRCkUERT93xvIAcjNyjsw5fuLnyVLx28alBqoigm3rD
9PkNTmBvq5ozL5vJ370n2laZKyCF1J7BadAjkF/MwlNMEtphUP27eEXriHsvC2f8
JB4DYIuSduTBkr/xusOdMIgjWHpLBpic8Rh0wwfFQJ+DQAS7NJ4s5Dl9J4N35wEy
F+VQciZPO3J1eGAVkPHG1bSQq+AVtSKtwz+shnsPAoC3OdKeYjPOtYB99Z11q0ph
2zTHRfdadb8mPF8bGEYGAxZpxgP3z/DuX2kr4DhHEzGtNlYMsa6srwHWqodZSCH4
yQDBFwYOL5aw/OrFmEC4OybAcXNAEiUUPjGTLF4DgY+SpFnMkHoh6SVMMyVF76il
q5MtjK3YIQa+pSol3cO9vVxmf+M3amJPnkck+GdK9iswsHO+Nwe3TW3lyj6d5Iok
MCU2kZkUq8aUHMk5N6KmgueMWcoHjgHqMeBn8Ur4L3Jfbx+wjjkApKR74JWGunNr
3Chzy13BCt6gdUzrcvB5hPv9wi1LK0kZ18R4QhxLZnFAybRFVeTlfw6e5R99djBr
eFhtjNEpPDBXmwqiu0ZCaofY1jFpKl+EPM6E2U2spBiHrtrbKIsJ+L+ZQkbSqB5B
Pz1/Ww/GWbcdMvatY0ZL2snb1d7GqJi2N6oBxE9T3Kn1+kWgZF0+1YGg5QNLDP0C
qlMx6YRXvyzrCwtp+mP63kpkg1CZRT2+yp7U+OWO7rbEzwbmH5vsbbZjNE6vuzky
ljaaeaDu7QGsuQHTB4OooPY0I9kPD/NsxL3UOjAfdpvmfnPZYV7JJCg5elBF5UvG
MQr6scS7WVdPeT92J1wtbhCIkUlmC5U1eeMJzJVS8iOcrIo4OKguPy9cwq9s0I4W
n4OhWuJ7LsfBISnsDEvsQBCUe6b+78ida+URuHmAvmsgpm5Uj8pS/yzNZ0d6p+AO
RZ+qyH9zF0tnd53iPCzIg/zb4clkKRFfEG2LghmCqyUBt5mtEKA7uDWY6gc79T/y
VL/QQqW3W0oMYq9+m9ZGBbqpxIfEF6Cfwj5PFd0DGQ4TsGvjS1P2C3DJck29sSWX
u45qihA+eNxNjXMkcZUXfFvIq6JN8K+t+ogu32AEH0RCE/GLtqssvHaeCppglfkg
UQVfZ7eS5kFNT5Er2UfZwPlY44ICGJ4KyQxCjl7vHSw3ItLvth90PIDAvPeIjKGo
DteSnDAxGcQbdFXX+elNvKvK1UA449zvv7kYwXzdtCYi4wwhzM2I/zc1dRUEp5g8
fqVtxwieQr88WmaV49E0BtSv5+JmiNVfz6L5on164hvfTLhSf7Zt0OwaBdovmEPK
EciVCd55JoLptQL/EYpbJvC8rNXoDUJy9hkRcWWy+vFgEGzwU/pqb+lgCvpM67vw
nT4XTAi9MJ5xiXBnrYJpVoFzqjyt1188ADIqy3INYQeIRCyS+BcUGOIDr/g7yZ/X
wcOTxUWtEPJxwtY2ce3MxUtcRIM4VJPxajNcfa6ld/G77o5OpRxVpm9dFxa+RFLT
fsiJTafui5u0NtluLUaC60atEoWAzc5R7rB6Wgd57ijG5SZUm5K9jBGUJ8qYU2/R
5jhfrkdbkMwSS7Kxg9AonpjghDDmE1eVhhGYut9+xjc7WtVGWSCH0yeyQlHicZ8B
E0MpUtRFSOvynKZdSLt9/GFBdoZDzY8z6BUbYOMlHoxEv2HoeYsl+73JXvHsAmpT
f604BTr3AJYVolCAy7LYUlRbBmBAFFq4VjnkGTYnL2DVptQywn9JHs3HyG9c5V5x
iH05bbdhvI2HC7IrvtldDG6nytpgwEs2ar00r1z7YqRYJx5hSDbRtY4zAiYtgrKw
glEz4YecXCFSfRn+Qx2lA4bY2uX/F5upVP18WDFM85fKYnyZl6tprMg+AMWLWCyf
Lm0aAfYupzJElc9Z8PHyKPR0YlZc8J1QVcE+W4+BGHG4ou4upHEa+jqx+JJfbWEA
EDQaTAa4edQbL8qAHytOUbrQO8vPBYEiL47o2AQfMqqNy/GZs9BmTqhqAUN53mpw
vxVaXz9z7sWmUVpOJ5cgAcZkPPn3oXudjR1l3OeFhkIQmM3KsXQjXf736U1B6dWI
TVz6AlCj+mBVQoZdBFc1QQMn1P6/4TnB6P2TkKgr7ONx8wdBKV4efEPyM/fcJ6gu
5cTtF5UhzFt6TZbrtFqQfMVteheV6MvCgIKpmbxbrF7+ZvMfMzOygUg7v00CQtPM
PZM3uejPpIq5H0l8WUG1lWeufF/lir+fjYYKvtMYlJJw9A5OskIPZJgsUj8lU3fI
9yB2GjkZmKnwu9Q7oDu4YkahnMcz3ZMIhsjE9xK/EOHqbclt76Qv9XatueFVhFbQ
xbPDSdmAkVFFbpoKv5ku+RSkWO8TVn+k1dQcAQ4GW1CQZOEQtPRCW6pj7Rsk4V8w
iVZxzbS7xNjSY8nNR/mIZRa9jeSqP6w6AwVSEbmaJlbrmD96eTf267eiOeSZ9SVU
MlRGs+kMtik0zclrC/y+093blkTJGEzgKPPiINxHinxTs3+qMB2+1loFlZvekBTw
R5lRS8smuLG2OiV5P2K4y16agX1rc4e2KRHj8bJsHBM6tvLz/dsDYnqe9JpC2+qD
PpBEevFRz6gB21g5n1pAB5fm4wTssMPFH7m2oNJHsG/igGsYfKw0CCz4i7gBTmoT
wAs58tzW4681ndKzzLA0L9KtUf7nG7wscJgeHyhCXjpRgK3+IqI7CAcQHb7KWVIB
iJ6g3kaZG8EbzSh2U3dtUfjiv6SPGWjWCo7ARXuHiAaTAFdf4WBS2C/uFLFiX4UN
MBw4EbTiLbXiXofi7gzk72H5OjjC43m1hl0GXaQIbP5wwj3/zcd4A+NdA65AUPV5
z1mwdEEfWet8S1H//986pnBJ+x4tFUsmdLO8XHSgSrZNYtQJB5fEhdVg4DUiO1kh
nTwv7eNsPO//1sas2GzqGGGeqwDGPOzULslf7Yukn29j+7Us0JNKSwBWYto5YNVn
S31HX1Baemeh5OhLe51opnUfEhpv6cSpuSsuWS6TSPlfZwo7emP3Gw7lk8dxPrII
uocs7guij9gzq1/hOygxgGWyld/7C5jNAtYsXpZo2z7qgoNCBcvIxy+3rPVzgl/l
lQUEVLrgrO2R9cCkGh/28wMvHQlh8H1HJHKfB1AGXgIo+oC2sWV15ITqHkUgPR3s
L6pKIIiXL3t1pV6soSi/9gpW4oQ4Lc9RPchhAnAGaLKCLmq1+R+SdvBKkuShD/XP
e/z+PwT2ItF13blQ0lRz9QEjJTGYesZU4bG0K79KT9NI7psS4Yz3LrvFCBENJwEF
pQnIhFRLxTzspNq+H2HxDnGJeS/3qyUxXqG1Z2KMAjapPi2Z/FX28OoGgU3LN6AP
kyF5ENsxozRK0x+rid6uUoTHqJU1hLjRHf3sjA3/pACdD+uQXQb0fuZAAvcTj75O
eTADRbrgbqljCqNhGH25DxL42c3v29pniF3Q6TF2Mihaai5FQPJ5o5MueDn7/5fe
s5KDo2eVlubf39uIbBKumie0sIfpolTxA93J1JRsfWto+Is89VKLB4JWLLHdJ5ta
RikwVkb67/z7xwwzMe2KMnL1CNsD1uSi0gnLMzlazQthstQy18ChM7sWSK8M12/r
jZUx+YQAoHe8I9sEGwGFreUcBShrmvoJHS/ImSWiP5NAg1HzBoyAl5tabDiJx63p
yeE4tlWxv0blzwKAgP52SsgbKaBFOgpHjj4BsPObraZvWX64JV3U68S9IQepn1fc
Wek5FXiqUSstj5W+9zEmDeNc5swjSov4fSNTSAJNN30ErWrmjIpimk2/ZIyDjurU
iy6cEKkLnGVX09s6G4+lFpDs+fc/Ydu28KsTkF1eWNDKdy/ukn46U6Wj+TOdX0C8
q6RfxBC/y7YWO7H5hhjT6ABgXoDIYHNXPp3T4LcsHR1xokq34jGMo2DHZx1k5+gU
qUIDZBiTv/9NFicLR/NdFFJ271Ki1GY7Afo8oM+SQoFd68pfc8Bnrsqs/Z0lgH3q
vWxXCGlZmPYDCaS++9T9+dXB04d2B91YICVrNTa78DBRkMOy6Yi4jU4rMeLQ+77i
pL/V8vMY8NgR2RUkebdObZfOkA+SdQ8n9O6cKpPibPTgNITHGqrExmMFURucpv+F
gX/HZw+ddha5bFOB8QkO8KZu0jMDfJ/4Z6z/4OuoI8Yt63UG011ZCBXWB4yAvkRN
rXHG2JLVvequMUgDy4+ch6cX0J98WRFvdRNj0ZqnZGHHCPt6auhJdELCHUvYCuL7
HrVxg+2HISdCdy3PGM1s0ZftltZV+mGLCgoMyj5yek5j+BVKvr5A8y+qIY5ZfCbL
ociPn8Rhsi1tlS2e5TbVewe9iblofNsO0l7z8sj/oJNYX3OFVCPsFEeqAWarlUA1
tSzarqyxKINc4o9/Fc+1lsEgNzATN9BNx67rIN8Qfa343OE78N+J1vc/9ZNnsc49
kCcCrBFKQjA/gUUPSxPK3kGOyOYu7xFeqOzWUuGvWiu9vHtkvuige5ynHt8+bVHo
Fl2YcZHjR5ZkYNJZey7cuOxAmYo71sEzDFvdamQUfNEs+xd1FEt9enxvOK4LpoHm
aWWxdq+glO5F2Y0IOI4ZJw/Z4aGyZJmEI0y/0X02ykThYy89l5wryW+YQZasfYvc
gS6gOaRfszbXNVZjSxm1EaqQzJSa7YHn4PMVq6amZ0VY1oYyIuQgvjjzwX4BeA0q
/Z+gZifPHKW0cesu4LG6mDWtH9w2eDmXNt+/PG54kvfLi0d0EjV39xmc+dm7tCyw
KPsOhgBC6qOGpoMgiThVK+m5uhHFclkN5JoC1oY28Xxwg5Y/8+kNfbzgybN2dY01
bE+/jobAsdM/+/qlaNlMxbfrR9/ByXyVycQpGZXUijXs0+KFXpjVTuLKKHP2suPp
7/k9wOTK0DRe7M2H0e3qPVt047nJRqR9B8LvZYUka7Ms3jj23MVr+34MvgWZ/T6G
+flMVsnat1FW2iCh8S1qYROEl/VNE3Wpihdbyb/pV+J7mJ1Y8OCLby0BjEif+5Zi
jGspoiPl4TrqmqRVGfSeFV+7mE3DpJrSIwk/oCtD9cXRTUyvADSfKcDJR9A3yktI
YKNPRXYHrDUcnSdM8xLUu91yH4RlD27DU8wm89P8RzThs+++//AGTLHhAHL+ZTfb
jtJ7MC6MFrSmAjsWKiE8j8p3lt2LrlI66KyOcjO6fzc=
`pragma protect end_protected
