// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+2o1j2TDkdxqP3MzD3BhRVYFPRIwn6AJ7HVpdeWGO8BkDYq/w4EqFAxwXtUHZGXB
77AXZ9+QUJ92taig9V3e/GVqA/jepC7RGGe521ZEj5TcRwTbbkqAZhtTmW2RfNP4
FDdYvwjXWOi9zeS8MBkckvwCalfqCSfHNdBUU/ubV53tO045gmby7Q==
//pragma protect end_key_block
//pragma protect digest_block
1snVRRU6CnQpF/zwehDbfB7cbUM=
//pragma protect end_digest_block
//pragma protect data_block
GxmXqKonGmtvHMB97/E4l7twIRTEZCXH4xGTYwZtg6JR3Lu3v2Qvl5qmR+oGguEl
NHyaiRGlpKpZaX3/HqftcnsDcGgYZzOwlSoQ03uHQVIquSrcq0wGWE4e0sWndIxI
sIywyyEShUXeg0tnKnxDwnuddWqyCisegW9NZopHaVXhyYFYJxj/PZTIeY0sU+2a
h3qu1tVGP0RKrP8Bv7mWrQXYTMJH4G1Ta5kwa9s4AyTtMwgvknTtsPLh2r0/yUeG
vQLFc0UVfukSVRpkuEf7GeDiTBpSHp0bbgT55OiPMJRHPSWPupZqGVDn/p87YgBN
7zS/odrM+She9TiHwYjS/PCixRms3zPHyFAU6EGmcX7xgMeWB3rPklxqcN8EzZzq
0JbkiT2P0CdpS+ZtUoElvs4HgVxu1m9KjEk8il8olnU297r5+hjL7OWTwOUNsJvu
K4ZcEeZtSzX3sMyErBUk4a26jC+ALrvs2mdyigtmdL5BxdGNwV4FEAknlQmzhDWZ
5jLRUE1HoO0k7qv5r1YeD5+ZjI77PS/vp4lGH75WQxGzGJCDfy/d+ozv31QM3E4R
l9hBCdwbfbReDU7TgkN48j9SzcTrtGLHqcFOKcJjsEuqnKINFgPVWu79wCWgIn6e
tTHGxnFXwZAj3CwVJnDGb5gE669a1EjASSK1nXzAx/+EI9RjMOkNpGuaGWeKaY9c
COlf9pz7Tg8Sk3qXgXtG+mJP1HX5B9jI/auWLBWPshB5Y3YS6DgR8o8bq628t5+u
bdb4wbaFi+yHFoHsdaAQtPGhE1srXDKtmbk9TP0D2zNuqTmFGIBAd64eY+IcOFBD
xMUvPU32APvr1zfUB/sYeK10EaCQR5DEtGU7QjCnS59t8rAaQFMu/+ioTl5NY/P9
8TzhM6emzwFmGOSrPAzwOBLEPOpXeZ9cO0x3unBavwLYr61PeedIbtqhhZi2zkyy
4D0Mt6lxRhQ+QksDnhmNijjSxVwW110VKmI66NNc+BN1HoHzNZyctjJVUk2alETC
aAxooiCKV3yGUgZffEvwA7Lgck16MO/WyEYNKZsmNgxIVeEQDJ7Lwv0tdGwnIRWf
WYa47Jn3aX9uMiW5bMDldpL3RxzOtSg460Kl07Wyycs+sliJDXrx5CFbXNqZfnyb
r6Rb4Pl0yQ8OynSrXVWtPZhq+zdOyIJwQ1imbDTb8ZJKoFRJwK4nmJhbYfBpYoUI
oao5t1tTWOhxz0ntiClIt7LqaLrycdT78lbyoM4WovKrBBiFyvdiTNXKFBXiuFR2
2xygBukymTDINPcFoAU9Rj6V5+yUija2w9H4U6eOd0ZqAfcn4zVGCVrVeGo7JFkY
NQEv1t7L/oSUn8sleyK1iPMfjZw7Xp09hCzcl51TKJ9tzK82V+1p7d+Cf+LF+Cfy
ejxK4OW7+QknoJU61YryBOA4UwMfeo/LkC/GoihnKzehC9cGEkBOc57cYBCeogJc
dQU1ONrQRT658ecYX0fsIRJ7BDeCmOexRFCF/g6dWfcdL2mVDhv4hxIlL9YaupBZ
h+c46xjozPCe8xPhRer4cnXCHpM5mEp1WYX4cLLZbvV68pqgHnVuSvYCpbU2etr0
pmiCuUXM2WJZ5WcdmIN8+oEjw7g/yVQET73CY6W3alxgy/YA7rn+d/u6wzmShr1L
iOE6Zb3QZ3tZKNnkXCD4DJ+QnHRFgKXE/F0zH1r9VM0gC6grW24O0ooidwRMQuL2
Usbh980XyOoZBBCfQ5vUPFGLDx6cyr29MW/nIwlotIUeQBASdZEwoEJXaCuCtv5m
wPaDxliS8B04scUGsnhanP/4T1VxHTVivR5guFXyZtitdtDAkR8tBGM0wA9oB22E
MZQkuapjaDCgMxCStxSD+cQjhxnRlQ1WZUz/ABITlBDImkgaQ0OG/GtCFaLOK5AG
S56o5GOCs6S+MTVlpn0PZINbzgsdfzQCyj514M8Fa6ngJkntxaSsvT6sk703Lhr4
P4+f652YkuDlAahVzAlIPFOj91IiiIHUM9YphxRFWW9ks9pfms4slnv17M74M9Ux
4dDjh6xDyDa1hu8M56zuVez9/mTkfjks+FifxQ+pSoxSqbk8DAUU7GJ3mBV9hMqE
gT0osSBOSOLZ4BsSZBr4F6SoU6NCkDn5Kzjey2OQhn9LI15FCMxtQqLXZ6nE9rOX
5JezzT552Fm4A8Wtby37Cx0r0JezXVlLtDejWJfNmrrlvr2qzuMOBXoEZNa+VhSd
59f9PA9sAjZoM6DXrE9ZqHHCf7ZM9jluhjqmaGSt1Mvmjw0/d9H+pinCJeRxB30T
bVgV4AvrqyEIhKeeSJRgJg0jEGbMkl38g6mB1JhCQvFmTHKsxYLZp1Nh+97gRM2x
ez4lFAB3Pzp32G+nIkDA0thE9bnKiVwrRgfBLZbclNcHOVs6OZLle6tV9cKglhhv
clkDWlU2I+OhFuoz8t0LvU8p1CwG7x/qnBk9gr1qV4R36kG+SmJAgapuWvxgI6ei
MQyExj/zvG3T21knpXN0u/05ZS8rrGXtHXZ3Sty33a4XfCh5+4lCZwxuXPZRtBQb
z/4Dcqb8a8tFRywgfi33OXNbl6xzdo/AQVs3hhNC/J4cnb7Rh9hYO7+A3WcsDg5M
NZbDQPRLPVPJsCzkiFsV+bzy8/nPq0pe3/s2V3IwFmJQjVJTL9UwK5lB7GhXertS
Qgl0KGeZU+8caJQvEsaDYkk4fUD37VfDV+jZO8qsfGWkLkq4FsGA9spznzCtWkVo
qhnmtsxYT+AF9zWbHGix+hdFe4dred0i9VC21rT6u9SyIls7I4PKOcNOdDB6R2y/
JYObPki5ZCe8uttoyxdzoDOksmw+GxeBFVGb+7SO/69toqOSAohn3YYXhB5+xa+s
qfW3QeK4yzYuCPIvK5kktyrIrVHgfpCfuQNVIRevSasG9XtK54emTcGODMVs/VDT
3i2corwvckr4cDjEtbGoOOjkrgMCilZnqdapBWgQM1hFT8la7htv50Oib/o3DVs+
73Ld1D65kdkg32t17I71/VftXlnI+uKYFI3DntY7pzHKmV4BxsfQikZDbtnSjxY7
ykPoCYHdFHXAh0//xb/9AFuun9djFH+9yLia28vPf/jTFyAQzkWhq7PHpGN9HYlr
b23uvyl4VYB1mCyv+inek0andv117NEd9rmTRuUB6NtAI3jEuO4EO/KuRsBHYpux
W5vfqJP2cWnBDQW9zTsDHCxA3/NMQEOwJmB9VJ58aPkf137xUrT8gX3CJvB1MY2m
K2U6gc1akmsc99HZqqHLwpca6tjDRc5jnBJQRVUvwOZabFu7WYE8vTTfo3dOEyE8
XyKSVXkeZ3dUEJ9xq2OzN8QhnJuW1IkHmkojs+HRj+OFpPEv1lgcLrHQIurB3rZF
3Q8Pt1AMOiE9oxR51+rwg9DVbKshQI3xTnpYg7Y6J9ihKC6vOih/u7SjuEdUS16P
b0Kl2ctcpJqkIc6B6Wzjs4CkZwJ0iFwWlnPCQXBzLxk8XyXrA+iLaw4xOVUVampt
gidt8WypZ4ClLVqfW/Z8LT2SYeW6Q7iCPmVeGtmuGorfV/dFFln8YtpMq/07gZTW
yHBj2srIfOFJlPMfhPa9U/AXdowmRA1GAbODKzxCK0uTZde/RqLMxBXEj7ksUAk7
zU9X4ywTMDt6LnEiJuY6ZahasgiDfab3UvAaJvNhbZsAq3qbCYg64KayzAGvjxd7
CNztFCC/wINY5EbceQn+KI+libUNZVEnLtlNrLq7b2A7aTiI7wh6Kc9Y/2fXVzLy
3LJBn7nbm+bfFVSq7Dl46+VMaunRZ7ORxABXudA/+wLRZRB/2oNUEPDgHUckSkrt
y8vnvYDRLSLvK/i4wBFxq5qrzATZtSjjHYCjwmN1WDNHp3cPdDTv88SQmwLoz+am
eGSESRJVwwTUleo6wTwK8rgajQbVgAO6YNBCL4wa6wFTGlBik5q//5Ab5GFGdFoj
xLE8CsNSKTPuRFyVNVCdbY//uQnrowBDY91AIpS7t7a70sdXCwZI6SaY2PJaV51E
IhwiiMgj9GphbZ41IqMBzeTL1VQD1EJ6jWFk5tBlPQZTwUi8VB7bMDoLc46Eb+Ty
2EYanbKD1Bwhyo3BG67uEVOxtQedmGKvLnHshDhAxeF+uSSc8b4m0Z2fYiRQ62UD
pe1MYAGEfusA/H3Px5ih80UWsXtq7hDMi9G/RzdTa8SKoA84rB+L+ziMp6MV4RlD
Ycz/Ebd1UB/8SnhLaqCwwqLdx51+j7IT13AF1ctWvW/XwU+577Y/0qh3u9PGyT+w
EolaQxLu25nRwwOgu4ZkUcGFtujq+wTvnaF4Khf32e8dccEil097LNyrhBZv7XOc
FHG5hxwQOAeZD/lc3eGCSVE+j2ZpB5m89SEYBABeuWzYdC9VcQVADSqKu94Yf98h
My0vr9DQNexTDVHfkg2nIsgEvrqtXDPBpy7oFcZ3RbDJZfuHcRK2Iix0IBdZJvIB
JDQTCsavAYuDUG/A4rex4SqcYjCgtWwDvvsO26JpoOFRGr0W4Q0Cph12H7fqQDP3
iRCHd7ew9jAG5kNKutdhqZuhaMW1SIkZKlxI4bnRYMp8J3PHER5iqFw/cdOy6naB
N6ryjT8V+u3kC0eL9OhWdKrxvPosmctwSM4ayO25thpIyCZ3wg1IcdZP2Vx3oo+6
YDjyVrDt61knDybKHNOJskbrlEt63RDv43UiZbAlIIBiwPyQY2EnFOy2w65aUl72
zt5IAhJwiPrpviNehvVyGJYuBTTwKWoUMYonvD+y16J8sLqZkNWcgsra/P9MRcBu
Xv9rlH3NPyMk4dNJ188+GWzID6DQ+t0v92FTR/UO85NOuatr2+YSyMUTnHzngpHV
rtJ1o7PZ61xH1D96HoTiUglVAG8eEVk4e1gztx8yAfDHkkeOgTBFLI9jkwWePl5t
GY9sBmWGYLACrLuXytPIqbsCNsltua5sekpmPOqTqz/hghY+O206unLMHHGMwSXV
3ohwBBwmuZa/hCYUaLJpP9Mrr91RBC/5FA6OLXrHcKu+0Y1bbYvdi9G4qyIzuzPJ
3es7h/SJePhbr9dK8PTbqTqKdThkneD2WoWSmJ2Yw+VUQZcwVHOJoEV7MBLlFbEp
OKNYt9BnSLKb/VTUixE4buA8dDLkdwxH+yQLARMXtYJ/q0WVV2367yQ191MMpqQF
JKhGkhwt6Cx+UMr+lehngsF4iml2g2eR7jx3QO05v565PuhCsx4kXw8Cy/rAMceW
gACv2LAOaiZEJyn0APdhlbEhi2Pa5a60oUdJqNuxOzb1oSS/Xm7myXiXBe/V4iIw
d2RqCdc62cit1hu7ok9qwaMhCNbEy4n/NoRo/kdg30/oBgYExJm+GKjNvY52O5G2
ooAVQuXFdY2j5ZrALylLUoF6mB7074m0xC4aL0NzjQLHnQb3LESqHNzAY3+/vBN7
8ar4YNNr6svxfGNl/UdJcu9XTtesZPzlgcjv5hhIQ1R0Ca6IJDKCNfpcURv6jVgt
xPJvt/jAXXf6OOxDCdsydsEFfIeZ5ykwacRrt63olKZmFu+PL6jS2pCNIILl+PXa
h+AcNyqxaTZW63nG8PiOWpM4VYYTJEvEbciWACpJ4f48/ao+Wcxl8FTCztwNVIV5
Zq1imZLVjvHSq6/hvX6BwXn71+FTwQJkxlGLmS6jrr6YKfGuUB06wCNTRXsStPB6
E6Zr4TBm8c/uqmKoTcqjkAqIfoIyMG23Otyeep3/aPP8Pl25Otd49H/JQcu/pLTI
phWm5yNvs67n1yPvb1g4SVbZ1QRJ8pMnDMDpUTSUYFRWTsjcWgKkZgim63qZ/JQr
3wfzaI3FY5UlER7cIbgNTDQd4OZEdpW7nz+X3vqJP1ubJCes2PcQ6jwh8I3hDeke
AGLCYZWCJOumjWUCtdjfl7GBHV2E7LA2AP9NQplNIzwvT2xUau3MPKu4Zrnn8plf
OkpPdlIU698XO2aTsjD7fG5QoYMc4xyd0gj5mCOrIW3F2mTOALXaLICzHYoull+k
BypLLoTf9r8zguP8zDWCuPv4lRJThZmvzblmaN8E2JQm5oy4VqrQXo1XdMlPE4/I
sOk0sxu5fJjKSiovpbH6tC9dOUrOxRKE7bL9jeA9DDZHSzFrXxvooVGoP/f8zEtx
ff+l6cpiB/2iAo04YGDn3UrSALZj4tSStaozDK0DjYPXqalyf132gxgLiQU3jFo7
HjtTEDn1om1FMuO0QxpD78ALfmFkBpH2TUQcMcesmn7NvJdA2hjRf4wRyyAApjTm
ewIwgyrexpiDy0PYBZaBz/QEyK6NRaNTQWHHuBgninl8Qk/8pYGQ2g4wtJh8aOo1
XOVfnee5s4WHz9rbyMvFWhBQhEY+tRVik/NFi1wvWOvQTMRUvRSmRVJVTxtjgevQ
YjLcXAR6kpt32+3hWhlh05Bnlv9bTH3PFyOSZlwtCeN5Wd50mvHgizwF8wMYAluG
5B7UWnYX36XjRGzjHJilmG2k+2Nn94tqtR2dijOxuZQRnFvugQm7r5NYkinGufN1
7cgPvPPIWN9eRfU3ffYSdVfvDXuY9HbG+8qpfQ3vqbSUQWBYmvnTtU+VDUqrdZ4g
tRchFDjL7r/1JJV9H3PN/k/T8U1p8NMPUHWHl9YA/2iKHBZjlY7hBY6O2HgMwnph
dEULAvjA4mr7FnVCWeeDvuDMZWvs6n+K0W2v4Urfn8CwdgD6nCW7RPncn0U3ftwm
m2hQK2geVA55LkxN2qRAwBrOn8i5vwfoAITUk4yGjULk/dpnH+7zgQuDdBn/NsiX
Eznrp9f3ztOPjYIzMWjJZw7VBNuZGd/YZHQvjfaqE1RXWZLzuOFGyLCNGZX/ULl1
4WHnOh2XfeShEAaD+9X39FPcHKOWHD+XrATqPRzw/zryL47ms1hWzYgXcDtFXIaT
ioAoC78hT74ZeMrrBwAbzq46+QgYSbREEydU3igNmKBXmXBNazK3olw+E+SVLcUc
irLcUuFxFFm/Fpgc+YPYhux4jeG1njrtgg/GAFsmRwBcd/MG1ml3622MExpHsmHY
8kgEXFAlTB1wgN4Ydx4oa/eLhZQxp0yOxO7TzobyEHnrnmD3FIXm2JNSlzEwzuLF
8Y+3FptheCRFTrSci/JEYudHlSpIr9K/9BjbvWLFHHQAZex3tHeyy1nZLulyHFjG
aOMRFdufSgs9gHwUYNlwER1+8lZuXmwfCkzSqzXEMLMe6uvBN+Z/W3NH6GLVGvO+
UiRRX2qbDynpNNrcKomEXxeg3abaPqdKHx75UVIHmBHzBdg3tyXGDL6hsKfuBHzN
rCp+p9ULwa7ugL2xer8wp5HntT19arFS3UCyYg1RyUCO4ONTEeP0nvB/tZWQMKXj
zyEhO5B8x2E5vgyh5djEKSL1xhxH0qPCuz01WhErMvGnFumbKmp2SRR/9uMZF/CK
0gWqmy2LUEOsrOu4b/fyXxCphaQugOrPtxpOOHfcVNp9IS3LTL3UHuX+EOxZM+ez
SSzeIjXNdTK24Q/w64uDlzybqw8fVc64xrrTpPkdm0UziqTNK70QvClvo+iPMZXE
hBq9EqDzErZVpI+A4ySsY3WB3JrjzxR/xQnk6M6FtjUzsEPYn6aVEa2q98N/0tfN
R2PFEUxySPpQNQlbObU3RTJlNoT8rj+pc1ob3bmcZRAWtjeH45iafiy9Cagnqjod
kW+muME2HkrwGvNagtYhUWq0uh89MWIIJFE9mgs/E3cG11nfKaM3lkpYpoKJbWuP
Pn2MIi79WMW0iVIrOPnIOIy9dKey6nvYnxiGbFyG04hlSbGjlAaR9zEA8vL11AsI
i9WtM47BroPuuuWZP+BcY5X2xIhsaKmziLf+626z0XD8T4wPAaLSwa/v6Hsym45K
MjIjqEXXykx+y5rqGf9tPbKgPMU2YxfWdlpn68PUZHc4upj/MHFU6EqxmqL0p0NX
C68UvB2+F4bxuqXpybfWjlnWanpfzSvWZzCd0mPFNITz933Skr25lD3SnVlZ6EhO
AX+ZdGkQ5zr3RDy+psHzRoai1a+Qihp2WbBRhFWO9l+jegkwDnw9BdnmkZVWINRT
1th2oB8LIf/iWpQWI1IisYOlOsFaImFhTMBL23/1hDVknUQ6AazQYcKToHfxeU+q
pe4B8N4e708RZpc3Bgb7H2hrq/xeNHwiYmQFoKrgIZCiqCbPAtAiHtUSd/C88st/
XXfEP5r52mylEwEuPywcQPEimffpXw1DXF6s93eGlJzyJsBDSgVv8Asl6UrO3c6s
wCDzL2+J5t61pdDc98ygkYvookoildeDFSW76GKziTs+XpfGByLsxvMgiw3CvknQ
cw9EF89eWdkoevcT5Xu2FN4WWpnfhw0gCICmk4EcOyoVIhM1PJNr6apSbXEfQO91
a7mUJGc1Gff8mmfOlHmgS0SOUvasOkvdn2ushvNKdu5qGrkEKS1X6K36wLtVYbrG
N7BEJAWQGZFqUVZ4qSyxnvifGET+Ui/09gXxO+xZ9cW0bOypPaFl3i/+bZ9ZzFC6
/8aeinEuH15YfzEwCLzTEa/GU/pNo3+mLPB8Pv3wNVhbTlpu6UBCAofL3SJ0HVam
DpmTXIIZyaBvgDXENxhg0//yOJnvDs17DS27NAEIjz+sVGtxjfLWEtpoZzWM4+tA
orjaHk7l9NjFZ6ZPJtxjqT6Z9GM19+ZBO1Cy/o4y4XsQOZbeIGFJ1YsMrjF6aRnF
RW5SXIBzUsa4LzjgOzqfN349hhCoySu8cKemw3nat+ttSFddnjMjMoMG1i/9eeZM
lvkbsGRxGENfH6YoxyCLxdhUtvVD1eMZ65KW6C3KMn15I0drWLHsOeg4BIXKMvyF
Dkk6hxOKz3Td/Q87rwKDDnf2MUBJXHH92nqfodzfzPr7PD/1d8wBuWYnKw+Q+JcR
zu8r4EMMBUBiOTIdQjRkm0B44MqhoNamjm4KamG7Fef+Q9jlvQw8vh5ekogmDb/s
iC5zW7MiD1nbVHTwPjSppYhA8NrTazDXsbGaeMTrJ5gV5ptgOR2O18l9+PnrKAle
U3Dr9Ny1SRG7ye+Vuo6sbziYOXoV1b8WPk//6XYnLEHCzIhRepF71tT/84t+xddI
VwNiOKYccdYmF/CAQPi7Dlk0vD7wg/XqER/tS/QOVPT7L8CnIwjZzvNxoWXVyT/G
c6M1lRfamC2L6VqAF3tiP3pr8RtxCiEwa+PrUPG7gNPP7p8gEWv9A1prTy4AYwMO
JKCt+ojdBIjMI1imnyqJQa8Xm+GvSYZsKG7yhC969Q6O9CSEBysKQQfTLBp1r8qe
Nmu15ECVm+fufgIW5cpZAAS2WSsFz6r2tr5dY1bMv6RShYCh8AteNC8gRgxOQ07S
icHegSesjWe1zOgMihBfU4nsr1RMYTK3q82FruRvHA16O9zCf1Lh1WuoKbW84YZG
1EK+CrxmwX7mugnJSPmyeAw420wtnXXjbb3SSb0HPqiQoNEMHDKbeQtzs2Vvd/LX
XQqgepD9vx4Hl46LneRKqWbFiPif6Yqbvwktv4c6DDX4e3fuwLhr7eDGqXR9GiTC
HOhOqQUvsRStDZIj6R3Jw3XCH9XObC/URjUhv2CgH2YOuoThpsR7q1ZYZJ4wWtij
2CIn8TQ8s7PXt1n1+rIrj4UT2xh4NkLm5N9w3Of0+bxltdZkh7ulY6fdxSF7O4EY
MS4E8EKZMgoQX4OIANOSZYe5n3S9H3/TOzO7xYPUe54mK1p/1wFFHiEhyyLnmPpN
otGJ7VeoBzpos+wiPirCtX99p1viit79vUpJkH4bqfBBk3evaF3UGIsRyp95Esoj
XzET6YMN9WwyLJSXKAOTfa8Xxwu66FdThpMK7nBt8YnNJ8P703DeTKi88LYuqboZ
tMboA/Ty0H7BfIeuwY7NkF5PsfSxY98f+6/mU7aA1ld9PEutAJJFLawvzN+tjFmH
mj0oHD1lj/UG6f/01q7QxyU1AO5hXTnQCzpxdNOUDw5UAnXrzL3YtEFRkXBzXmno
d1Bz5G0QW+pNaXBD3wqaiMGKFxNpVgmJgTmqxYrBQiz3Q+bh5zjVVGVhlj97PFvh
Ncmh3QG5hUZoP1xgqUgGPcnVNXjgpL1QpLcI/xuLLCuHb1vIROB1mWYhbrdCZlaz
vfMECO+uF/3Gy0KYenCFblKY0HGb1P6pWI0t9Pn8l6LBh625dh9bOspd0EOiIol0
wxwtcHOpeZPYq1hXv5EKoK1sTd9y0fYn/Kb5u2rRp5V8tS+xfRjVQ/tZX9tvdLgh
Mk7JSX/X67umBdi7sTxeRQ+ysoDU8cDABRNdaL0J1XurKd+Cnqe848hMycFHuwbG
UClD/b2ayMc+S+pVLGwxAQk0CNg0/e+H8fFx8HUPgKigAH4v1nx9sBs3VTG84c9A
T/26CH6r4+J7G1QkBKB5N1hjD/d73rhdKYsHwEPvXSwy//ZxZBFHkRDujyvrGIxq
srgXhYdKc/MVccBQmivQPSiO+LcALMb2ZRrNDxm1Op5aYEX33tB0PM+aNVB/Gq8S
/EwSdDiVFclikd2QS9Vrmgqn8Y7ZJogyVswPfmzEZXWn/qKsF0DVmoYBzf56UZ77
uyqK7aTESzulTnSWvy8nAjW2q01aJtrogipE9e622RIrGS9Ta6hRje3IAwbel9gH
hzU+y9XNd77hizRZqZVBBfyfySc3tHJhcYRiJ/A6XtVAG1WiXiH7vpCrak2XGg5T
2AEmAKkA2QSaCui+1ZevyuIu+jqNj5YVWbqJQiWwqx9IjsQEnuzeZdezhzza45ba
AB4sMsqOuCT+8dTpxGXuaHo1LLq8rcrVFnfoiAjgX1m0K2AuifGpBg8WlI7qvyxV
XSe0G6vhcmgdY7Tp8VH/6+AdEGv/feJfCKCyg++fjZGfDajOEpfcxcTPMlpG7isi
15tSVTXtF/CRAH1Sp7WWowTqKCPKd+WjrXKD0r+Zsh/hYG36BD3hRcEeV1biTskG
P2QO11ru1w8rTX6jr0f85xgh1bLF7+0Dd926Mi8nuz5vSkjPmO9lvFexJilOmcA9
H5ESrAOQBJTebtP2CLKGc4h2+nealWlXRkJc/+fZnpYIfCCCOfn6a38ZYYZ9q16g
wa3IDw2Gcu77C5KBqK3X+gXEsmUVUG6uqu61j77g3649laP0xgYGPzPa983m4hW1
q7XCNSpmOt8CCwic6uCIpkZv1HPq6P91Q/Sqa82HidpgKDDTS9Kie7sCg/LJ2BTM
3+W5nhN6iOAuhx3Va6hBNFRH3fC4hzuBxb5HqYfhGP4bNXckhnAFcrqTfmzuuv8g
kRbjaMoLZTddfIHWVytsquLZTYi39OlcDfZKYlybRlTySMO3iUjlLG8eo3VDFTW0
jJdYGqs14xHQAebK/zXZjVeX5U5suvuBav7Ei2FFxkavrdnVRPDztkYMOftjlVug
eGhW8UKI7+GOm8cYyPJnI9XE7Hp0k2LpOMae4xbx42hg75N31rsMu8bTwUBlLkRI
xaIfL8RersD3jJwi9fad9wp/C7+iLeOCYtC+Alz9Cp+elPbFdMIguYI4UoTGyL0X
6tiRQVh80S+b8M4wXivOIPSFtRaUrHl34lj52ZCJHFmk8L+gDXE6B/lF83Ym2LbS
foIAQaaNjN/u1C0lVHRPScxfgYWYe4az6Q2hmeSpjAE43QZuvLFAAnlD5vQb873a
AJZJ1B3FsYPuOo4RPoHCy4afJt6Klp2YoaiGA7UikpA6au17pHqb3G8K9BTYEass
PlmTJ8GCpYU6XMXn4Oj6JGUTm+5yPuqwKWpX0qJB3P/3IB6cDB8+VxQRqqyfQ6Uv
Tf+A0lXRKtHE7LhbQpwvziutOTzVhrm0SmCs1XyqhvJs64lEKTNKgtKVW1GhO1dE
8kBT/H2VPya18L8cE7ata1PpvHRHx0HbtmBl8i9WbZHILEsvuwYV1tIpmCenHbzk
TpkPELQI3dCgUPZ2Boar7t+goaZnrTgobKTdjHkbY2mZEdK+fV6wnCtgxBkOZmLc
mkTMMF374x6pw5EVH1zC8vZ7ZWLz3170o5pUJasrSev5CLRrFm8lp3C1J+0k78ko
cby1AGL91ci4ibACzE70iGyDkGCLEb1P/oz6Ll0gVSlANQIbNhogIxBcptJxFco5
k6bvhe3HfGVlhXbo9/CyI24UfatszOVodjRoApbFokq6x5NqKs3iP8lJL2SYMnR3
wn593Lz0sheK4hF3mAvkGqK/WotMiNlGTUIwGRisFAesD7aLyG3Zckoco0Ta/Rkv
r1HXvgb28Tyi13eSm/skv4clrLMsEYftvCShp6oo6RSb7uOpgaBMkEnTqXWhSfVe
L3b2DozA6whVxKxYr9ypsFALFDT6EOuxo+t4UKI90aRqoGSoZ0P3u32Bs6mcmePn
KIKS/IfIWNGVVKtB+D6+XvHx77IfDzk4AwvKzXUboKlgAv7FZ5ZdjSJXtK/3RsHG
JCDlQRvDK6FQWfdbxRF8ELvadXDWwrCJbm+NLOmhLmnEylC5J9i4MG+5NB+GSb2X
pORITKIqYDNdVAoR3sAQiaAuz5AsPyDrsYJTg1xnutW5MJH10kEtnNeYXcW4htW0
a5NSq9Tcm/RmHXwlTpcxQWuAgf0A7FId/ygOIGNRwU8GHrSgzKUGjql6eA3xkcyc
e6u5vmNOKNrxHpITg+ly6LtPhQFAZxY9rbjz52v4mkQSk1Dt7LiPb6YPYh1/JXzh
aMlf1Iv2hTMeApjHqjNQPVgKL1A3jnHm8UTWiy+L7dmi+sGqorcepVvBEWL9eML5
l4bh6BADHnV5Xbxvh0cW3wkiKhxfHtbpVn2R/lndgFjL8WEHccTJWLwLt+6//oLT
f7lHTK+zA/B/JIo9G2wawpAbY5nGlx8+rms+VZCmQTxOiZAI3+xoQKinODanoJ/O
tyVVUGE5MGOUts17JV14zBExclm8T8lxnaifWoaqGx17dW4ZOZFlhJWD0z0bD4Na
fbeqbAslrVCPwD3oz5qZlEvM7Ce646+mQbNzGGGN9z74946Q1HVRrrBJ4bqrSjDw
Q9yl40fullhpFLD/4uqirRAsEqjBG5hqFa0YiQ96lG8t2DXBR/k1pVx1rcVpYuOa
l67SS02+9l0Kht8dubBPZYd9Z43N9eBVoh8nDjIwbOzM4JNwxmvzLZOXR1Fhgp0i
xv3uBDf0l2hA6z5bdUiIz1yEnfHU53/vY/WJE3hkIpobddnvPotXGCGrvl3e1D2t
loI5oDSU8hI6eTZpwwyCp2R2AI6JhyrzUYezcRBkzhZ2lvaMp6cQN5Cp41ViB+mQ
Wnx+wqhDd3P0pROAUutddfsnu+cp0dlNQ/Lh3mGHMN4WnEnc+w1lE3e59zAmA/M0
JV0lK6bg/Ldh26MJQrGp0LntvrmezcfWZ0iR6AJXY9Ix0UAOeJf/nmwanQWVPBkG
VC/LDBqesFKWhmnrTSvVlkiWdV5xMWOz0CJbPtR4hCY+wRhF+4LS1VsnO8BK8N/a
f6CSxkL3yzg2M7HatQrhnFJvoMqGPD9tSCqVhDXAABhLhET1ARPi6GtnhSeriRVi
KK3KE6Ud9p8kUEFv4qIYbzWE9VnQOrt+rcrqysEvnv4kio0TjHaX+0VXDYYPRasS
Uf96t8VeOWr2WKBgCRBTr6vaMFUZv3BNsyRVRfvUHCC5k6g0GLw+321FoI6zVIA9
CWEBj8SW+qEN4hM6dt9ZVuiLKsO31y/lUmWTTTlTuxb6O0HapzVSfqNskd6lk3KS
59geI826I8iSBNkzdqfnOBS6hZZwtYcN3ol0MdvLg9LoQJWW0kzIQ2jPcARC89Qw
ZFFdOQp/VVBlyJmY6Jp3fbdBWLslcSvwpJCsWiXaJBP3/6biIVqnlHbboqBw29yJ
PCleV/+Ah6tLa2LLBIAxRWdSkBJzJdLtJq/3/AWJKNRGeA4djMm2yYig+cHyy/t2
VV3gSsWOIhGBalRqEruemkuH3DEDLMvi1qzC2SSupSmiu08PFnWqP8e9ttb0h39i
LaIpQNWhk4a1gFDPJFSfGdqIIrZkIWUh9RAwegLFJHvj5Pxgs6Q8EZZU4C6W4x0D
oHFmsX5/lVpn3QqZnn3zLZIF//gfDkzhH42iGiocd59NWmpvMLB2Ri7OKWdlqgXh
xX30LwO3GlRqGZ24fbhYCT5ar+pz+yDuThxfBLdrdCqWHhnUToIjnMabce4LinvX
aMI4xv0Lbv8hSpCPBny+QulVAeYYLW7uymk7B7q7QTvJYu8AYlPNvlYWfi+ljM8x
lxoi5H+9BD3aGi56z0CP40EsabU3I6FTGcG13NsMqGjp2NA7IuNxWhr5qYzksQgH
+gXZSSFJ/Rxyhj/qoxLuzcnefMK7tLvuyVf4YSudCtpn1ACtv1RPSJs2wa1Q6goP
0Tsqqq+P+il16W4uNYfHG1U700xCvvdtsbVvyNZI1tgM7/lAJjqdX2wfs40qLocG
ue+F9I0bReqgZJWthGQ38kDWyp8EvGa0f9HlgfKiNaPFVL1mG5uliV1R9t5mOLhh
xkYDKuiG9ZmYiBClcRXbf0/nwqKF+duK9xvRQsAQ0yo1C+zcQH0K8/+xzyW5Fe2E
eRd2661mBFsDBukMRjujPQ==
//pragma protect end_data_block
//pragma protect digest_block
+DHB3U1YqUMjKrZVe/NWYOKSz0A=
//pragma protect end_digest_block
//pragma protect end_protected
