// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i4AwxZnNPFmm2OWfYTh79zjQ7c7lsVx9En6QQSKrtHMpuyEei/CGmSnBkneK4fhQ
a5C3YXM7QJfvIinu7/op2Jg6hIwEJj5vUnI3Lpw9x57OnSADBClPx2pNfDSnfGNa
3LGp3jrI+POXe7zRXTir2FlzAUj7eATcLykwdTLUPD4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22000)
sW6AtKWdRstN8JmbaHSuFV77h39bDdsCxoPMPm8c08YrtA1RbaMeHfzNt258Hd76
lLvMUcALJdCIusThGHu7wvlNnSIQebBXpL2lDXivCA4o/rmZnw1oz0/4OL/ERjff
V0efki4pi5JOZrQ2oiblkbhreiM17KiZ64O1vjljpogdR42hxv9j9yhlThLQtJOD
Cx2I4pcpBOYEpPUp2QioS435nrA2dQunq/C4+htAzcwIPThPn+088vzkOoemv07N
ZEOP24Spui9Gqd1Vs7Y3DcLGi4/6CikBlp/gJPfZuRU7IA+s4R+b0TfGzXqpub/W
dJAZ6qIl9ik29GUkOiRSmDDkOIHhdEzu1ZsfqbdTIRUULBVK0+dgv9JEfNpRdlUz
uzo5RUx3bswwx7q94NDGY+5r/NPn3a6KU0CI5Ns1CwAM/YbaizGua0sfsFACVzup
GFsgvVoQ+R4xpHoZK4DvI7lRxn1k6Nhl89BHWufkQ8s9drfy6zsGvigcoXB+vzAp
EnjhCsxNRpEtjZwzQr+rfDpcREJpoS66+GzgDd/W7vGxZ1K67bBz+Mufdpysr/Tt
5QOODRi37nnO2GA+D5qaJPsywQ5qa9PaPV3fgwVfGSAQty5obpY94Gk7/svO6hFS
fO6XoTBCIO/DpJ17d/is/3hR8BFBxvbXear+45DMs7Y67gCVtj3NgIb0upsxamas
H+eYLi4vSJWn+W/kmnucjmNiX4GsDYIKFlt4k39oo/QERci1DuNYsLXXFImLXuZf
BZ6tfTRFWKdB6zJO/6OTGkfhhnCpdcpX/oICMR5QioPD7G6BDEqGZE5iFZONyCW1
heuaNV8P1gPoGeTYKP4HqNsvGjrLk9wzkLdRNrRsOArNOg4SZtSbk1xyHNuCrQZN
lEt5SCaCeXRslwfG/6dMDOrpI3AAq8+nFDdXxKHsuN1ahJgynCXrjvpuh6oZdVd2
9RKDTCUfGuaa9cD+dD03c/cqVMmFmU7kM+JuBQtjXmqeR6RaX1MFWqB8Blzcrd8u
lG9mi4beRbKphZuC3hDPOz6nSYekofDebYcD+rt9IPFXc4x7pcCi8j91dkKLrLCa
imXqNsbukBDWQ1kSZAzvfxfo/t7K6q7T1O090UjVZGXXfIM4xVRWu5I8NMzBGH2c
e7vL5rUWnt9aBTKNGIPZFWNExcNmrqfZawo5Q3qwslhzyy7yg6UIG8Rz7HDSoMB2
cyJ3Jwloln5kajIep8UlfU2gcoruIKiFcX6lcWOsRWe44XjGHWKrkHh5B7Ji2IhW
onoWqC0hFlv0c3HkaqL2QNnEwEvH2zPkwSX9qsShFC0pOSfRb/WprMjcNI+qLim3
ZEFqppTkmgGwWVEcHOb1PVmP3bIP1GZbgDwqVJrbFsHvaQAYQYufeibeUWJNE1iJ
WeuQKFX5bB/ShyH+x+pCUwa09e6OixpZEBhNrGScchI1mqu3W8uHxWYsU8FnFggA
93+jANeeNodxIfllR3+aCWV65HRXlY9stem1H4+DeqKH4KUaakubFF3AGlp1vFJ3
U8zqZEwwbgxSeYGqNHouPN6LZXDb+uKUnlcl0aufLV99mdDdTacYnb5cgiBF9kRF
GrCrFxTcrvqgp1S9g7v5q/hksPH8iXFar5P7wr1Bz7+IMPSxX3qH8SkOxrKMa6Y9
KzW2ruLL0/fchJ5KuhN3GW3GeqFMKxeaLeDxZO9rmVmDvhAUXTtqlqHJQ8MXOeAc
OxdsLnUDTjp9UQHIEooArprUUqtqVTsUac51VG5PSpSwF5844+x9hUrdIXOVrjqt
Bzv6uMX06nNVIj692UpYyT1SsBhvMGwm+YsWsd9cOSOJwpPoSfGlsPmRmSn/yoIK
4ALLrXiihGZg+3GD5fd0ACig1IdofHDhPW4wp8NYaK3UhiMF56oneLdPvbsr7rWM
hqsBSQtSkoWCZQD9Uc61WWJlDTbqjTaEizcdv75+bxijjjV1bGqGVEfMzUjnY9n7
FbLYKdIhMw2RqtHuOURM348jcQ88h16X0tf8Q5LuS4sBArx+Vik4b0JYM2Fyxnpj
0ADv865gGSS8kObGWhdVpLfw0TGEZTNfdvrwiDKEmuz/Ia/yNsHJwWxEhYQRRVca
vOf0HlC1ZvumZp9Q0OKva2wB2Myln42RmMwHN3lhZgZeLr38SccZtm1W4LwX6/TD
FdZmJELDuQmBkTzPygZAIeqBpqAXaHVd9F06D1AYHZzSRVvB+u644irVipMYY/yZ
cWTPFLyXOQ7HKYXcstev+s/t4Ttrcn0Dyl+wKSEGWM1JjmtmdC1wQM0IBJj3zb00
IQcHNP/MG+p56cw9Us6ZThGjEDhz+T9D99yW0pjzsMh5AirAaI02Z4qB5RRC5hT1
HkDgvvQBj5NI3K/kY8hmJUlPivesEzW2FDTJrS6WT91XUf8abfelG5GIPEMLI01h
fA7JpdFB1vowcCZtxW0WE6Bbg7jfMbA4FqndzHbur6M1dx7niIaG28oHpGa7gIp4
jWvu8gWKs1TrtGd7w8VozCSvl/VPswSjPMPSXvBOmTnUaEPlkWU2u1Zx+PwekZPZ
usRw+dCNXqKASD1AQIdor0aCXg4KNm2VWk/bce3PblhvXm90lCAr7OIPWf60cCbS
gPh9pDJUA8XaZFLHM3mhFiDM41E0JRGbrJR1JZaW8SenON7UOJrmZSOFamO/DfHO
Zu1BE9e/+bTP91F1ktviXMW0p8rb7rTK7zewqv4bplzO+C+bvffMwbK0mc9wQZaG
8ZmVGOefAwc4+ud41GbPSUxYwo7TA/uan+sMpiCjSAhfbP+aCMQN5Ffb/M5ZSOIF
lPx0x63IDxoAiEF1qzCvLflSnpGq6+XMyVXnvI4jKyI9T/4M6PRqw3++TqTvOnp4
JcctADnteQM4dwIUn0HekyztuKN1F/R42YwncSZcmYv+Y+p56Qrq9zVXbJbWvhx2
Qsc1bBpr8S+bQOQzwdCbssNDDtUF1lvtozv4RZK7VqpgJ12NMZpK106M0XN4991b
DMZQ9lLRTYyBX3Wf7UyGNUnabci5mafxTQK2i3llvP0iFJDngoR4rdiYhmytXdB1
TwjoMXCd5CYY1OdiJf0i6rRT1dC/P4jmcAjH7uPymihyVOGTNYnGmIoqHLpHbl8D
tS7AiCCncpo3IYWb0665b4i1rPVMhbRpa4Auigy4k17o8pxekd8AQV0nArJnZ7Fb
WVpckT1CHiGjzxj5UAEoloMD724S2KDa0p9COEPTgSJbnOB51okwvTAJ4mE3+15n
at1XMw+Ug7bWitk8fhlleS3lbM7I711EHUU2IJnzloxpcVflHgJD8bUuoEkC5a6b
F4kb5XhJAf4dbnn/nCyXORRO5LYbOnQ9kU7ReT7en7NYWj8g14UsVqIZOLOGnV+1
cUeYZGigHmYjsZEAUQ8cAXgbp2Gcd1LBkZleshA+mNRTeuRP+HCF+6H33KfHl/cj
eKrJ89afDFzBcoCuL3Dxj+mY42QADh7H9ZwIYsxE+3cJUNBL4iFEmXjwRw6BhkYY
jdaPFDhseaBIKo7cyS0xaETuNWfXgS3EXs0VfY6aK22xmEnPfQ6fBeWLukSSz4Oo
KwRFw/WDiwN1YJNz0/UXYYUiNna/yPkS8eb1UvY3jV4do+96QwVt1LDyvCBYrztZ
0qF6LbgQKdTf33FXXzC+j0ZorPq03NeCclDfKawgh2IB/rZ1f8wtbi3jl2TcCVTb
Il6S3FArV0qgQ37fhCeDDUxxo8iWZ+b3r7+Kga8Ux6KtNaVSZfGQsSL/rHJsKmPL
+ttbCWpBEJq80falAW92CWeekfyTbzQQwWHvN8L0ASCX2dZPNkC3vWnamyteuqcV
Y9u9yxrmC+Sa0Ys6XLCiLV2NyWTPoybJ7y5MKW/pNdEBnYlThFt0bBiai276uhrn
SEUp1gRv3vk5NeNJxzG5KDRu2+bShvBSoe+cQBcCl64a+0m0N6SRidBRAgMZ5SZG
/Yv3UOyhJ5yejIcjQVdGOjIxBibn2lbAUU/QbH4Aph4QAP4287A2pgSO8wPsqehA
UesoPM2aor8tzz8oF4Zz+mL35nggaF/o0t1leBGdLKAeJz60wU5JNfhmDl0RlaeB
GWVtwfKYbcpmqKvli4avOsvrjk67e9Pw+obNBFv7gycdD3M4sCLryzaokvMBTWrM
hovfXG5zlXgglg/zX9Oo2CBeLctlA28Yop5WB4ZIaTL1OsSuUZWT783FPtL457ZX
nUhJre3eFo0Dt6M8LlGsFQmg0aXLivKN9UWeeexw2mSmU+0Po9KLSLKaz765Ywwz
MgHUY0x6jI10s7dDTJmzjxPe7T2sNOEq8eV20TL5duHfCxE+jMDlaYj2bXGShTgz
f8KQ4nckSJwwex4qbjem4YmPuHJgrfJWR+S7lesdh8kBI9qn2R6FExpWWloFd9o9
ZXm8Zftc18LA3WJq+tpy/JWxAtRJxLgV1ZkttA+pmrE+Y1oaW3Z8t0M70FHXykyw
dvUpnKyUvpEe0BjpecnZWYORwIaqSqEjErJ9BxAAr7tQ9PDLqv+q8AaQol0vSf8b
PPjZDgVqGLpl8gIfV6blIN7+y+DhDAw8db6lIR8Q1NiE5AKKZsv8qsRDUKQhZQzk
cHzCp4+ztvC2ZyEqBVg9Hjx5utReucamvAtG+N9ZHEKJYPddPxge99SbrJu4RNN1
ld5B2s3uLiUK7N/9CmY2lnNe4T8sVJhX78+re7YTOa02MZENQMwdfwSYtAx7tvH9
uJJbUdFCFI0HnzCWiMHscOBGmOLfNfLGPtIh/e+Py3XpIDz3lC+gYaN8+JKd5HJ2
fFCHVrZaSjkhGLcZ+WaU3Z3Wrc3sx7ubyL+2u9f5zKe0v8hlMkEWFMd/f84xaJ6U
dliljTYep8pxFt5TeXnYzoC6A+ONva1jc+elu4r+jT7HZrj335SmR8vBopHTZhJg
N3ad9CjKtrGg4hDD6mdD74m7sY95Sab4Aq0K5r0owS4Uu08557qeUan/4pEj+XlL
Ib1OlrTNsksEOlOnmCaU59t1ZA3l8JmymlhJIaKSKZ6naLi+DXrdwmOBhMRCoifh
m1yyqD8tTKKszgYjrLKghLDEHztJ74UWzDMIfG+7BcJ8TacW1D9BNVGGY2Q6Xlp3
KBR4oiclGpcTjA8Y8JVQ/av2Vd7Qw9ZsnJ0zM3qMvoeny2h2B2VdRYYSTnm88jp/
TsMa57LxLBNg90q3LnmTFe6ds/WufxBOxJkB4HuRIwRX16gnU1XoihVtYTgaMmEf
2zDsih2sh2osJQP0ds1U6TfT8gRogUcPMbNjbiCxtZQlC/hQQ8JJVWGKyaJqRpZr
Gqc+/k1kPDmScEWg1I4F1st8ZGhEffAjK7d7Pz8BESdMS+vEMX9TPEyMSkS56oSB
s9mnI+YmieYCt/4BBrvSh7KonPi9lIvt1nigneR4v0iBSGbWmmEeLHoskQWeQE8n
lcZOrpVh+a4wNugkyam0TWL4Oh377mD5nS0+4VX6yQ010Op/K3w8/T1YZ/BtiftT
t2Ov4f3fy2QQDZZ60xBWw8wBFUlnz+9/s0ajaxXTQw4bTeMJ33yF3SW0aaeWf3XK
UOgEyrff/n++9GEk5PNbdIR3bOmsC5EUq2y59CG4CWMj+fw1I2gbb1eavlQYuums
C6tZizzWRfR+OnMQi1ZWY3aOXZ9XvH/8nKO1ObMKztMB+s0DAMKDqcRk9nDMw09h
b5CRqlmxJf8gRLhRKw3NwcAYi2cYW39kUvvC/Ch7KsYgCIyN+DNjqLcjlpCkOzAm
pd0sTAFMLBWz6stijgddmeqjT2c70caeK2n7MDb+R35/e/1tk4fkQ/HQF4iwXPJO
4kALynmksRWmDZmon/E7/bNsgJr5D45sLIDmSX1P/084Y4jdz+u2mY0Fioe0npzX
n9CiwUJWsnK55p8e/Tk4AI+M02GCnTdpLyuqw5/mEy6dtdhVtOaGbzoCIdGAcWar
nkstrNzAEslpD28a+KpcBDtuiINwEcmjkjxR3r59H/TEzV7+m1vbnDGENnMZCg9m
D7v+RoKuGTxF16AF81vxNSgeorCozxenMbMiBhdLGfmcxcB17IKHXSMxSOnL7B7R
qBjGXNZmLg5sD1FXPlyiNjRbzJorDNlGN7FttSUJwG1iVl20SKcgAsF6TnBCxGVW
Xc4zbdLN8DpTJq1z6uyxMpP2oG4ryTNspQCFdxxGyucNadf6ASa0Y8Jd4VxaGal5
jvc3KbiAXd/jgi+5l1zOcEvvnV5H4oH71QXop+lk7vIdiXAWlRZS2bu5S7X2XcPp
iAp2fdPwjX7ktXD1sZNikCGx7mqrR4H+5qVROtIv38RaZXqQzCuoAEJAL2BbCuTp
HZVfaZ+xjxAGJ8PJp9Vi7atbTtUoCVTLfQq7anBNmqS7/ZVvZYOG/Bz+C1HvCvUb
oWdmqXc1k4f3OLH257xcilr1i0DzDbGCYeQX5+4MZoWOlN90KS97mFc/lsRdCRY9
vVdZttCRB7kK71Ymjmt7bsboqznCw8EIMGv1lbyK6WpSzZVGJzEUvDaUMv2sj95o
wTM++SKC4JoxNlzltEt6rLcID94VffXN2eY3SmBoUu+XvMTkegsgTCZ9xY8yQBOo
7UWE/SCsVzFGCJDFPoddfM1iCBpmfB27820ih5VQSMvN0j+1N5N5batTswkkG005
PLpwTqgrP4tFISsGqLTReZ04zuw5ciFY1mm0cjlfmVLitb3+amejfPBkqfuq9/LK
FZr+7jWP2idTqCEnSXHJwnUlFLdXjFhIlPEaLzMJiV9ntp9q37STd99K5AkXaq3r
83deVZS9sTQFSKSWCgMQTTkYRWEdqCzNJ4v2sA69sxJjCRhaAPun53qwPH01R2I4
3sxY5NL2ar/242KO5bQBCPfQTtDtELd3vU2iYq6UklnXq9Ny1VvommSavqMJvO2Z
Olc4ggiRwgQjIAt3gbR1kA2o9vHURVrg53lOu1Qgn//R+3JWniDmjnWn3nelNOGt
3bM8IBtwNGyFzRmdvwy6DiVQqkq9/oBuPDcIGratudv/ksifWbru310JL2lX3pvi
JdSXP7q1OnGas/gwi507kSyvxDlgCXF7xy+HBvWEbH8IgiHK+EhsA0OMF3qSZIvQ
7o8dQ6VLiFfaou8fqroXVllVkXUKXzyRrf0ytaZ4xnpYj6/gFv9iwnoUch6bMIhg
935WV2CuYzt+aqNHY0vCyb/9xIxl8qkXOP5WE1n1ohYerbfSnlPvKdPuJyQJJREu
KAE33Jp/A0+Or0Sicbo+bV1kBg+QbA9ygxSrtUrUTe4hgcLnvNHCtEygN87KdOdx
hL3/S6+OdZUSVF2cdfHI6CpEBbTI5fR1Sjr/avIy7C1SEvj7O0IcqdQlpIgwbQik
LylwDw0mZz3Dru99k20RVJ99CjCfw87709zB7K1mU0cACB6rSzjxkaMDsKYsExRb
bUdD7vqaWyAJ/9IlhtR0kOgEi9dsIpACFJJ6AxYV2UCLEV15z91u31NOf8MjF8Cw
YzSfIsx1oKNfIXiB2etO7rfCQV5yfTYPy+JkhYGzsP0a6NMx+WOARKFFfr2jq7yE
T1HVH8jgoVi3SraFCs4pdGFbmaMESpvhIJOc2n47zhNJQ6S+SzE9R0T/MWqv03rc
8HtI5Dkoe7a7Q9KyGE3V5c0hljaxFnMKVzPzRXdhh2uNBJjH5+gBFhfJjSWW2uu5
SsCPaOs27S7zoElgxQgoEcf/oCGvNCgb4X15HBN+J3nG8uQ7p5XIX3MRyTaBvVTt
MA92601bwLhfqK21mITh4SmyAlTOhlCrxP225CnMO19dWtewYIbfQloufvQZT9me
3LV7prnwB6Y7QjNGrQKG62fXeOT1fTENvjIZXGFs5KM2KR2CdhnMu1/aCaDPiQRS
ZW+HXCwrNEbvt4Rt3wViBrFzNb7pFZkIYV29L6c6CwSUIApQ43vo18KI9NLPwb2f
sULKv2Hgfz+6HLw9PNDTYhg2fHYbPk25CWW7izzTmtQHW6v/Su/K2MN+W7jFoV+u
L0k7JCWUaao1ccZYEMD0/0RlCvpneCAM5ue/452MtjutZKv4U5gPou3gCqAtjjPC
HI3Khd8kntsvL3dLsGHZgPjVmCSYYXmbcASBths/PmjokUp137V2ar6tj+tbwZ+t
CjF5jaDIOo68NSifiEdYwm2ISiYdsI4J+2UQ4+FRsz/DzPJwb/y258sGbbD9Turh
KFNAF9hmCo91ZZJqxpVxeb0e4QiW4ZRbprvk/NkUFFrYeYyYebC/tLDXVdavuOS9
Ljq0Ugl/2UwKnsMj7ApZbRSixM1mUmTDxjkU1MoYNREqmz+eaUEzSwA5Nca3DhKd
Ph9L8SE5+GE9I1z1Bm7UvYlAgbrXhYbvGHS9mVvy9j0XjI4xP0lzw6hqujHnUDzm
ZQpfFrdkbI8iiUUk/Ho2favlG7zkaJ85LlQaPpphv1VmkOwBmGYx1Iukl3t771Xz
SJDKdhDFN7QEba3O4J269y+3icv5y2hlwJJRt0XMwnkIDw04pOdd64usZwA6AjvI
HSDysalAHq7xCWa2hX5vkAICxKlhX5rO8WWabwU2zVyGezs+2kV/DQIf1DCDc0Io
sZwFpQfcI4fyErQ7Vpz+yS56IAp9cC5GbLFTFzuotamlpYtOo+bs6QY7ttw3KxOe
KIo5TzQulywXcHMaDHpUiKJqsc7yrcl+8qB/BecWZVGPfs+T1sdfjscVt6/cuSRY
Q2MaMk9T4rxEtpcU01PIe9pKQ/urAv0ehLzqE4kFGXRoOluPNplNJVq8eYNEgYcX
Uq1ZL4DF7Zweu5YhhXoLaSomCwP63nLTE62Ya0yRU2lzhrJuPQDr9bHfWIsHcQjs
/lWZwwhnEeNHxVxoVvx86HsEOhu4U/zWFG4icm3diuVN5K97N9mDJsjkKi9+mRby
hZscX89F6H9CpHLiI+tdD4lDEUfuhFDFgU0gn5eu6CiSMF7YTNQwRQO1a9bIvt6C
TeCxyWcHeEF8FNJC5tRLMoNqDicix1D8Bj1dXwf9GTEpAchnc2wQMIblDJni4gBw
vAOuj95R4mFEVa7YJY5x6OIPT3AJ8keX6MY0gThdyvCkYB7XM7+GZs3ExmKDUDGd
OBav9RpORc8Xq7eyrmzaNJ4aJnS8qxOMz5O8op3l5o9B1O24RO8sHe006DxoZd2g
gVYd/QEKe5ucN9lJvif/U+vIB9mioSJvUOvbzgZumghC7XrE5L7reOP2fw4pqOA5
UwinGu2ZcBvI08XLJ9E3WPrFlSBGDq3jRLoTOOqAsTpfKp9N2JkVa+zTwnDR9nr5
meE/imTzNFxdluEnrhJ5IMoAKkvwJo5qhFqI+hzY4FHy3FuV+QmGF130WzrMCILf
g9F6qtOJIg+rUx/vOvI3HjZ08iPfFz8BVh/q1Qpgd0hf8TduF3uWGZSslgkvB2bL
NXANewgavWa/ok/1R0/zfkip8D6yFlDabdScCNsfrcoLObjTQcE4cSmzXez5UB4K
7VjsLSlav29Ewy4gWHGW8VXmw+6EFQPHh+yQp991FmR6bhiN8s2E+H5f1h/2uZZv
xDeecvkhdsCPCdlt04zY9HWqPZ0vyt2ZDFc8VEvHbfI3mzuV9XnrD6jGLh7U2r8A
ozh7xW3SpHVQa/4+bwLCiZgJZtarfL1d/4J+yVy+a37Chz77dGCCT42Twtclyom9
JX/c4a6t9epdcLY4v6aCqnOnZ2HleO+qjqD81LrM/2NWDo0Gp91lZOy3w8t/sj1S
j437YY1nGFdygOyhxQLL9jIfs67SfC2N3zN5ODnq1C2CSOlrJEdfg2jbdOsOot60
msU8UbMJ65HYdbWt2T3kzD/gXwO6314RiMiRTbAJxmDMX09T7DoW1Nhgh1P/q9aM
jXISsfTePC5I6LgykhW6dVZCaR0vPblS+q2MHxCLvB2GsZUhICnv6pGanql4gsVd
McsCjnidLMFi6l0C4fdpJqUM1BVQrW4i4hok4xTCzhriVhDmLNbxGDpLM/YDtdHK
PjdNrxLfhZ6TpXOq9uraXJ0TvCZlotw2BCXYcsHRkVYvJwTlnO8TqEwOSDVYqpLY
aPPkYWjnbGonzUzwkYJZrj5AKsA9jdljtrON9+0A9XHJ+QEPPTr68ib3ESbDyEJP
lLQCc1bNKAa5h3xjU+IZxCfam6v4360vTbHrZXp7De9EbL4x9/yoY0DfnkfhxIq5
3xp3lD1qQHFHclSr91riqcIM0QL/O2+QUI+uYTWU8rPnYhVN7ufqx+f+nhr/Wq6f
x3AubDmlHmFyGMngu9bSRekEVQCHNmjKUiFjXqByJ5CubeymykN8oK5WtqXcGRB5
QqrS8vCe5svSnD5OefKLKs6lVFG8DlyGBXC8pY+M9XyJCZMwArlQ1dgiFYs9e+MF
E4amBC7LjqrgoeOCV3aRdwPz2qi0FOv3xi4xYTs3/5WLLHxkICC4jDM18eyYz0+A
HEOgAzC0ZhwiALLe0mNJgB3+4/FjH8B9X0EfHRa71+B2T+SZUCPORoce559W1VmT
4oVzPH0XD4/SHjoOT7rqEv2aRZITqNnh0vv1cC+baGCCTSvhBI26NDfyiH+wba7V
IGCApVVaiPneAjD31MmRwvDy/AO+Ovtd0nE1dOMF+R/NzM3D1BiaWlEqCa6cCpg/
km7rS1FKFEyZX9x/5BECyUb1sCcHxyqpXK50EWbmU17toQQktchMQhbD/XFwZ+zt
ySnmoUu+FvgqCA2y64gygMFrJgEZGstSvHchguo4bQNG8PBIOVtkqWOkLlVf3QuU
PY8g74Ds+dPjaLMRTF22Zl0nVuHxf8vTHmOpGCNgfGXSAW3gbx+7mk6tfdMZB1Gq
ePkNaJH+6uwnMBFr52PwDnGSNlm9+LI/hjNxppFPDrkdN7o8i35pX55Pv70fwED8
jNosAfp2gbsX1xQ9OLQgu4xqSmKnQSilGRWS05ea51CUWT6gEZFvQsOYiB4MuwdE
dQq6InOr7Fx4vUvR7nQXw2iovqYOCd6tzCHsn3MrKv+i36DrG5/eOpR2/EQegTNT
zNPAgsvwp1Yrb5eLoKAlPkYZXZVNY4eAphvkmrN1+RHyc6cKJs1so4MWsAelpmu6
lV273OppSgpyK07PErGlwww634QlJgDvz7e7jp+1JVUCDG+zv57u9nDUs4Wpe6Zr
cMv8BU0JCUs5NxEfQoE2xi4CaiVMw8YfXg4UHRTb03B5QhzePObfzzHl7izcYTXp
i2PcPisJlBPK1RcGtNRNCyfSLTI/8GcmVNIZO7YR1GqvBzOnqddw1w8ZRMF2KkI2
QY33bmXQAqnh+ZbSYL5jyZwDP9vy0cjsYC69nhpmhI1xFGytXee/UkRsllqQpdo9
PrSZs5jnsYCBSDvFiERIt37wpost656B3qqIL9g5yukfiij/jXmAk64HpuH1rpx9
wj5MMZGlPZfwU03xsPN6gPZ2wns8TH469Hmgo7BRHlBXf2KU6itb1Hc0PglOgOhG
WrQI1J+k8TFRl4nZmHyXSQpVQaps1LhzuK1cVEGuyoAzRFWIOiLoTjmXIHz2hb0F
fl9oheSCkROMN+AqzxgQjCuXUZQ5WEDm9brk7Kt+Fu36k7WV2sQ6gzuMKOrZCaXz
BtZpLeyOSrJtX1pVgad35iZZzDM8nNHdO+05+MFFYfrUQ/e/iw+0OdJ7nLCpT5ff
ez+fSFeuoWJzEkbrsluRysodmPWeXQWTaZUJx5VH5BtSdjBnFUc97eME72glSLR2
ZlgbbJ2qodJFvBtLEk3WmRREqMEHCCr0fTYibNAk1s36xQR+2pQXifABK0o54X7/
WDLQFjCUKLxjEPJWdJsrMB6BvF6YadCzbQBdxoBBQNPMH8MdlMasR3XtPCSmOaQA
Vmk0leUxZEiJh7UNj2fDI5vvo7RKIOWPPEri74aOd+jqN/4/S3EFLmI7nNV2CMKA
dAupkJZ/RfiiRUrEmTqakY4msIf5A5UV3zkQY89ijwElQTh+8ir2V6134xhV4taB
2dhPqBo9g9QdHj+1MltGarIeg5GXb1BJ83v3wVw9dhCDsYZq2JdTDdxWv/CQfR2N
V7oA6E4iKYv95UJtWZ6YjhfNTJJiENgsn1r3Arkm+RyngFfbnmEnEWruKN8k2k/8
ynQpW7G0V21Ur1RWlyKCEXJoH9kzdWUoBjZ8EpK1Jte8clNTToPSMKa9BrcL8gBJ
QLlYkiqaRX6pEwTVeKIQk0zL/qykVLQ2HANMerPpVE6OW+gSzoi0QNkSeiOmH9XN
pMiakYr/xcwJp2EYlWbjs76c1eLKjRNUsgk1VBcwccR8SpqUXo3SRfjuRWuXaCjr
ARl5hJBkAkC0Lz4UMJvnVwu4mCTNqhbzDFgf7KRLjnYexcq77nePeR+9wNLPfrcu
VBaL7QA/V+Cw/KPmucVeLOSqSUdReVKf9Cpp+ID07xrWmcQC+coCFi/mDecwPyFq
m1DwjJhPtt8lokVh6dI9/Y/ME37b9lZLLwnswSMYm/fREqLZH/fIyixq7tI9IFdh
f0zQo/aeo/b2njyDnRmygRo0kJ+H9LRTThnZ7rGwOfz30DmBezDTuJBhN5AhixJ/
w5J1eDgiyAdEwpOam3WdtVTIPnUvGmyyBDaPDZ3DXY3xJrn+Brn5bqSkE26Y2Rcb
kQ3NvQnCABiUW284Bo77Uzr97VxLci5hzCLi8BvoxFXjLxv7Dr3rNBnm8UOIs333
ATLp8ys2epZ82W00zQLU4MDnvbvEfjKHZK81jALtsl0BePY01+9dJelOOoDitagJ
g9HKGqNNQZv4WD+MveJTml0yXldHy67xsPyyqTc2dErR8cWJoOPOYO/tHekSJkoR
4Oo2OAQW52hooSGqlCeLKJONoAgu3QorzcG/2117gwD4pnarmhwJ3/kuSf4iWdtP
eWQiKQ66Ww4tkmIeUt1bzJ05vMHrjV2G5o1h3VrrPltSu7ZQC3Jkd0C3vBcFIgeT
3CUKG1IrTQMC3NtqB5aINvT66ENlqhzsGRw+5VtcsmxQpb8q0BjDdz3vTzDwpP2F
16h3DtwnMPKFrAn4E4MgaiI4pUtGcQKAd1gam68sJsMzd2nyTCvKNxxwjftmXJ0l
0+2o9zWY9oQjWF4/A+s1xtjk/TZQnA5VDdp+xA2If3Hc2oM0WHej7b8/V15/SM+h
bgvL1VpIJ0GHsWw+TUZaApfpnB4Do3T4kjUB88d7BFO+DKOyrHBL85XaH1Z4hkfN
QwSsRcWlMC3tJUnmGLoMTEtHQmwYr//C5C4Q3IBbh86VVHOuasO02IRbSZ8UDgJM
uV1y1U4lCRDKI8l5V/hSZqJ7/Ia8zzYN872Trr5l/F+Rz/R865iQ5mpRFMkSFPxm
lR+Au2OKQJ3yZUnlkT00CUZZkWyzmnV8zkFEbkqGhdyTFteb5zsSNhdq0EreApU5
Jav81mdvya6Ahz9HnM3B/Oy37JmPcjMT7G0hN8w4AYwkYG3ZzTH229RpmdzP4y/V
tpD/RexuxYK3ZVw0aDrelDyFdtcFv1hvF5k7UfSII7Op/x4UQLuh4W84Y+XGugGj
V7BXml3gZFuLbC5tZ2F3sl1l5wBktuIRmWnGkK/NYQgswxgpQnDlFbzrC+ESCs9y
NOjg0duHVYueZNxSAqlOK9ZEGQ3TLRT2KjNg76mOBlX7h3UvNrKpJuud1eVdm1VL
a+yvvAOI2MRLuEDYfI+m6bm6RTrj2f4NOrzxUWtVHmb0xx+4m30m6CJu/OQsnk7k
PSAuSJBc9ZfpmMGq+JFFMGFoETHRNfZ7FM/1YlSAkyavSjqD034A7I1eE7bBd6ba
mAqhF3LDG3ugFEYh/NasQ+HzNhEGAN4ryMdhWXLP+UUIRIlYmcxiNoVmmWGJy4BF
szIh1UNOymkJQOwzWlu07xlmBSQFrMpnGR/cMZ3xL/doxuf+f927SkMUdigYVhO7
6N9hQZzBlXu87Oj0KJdqMQks14Sa85dBVHjOd9tfSjtfIvAhaFfZrqVZHb347GCP
S6rRXvLXPkXoUXcrQjwYx+wUPSE5MEgI4mOxQ/tBxr82KKnA1HjHyQMwBY1ZFPLy
IcuIbTMoB3sGOFuXlMlO+apAsSa/fjL2CXMGgaatmdvTcNwc6zmr3ZFdVE2rwHXs
3DhDJC123qiVekkbSMmm3mJnbmdQPKAybCXnvWdiVSRnIo/BHva+GozGxVJqlC4s
RuES5risWFC94/LywfpZr261bnRawhNsa17kBHOqqL5bzzxvzMyFKn+3RGmozV1f
TGwTsZ7uUYeYI+35QU3ECH1Dpoa87J7Wh6e3KqQdx2vgUEByb1MgVdKhQyiYdlS1
eKBq3KaxnhydWTRSyh59x2OlqdsSFYYPE3FVLrFR1sRK6fld35zrFbXaSTx6zIzS
IBsLTbdN+rxOVZp+K9F2wc7kKAUSc/TJxCW9fVReOSuIYQ3nraPPSxVTx/RQ/mqy
AALsYs+nQjskJGeIIqXvWEIwuX0dcQ3vnFHVw9f3cUK1794k9wA+NfmAmmthnIKh
shXG9Hmqut9+CPdV5a8iABN+kIi1lv3ajIAeKHxuiYAcN8zF8mLz4Jjue/y78j2H
LlVW3ZlgzlSYZsyu6U2CH2rax4HAaXOUw+YE+RcIqIrLRMytnG/zOK9bTmdv75Ue
9W19jYOl9yaUznpbhMWaVNGDGVaFxvzNqWWXJeFc21iZv+BSqIBIZ529ueM1ZuCW
oMU4SiOMvrYME11vuUPReVPxZRN2kZd/yeomlqnaZQ9LE6IxOQt6aLa1ezPbdpwJ
RTQlx+cKjym/AlrGUx8puf7GN4szGXXkTplJkbtdn6MEPqrGOPPW3hY2Eqn6s7x9
ScyOUMUS7TPBq05S24rmAo5Uu3TOWc4u5YCoA5Wytdo3L05u7B40O2UnkDVorcZm
wRg7M4nA/R67lfVKX0h0mykjMrLT93bXsTHQwZYicG+yQ1tE6WGANUDKM5PU3bdK
A4u+CH0jB43m6apbaedtgchGp0k3S/9Cn9ObmtoR5gwmYAl5mb5Iy/ir3W8YQ5JE
PtjWoujM0RHKAL+CXddi5k+nBlbBRVpQ2E125yovTmqBWqBQstNtLXmPwg2junGN
tlCtj2Xt6Pe8xgCfodvGIqA9sk3U3XSIEMGW7QoAwEjXFPrywpeyTYp+P1Jv+uix
wkAObsMVULbkPGx77bmm9mZcFvQyI70pCQ3RKnOY0XKirXFOY1wUSA5jWhHBmzTm
SROWRyebcTJyD2+85lqaaGnBpPNFsnIpm4KuZLB1sfJ08rZekerFuMaSM0YgPPgr
mhqi7WUD7LkVuvZV4abLXMGvusQrqPhhcp/ake0YRswXnLujZx6wtLgVqn+uUndy
c4iw/fg0mgGxOmm2Nbx7a0M47HMyoIAP7DWvNrCDzYE/BhEr/k7lJ493e2pvLnP2
PJ0CS2TmvK4UEEz6299gh34DY3hwcAsM1m/u9VhHibpUU9OT25qotPoImXQ6q0rH
frvaOdl+QPDsavpLzKzYnutMFtVHe+m61oRP+1ChS6i2qZuIv6APHjfx7PAqOGOj
LEBJ15kGx4BlipP/t6QwfEn+B98oOBe2AinhzF4E+H09KxdbmtKHmBucRqkPg6J6
2Zo3EQ/sfl6I4vwSTIW/cdUT6KUKvemrCmqCXhsAEjRjPsZCuTMy5604xSYpWaHo
TqZmBbydYwJce0uCUBkDcKcgSYj7oCBuV8HSjF5s927+7cJiBR4p30RFM8YFeNj0
9VAxgm0v6uB1SNnFAoLTjYYmGYFxJIpUaGvLnwiC6koDbSpag1g8/8qGcxtU8iVW
Z9WctXl9mixmkO+uOLfuqIzOXErOupgG+wJUaDCds4qsOyFEtAN8upYqZxjJU9q2
P1IKFvThumgI38g2Eb1hvHhw6ZrgnZbmmgcG7EeecW21bORYNGzhCyLkO7yyIDXz
MXLzAPT9513YVnuITPP5F/Y5ITQWzlYLcJbFS3cdFV6GAxQ7qdYeKcOqAtN2vLFX
ANYGmCxfsJ3lB32OcFjB35fCzybkYYyms1FB/IQT1RIxb/Hvom4SEWebPdsmwX6U
eD294C1i6bygseQ8GWRRmWQKbmfCDWmhcPy59IKkPWanNUSRuXuOU83GFSdRIzH4
q0X7gJi1rE9mjWd++mwsMc6+WjDHmkE+QPxswLRGtOdPIS/bkcbV+7fJVr3gyT44
P/i35GIKR3cayQIGh6EdRHUCYIrC0G9iKi+00vX8jPG4e0cHthJRXE+sOicQP6Z5
HfLOIiHOd1IzE3HcWuf0roQLpnOZBu4dy6zVuMzcNzrwtP50Bp4x/ZR0aR0wQtUD
cYKoaEVDYl2svWzbCdcVO1WKVjMUceM6hqYfMTd15Lh1igZAdtpxjVUE+5opPnzL
kQUEIBqRVGHbJO0fbP0oUDGnAkshxgWgGYHqIz0yfvn9CUz78h7FIuGiOqvjb/sg
bl8J1XeWlsg0nN8Gt4PsDD+3Nufog/5LRcjZNiVcYzbrX5EXKyuZgHZ73fjZ7rYt
waKwlOQAabb7uRBJgLpXu1OHxEBANOq96Yyel97ujamD/TC9XpA9D4qv37az9zYd
MshmfJxN4pjM8nD26bbOWz8e0tIf0tQyn//mNe6aORkHPX+9EFBYka6L0IoLsJKG
qxpXW2MiGMj16ENeCd/vzlSWIThP3LHNcssX9eCc2ko6N3CQgJhvhSZNprUwHsBO
rp0IeE4BrhOjZWKTfHXShAoBZ+xJNmDMzIzGwEM873nbBLAghnpfvbh7yWFkzIMM
boUBoPLXjMhO+tvT458iAfCz5NAKJdrQNB8DptShDKxC1q9xru/o4qDs3KmTXd8a
lALt5sCNyV9+yYjJDleN+Mq8OnKhb0gUSoLBGfRhmHYR8cTVRoe4EX5qUWgUkpkB
R1Z63i/Gw/jIc9N2Bm1QTbzQkEJ7Gv4RxWeNT5Z5y8NM99LQ6lmBSVkctpss8kVI
OJm/R5VbsRXwHonPzMaL7pOpqAjITXmidI8HivtwIK/bdlsDBxojnjtXizNEjbxB
1WUolQaZf1DN19IW614ArJvTH1u1q74rlN7jmy24oRa2g1jIFJTp1w0QPxj7lPCM
HtJjcwh0hSy2DlHbfrGFOg9wacODi0thianiJ5/ACwwVs8r0l7CWgIGzUmvxad1u
A6sVki3YkZ+8zGZ6sMU1wfUjq851aJioUMeJG6Rw+BnkiyV2zzgRZ2va5Ytwav0G
lDNtrxP8a8hxm3l+9Jomt8Kbgg8y3E/Vy0+ExEdULGB2wM+/+vy6xz6hxfhe6rbJ
cVbnqV3HfT2P9kQOHGOV/i9YyzhoIiYU/eyjI+MvY/G6ZpVsjgkklJjXdWh+nK8B
YSH5otHYIE7b2cLSLAITgJoMCqzljW1Y2tL1Akj7hNpS/zC5Rx6JQxKEHxmQHXIq
Accs9mWFZhyDI7SAPTifbgmxZ5JCHaq54XHWh7N0XWCJKGorCsCN/0hXpAUrMjLg
LT0ETiNlXzERjcx8ZEo67MoF461h/FNhiVqzbrTJpCoEvHrSJNP0+Oz3+AoiBHEY
YPfroTJkr+26lEBjyCuReaRmDIsnzCK4fvlUZYWIyV/bGOsuGt+rEPG0K8yyDQpn
oBkvj50WvKJ/aFBUw2r3ZvgfgahFJC517USccD/AHeUoHvmNwiQ0vciVxbKhfpKW
gP1OGf2lh7m+1qhQ5SiybE+YOzH8AFOeeBt7gj515EiNvKSY5QQLnB5phKQRXiOq
Ht+ypFq5ZhrA1YKoQF8xVM99qJbw9wQzoqbLN/LfbiFDJd5V1/0WKMzTF02YctDs
j2xt2XWbbs7PQq11iwAQq8qiTtUC2voO4vLJ5LK4uMtPxDl7ow5Dtw1yrmklKytQ
HNtXw3hpxqa67GB/28LwzJd5zWK+NhpSIhhA+HuKb9wdVVRIfcnF0Kd4h+YmB0fg
pye2KLi7mKTBbaEDEzEwLHruZWHDmNBpLT58STw0LSy7A8HADc/7w/yuS3Y3NPXY
rRZeEpNyhvO7pSK1AZ8SXIiMUlU6mmiOszJJGkl93bHdlFZ630/Ejo1lDq3XOPs1
6bXtGPTwEXlG8vQaxeHDUU/cDwR1p1STx5HFshXae4DTXezvUU53Pklx9PVwgbVc
JwznNb/kQFNbLvvR6tP2weGxtY6CTU8mcWnKMkFqg7IZoLFfYLL4B/N7nAdENkv+
TCBVN/AMRXjzXSoz/OYzncl4qRMOKVuVDvVgQJRzMc8V+V7tKMkKRArgMYgEUm2G
ZSxHWu6c8ZzRiVrk3qC5ItQP1zXFKP+1JxFfWoA3OvOD3Wnl6Fe4IWJJ37m4qRYI
l98UtSkO8Djr5ONbBcg2b4QoT/b9iRqNlSmyeNASZ2VzRWAmfXXBxYq6+dMO9Fmb
vFJzwDnE9+F5t+HEu9tTPsLnK3GgAfRmZlMDwMo0DFSqtLot5t4GeNq2dmipZ6E7
4Al6BM9AnmELZhz9IGYP5voSjxH8HAw3vvRXJLf+qq8iL+6rk9+hBlvGh2VXbVfW
pd6ZSbZXTNpz3aSuM19stUa1uFtRNDj/ARw0CIQkssf1D15v1LMUpPbyls2e41UZ
P+9oseYFbCthd8qnf5OjNxv9UpBI1k2AUD9JAFbp1rilD93C42MJEONtOXkbwflX
2PWn8qmnSOJASz13cKuD9PAmRfz0etipj+3YOw9vTN5BVppMEXuFZdMW7FFw+qPV
H0GvDWTJCXRs0ar1eqeUpEJGVyvDwfImHwBSI4lvmecyw6Gn+nGgGKPAXIQZlDzw
JGxqZnzw+oE6W6On2//XuC0zpdWK/MuoT+HGvbxsZZ+Q/WlYjQWPFUV/TKQKjaev
yowopCGFL1bmCDSVcpxxdzyT/f9tzXFb+jyfifqbcFcfys4FSz/Arlh0etMMi1fv
n+z8jV4bn7BO1d4od5s+EuNC3afdz8LoZNhD6rlJszhOjnsYBV8CAeSCJ63+fgI+
a9qFFrr7q8ntxJrTPgCQ8aS6/Rksd+mQ4UhIom4hbOUR9lImsjGq1B3wdzSFjbdc
EtIoN++GXO/yxTTPNsm5C0le2uKFzA6RSbQuhxnudeD0Ci/cn3QrXqd8+f2S/STl
hXOAOSUozLm7RdXGnm0Mww66C37QbvbAfVC7K6oVUUdz0/dZo26b3HfcPre7JWH9
4r8wdTcI6HdmrtHC0pdoMULSX44lIpIHytPwC5Rp0R5OnjArhUx72tx0TOJu8Pyv
BhuTVIS/VTAe5Gml6cclpU9RvGCtzKV1sSOXyMiaVe/MdRt1ygl0srx4oaM2JCbP
1ZdYy++ANDFb9O5XUY4sDhjFKYmCG34dDbFD1eYAPWjGx6430N/gUpMWecPPQ2eT
HpsrOegS/pHoHwK4d6MjhzUUpLpzj23TUVQ18xj1IJog+6FPKfE71Q+5AqYx86jJ
RwDIrZy6cWaQ4rbOx68PpAM4fUPaPFTSQWlUUb4AB08lozSp1enif1tX7GflEYCt
U+q2l1lSTG8PYfoSh6PEDqGs7pDscjMy8MlJz1qO8zeKDOG4IA19+m6xKJ0uwyD3
IX5zQKxoJQ/nBfm0CNMT2aJiG0vdnNzC7aLd8kRp55GmCcSlpF2HsAJXm2DrtMeb
kLMsJpphl37rVVWgQVTYAYQEmYB901IERC2o9g9coUqjxhsCrB7GX55FE8P0awTM
9RJzEhngWD5uHShIUaQLvB9SXSiHnuMOBVDeIyfNNuxiIGtThrU9j9ASEkyaXdQ3
jlUGRkDYTlgWCBIOiXvn2vrDbDJysolhxF8VAqp8pi6C5ite7wy5LBJEhwfL7NQn
Mxa4trsBWUbPFyc+Z80wXqEdYK/ji7ms7wuBPNX/NkzrM2E/LtLNSBd9ZThOwSOZ
xCX0ryw8trsjHSTYcmbeMPo355TLyPTIxxepROqGYCVcVD0klqZMCbRihOuKHSU7
XaSbfHmWJjpJ8hWQ1TE3Pr7d1fGWYPb+lAqO7FCvInq6Y8AXlNZL85uaTXUbJsTC
/F1J1/vB84b7SohN+h6hDOizExZkrSyIjfs2l6FsICyaKzTAO9NLxskqXZvRGL4L
9u5GuoigLvmX9JOqQNFj5bSsfyp+BKai7l+0sPJfaCNkDZgXf0mD24nJ9/St3/m0
EtWIDeiph/iPkeca74rXacZFQqceijElEVNmmfoLZZGX+1BOeGOQXxOIerMdrcRU
01mKEHNyuxbxM9Kx44vYDxC7yfS8qOJHmTuMSn7zsG5GKX7wBBGddxFNWP6wWZj6
zRVFAm/icEpCrBtAIqbDWZ+urGXh4v/XRttjFQdXywNkRMWtHXVIt6r0RBGydRUl
1VsNH+hqvr1kVC8dE3ydqwQ3ZRoqMs2mq/IC6ci6vYvJFs9Hi/1kDMkQcPN3bmQp
48t/KKwgwtrcjbsgU0aDu3O0Gv1PWhjOJjJEToE1G28T/j2oB5YlzNcucpnKQLUr
1ryP+4eOQ7WUy0plDCLgKOG4zHv5rjUeiYP/OqydmQsQPlSGxm1cHuSrrXetVsXS
7E2EI4E9OiqlgDGI5kcS4HXB/dsqWoIKRD87GbVMgpiRfOWeFq4Uh/DBqnP959jw
rGlx8aKHZY9X/dvVNymL9fUi474oxoLRTGo4+9fGYDaO7a3tk1ZecKyThsCj6BaD
RF9Y5WyUXGHGZH1mjbnnrXrtY/eH7j65XEqZBUm3/kHi9m2O7E2jB/ShX/JoXSlz
OUi/Qoztyf9R3VdBYb/aE8lh9hF+Mh6DuuL/7XRxYhawb+NNShy//RsG80ZtljJq
0Nh5ICRrz1+4+9DmQPQvbMjzl9R32ZbVwiW2KzWX80JYqrKGPMYwWxRx6nekm4oe
Vw0uCaAqwSaAxJ7ch55Y4Mk6d1AOWeIUFejYajXD+hie7EmG2pR9305SP3f6c8kN
ySdFCA5mjfXs6RQEYocLtiXzKZ4J2IhLj8VYOit0dO2qlHdUgaX54CFCytAT8hQR
ag0oNJl7h9+vZ6uG64LWyZMHcPOqhgzBIv9HS5TR0yu+AglqhrdSb3SUIlpVe2Ws
JSl6HLG4EntWbtfSe+9H6aVwMGuPkHZo5amSwRgjkq1O7qZ0JomGM15KcmZ1q61I
VSJ3OwMa3H1UWmqP7n0U/qVdk3R455AMJbuH9MIwIqPf8Vqeg610TodQ/mCdVJ6h
tLgyBS0bHzwmcaBfdfX2AzLqJKij91CGb1zocGTQYVeueJjnvYRRnH9LvdQvNMRR
Gb2aGGyuH4P4LVZbVN2XP/2pfweJQ2k9+lJZGNIhFhHohRBEsjzcBSP/fyR/zG2x
KqMoamk4hJv+wyp++t8cUi2QjRLg80K5eeRgdm3d13UAbkGRXV6kxMvMkCQFnm9+
aMOkRIraRI2rshFL62wNWOwP8c8GbjYLrzrDazkKcFUkgDspk8j0ufX6yJPZS9/g
rdXDHhkfdR0AGVXL+xeei0B2rUX6pCKQZ5Tde0ptusH6xqk3gdg8GJ1y/KxPZ4F/
9hG+vwcyhSbf2Igejguau0n/TDsirc40ZNUlwz089ntMymcPCxD8Z5uH0y/z319a
Y8nm46gcSfIFvbdY7P+Lc3mUeXjPlshqonDQVT+v4p3TlbiDgVPhhRqLI1WAFMZA
Omsh62P+uT7xgAcd36dAS/wNFGq8tyMe3HV8PqjLhofEqRBriy2OD/AWiMaYFDiU
PYgejl6CEGcxPrnK4KSmATKmKLf1pF2y7IZXaIny8cKtVY7h9Oxmp4syp2lM/lDh
w+YFzSmJSBugPP+jvh3onj78LogJUT5C+EDuMiJQ3aEkOB3Uxc9c7XT7cshtX2OO
px3DXhRV5v5iTEw/9lnMe/2L5Ufb8HMAslhFE57JDuxY60v9mLJV07RCdKOYt2jj
JKvshS1hIBfaMO5vz2z/2OSvSjFPZRrSlPFlmM0mQW2eDTr5RjuBkIGfUlWxGVvs
c1axLB/3wjlhi0XurClb+RCvy6tU9mYKkxE/Su0613kCmrQ4ZAUT8uVO0FhQ2kNf
3oGeVgPp2CdaX80NEVXegcouWtRA3atWFaePh2cdWwrgZWZMRvoq4urnZwDNQ3Qs
H2AxgRf9UCBXQrb/aT9rvYWewiHVqq7UCl4eR8Opw8bUXVaUf8vq27pX7pUIEu2Q
WoLbKgFEeopHeugHcjmlWA+pQofayJ7qL93DhE5FVw+yeD/yLIOAHSaVoBC/z7CA
k6j+deoQCSb2F6UGb5oaC0dgFibMXPzNd0Re8xG7yMB/U5yytbEZ1qcCGkOgw8/b
VC1rLOZ6PQHcDHAjt0hyiyOrt73ps7ehPR38lQTfslTbRxuIEYIeKmlYJLY+3lhS
qpho2RDTqva/IxMP5jXcgskZuVpBdH+HRe+Uo6pjah0fwauAsi9MjE0k1eyIS3Mh
lLTHLbaInu1GdM6uPHxMoIpKUNxmNUD0B+P84cK7rVR0ltDG38DIT/dCsUZXcmQr
GDhHg62JzupRufg1D6VfTdvbfUhcmk3BD3IM8DoaYPCxCob3Up5Ai+FKM9GPJqaQ
PWZvmKgXOSJi5RgwreCW0Mu8A52X1Rfkfq7+mIMtdM+Z0xKBR+iwvSxAkoXIOFEP
qGDgbO/QtaVehJIKsHfRMeCCYIq9e5aW6bcFgLgkxvUnzYjj4/ziv+mBRQ5FvY/A
uhnxJOAtdIo6kW6EnWnDzYxQtxJXSswvRYdrDp6FgnM1DGCuVAdPycbK0ZvlWrg4
I5fuBPk44eyB+vednr7OiGc6y1MCfoxOUYfnKhASeVGelO6b/3EcJjt6sBznPFZz
Syf5rXxhpsveiYgltVS3K/KtFBBhNAcac7YF1KJCYeZikDJqLQhgvbgU1NeRG9FV
cjzj84u8HqMP1xXr7ZDyGfXJq/JH8gLveWAyI+aqndSrFKMe4zI4HoDfNk1SbCvk
FGsZRjjefytLQq1bVwyQMwkoaz67WrtyNX7RDTiPh0U+layX6k98gGBbZkgSh6pP
Ddw1AA3sBEvi4wwvMMgu1BJe9VcLkJqN5moavCHa1cOSiUbBUDC0xDcp9agRYGlu
e9yHuwkkuecj29Q5mGKh5dwv/byXPmq17tUsFj+5dBhBiUb13Z8hGRPFjgGLckE2
gB8MiB4GcWEqRM+PpaJ79YyHgybiiqpJpZcDM5B0X80Be1Ws2upUzrubfVVKVodj
INn5B3ngYZBcRGARksQZpKRl8scHYaU9+8iIR3Rw9LY35Oa7e0O8LbYYOWWi2K1G
rZD98KLjVmgkIZyAIRp8rSKRG4Xe82bnX0aMbMNNxRrctyg+FsH51bmzazqBDllJ
zzDMQhun0CkD+99wXj3W9Mg0GvGEE2tIUm1cB9cooiYyIZusRh30uUvwyy2RXHhB
P+2gJYItH1D/De5SO3NoJbWg5PXZhGDnkGRAmzdU9EUqq1+L1K4Vj1pN1/tplwWV
pHZh5bg95lodsfv+3vLpvapcMUABoS5gylpQxdFoVD13dJ9XYdiFpH7CKp6K4LoJ
JKx0JaP2jHlcy3B/yrj2WtGdC5nIXQmWISFtcQS+5qzULoIoBp+qDGKmvIijlari
GRakEkI0gEONdCD+wFWyx+iR//iefoF/zUNXtTCwSernY/Io+fH2O5MVx9PUpHyA
wRaKPr8S+9upJPywVHRRUPh7W4ILLe+lOx27Z+glkfyY8HtlolbIZOmsiziupIA7
GT4XYjkdrbvvA0zV0yffkIsSk45aIceT2vMyGgQp58MueLSHTprsuL6USQbvRu1g
77v/N8BMnsers5S0elbiE6k8k0bUbRhlzap3LPiyuyvVQFdQ08HQM118ftq5kcEc
IPCJPyiwVrCfNvlqvyENyEEKJZ6PzKbE/ckYHKR4EzYACogyVdboLULQPNQfGEeM
Fky86K7G/0Hl4Snl+yvsBdhRFInAGMo9FFj5P0n2XKrBjg1QXEa773qEvsKkr99F
/lqth0f9Yr5uJsppcX+qeS7PkWm4vsc40RLqqMjDRuqNqNDjPD0fmVOlnia0qQvT
uj+/k7nVlFCEdAqgQJj+ZtF+UTonM/grQPrbymjGIqySH8yoJBNDwEFJPhubkbdl
C1qUWuDAivypxiOtpW16MtD449kqWL9NBhH+oFsNaxAo3f1YIcCVC/nvLg9K6fcD
OLulF/ZQgIlpBNEts0AJFoNRyK+7gJP3+oODNOAIX26uRecD1mrOyMJ34QD1h+it
YwPEfP4YlUk4PaEQRtE4dn4IK+2YnbhErfU18ueccWkchxIxtgx56r83jI7prxxF
yHhU2UywW6X++cJcN2X6aTFOA1Wcn37L3uimv3/YHSjZRifqeA/7Gdvm2/gjOtRr
5Vq5GVjHasHIK484HIWSiCqH68S2ymYJY+15PkSGp32A6nEGd6ADfxYS4AteSrPt
Eb5M6VvMNAZaZUiRHCc9+ZkkLP33zUV3yMPCGg4w3UhjeXA3A7FkFPCc9h6KD+hh
KIh1/dXYLj+JcESBXtPAXaFca00m2G3XQbW6z+4ANOmfyqYNCPgw1Qs6OQXK4US3
x04aepzDQyIZJscMCnMbgt9Vj2QIbPhLWooyeDP0DyUOTEzQBBeY7fl5VaxF0S1T
sWel2AtkBWD4San3FfXhHyYVOYwXLmjL5+ENuxb+//Bnd45gYFkrg4iDmNv3UTF8
Nls9ZnkZczX/ppBhdKXn2XxTNPMzpUiqbB8szEDAyh7QtkCwGqm1cZqCZa/9HH4S
vLxZgl9HnjZ/wSnav6GqUOALuBdFcSxfoV3TLrAxTAZRTMN1HA/+xo0oyHXn64vH
tdSvIGNxbX2EKDURbeb9uOKDlrbqLXjWSUU5BWVuuqfu1lcSI0X7qCdSiMTm3dJX
WdDdIUB6LgKyvqhP8f7c4KpCOeyzPLW0lnasW9DLY75nykyzxHlT6jofVOyGC/EJ
1Jut6efO3MnxyzLMvoVQkahRXrar7zFeGH6vdslSpfIA//r+bVXE/4TRZUbRDpIp
ZY4Uokjbfk+UWucel2LAmKO8Kv5+AtbgTDBMShLESLlQt0P8P2klhDRoiHugWztU
XttgQRCGGH7h6a6Sf7+ktHfWrkP94GTZW//2VNB0QDTCcTu/AWktaCiWaBNs77Nu
mGmyC4VZNWUiR24m66TC7njkHZ17vYnUWCEoRvPWkmHckyZDsjJ+r1RUIbElzXXs
fD05x/x8wakbyNZvokK2HRo0Kt1+tWvIbHajmzqOK/cryqQIzku9IvCzRSj0PoER
VU57O5BnV+Sodv+0UvwMm3duirgyrdWri49f4zxuYd/wal6UiT+BTx52bTNSS5J6
/naxZ1oFI6G85+2/QcnGat7PZFZNudDPGudY9XAmuvZsALBKWUD3PAcuTSqFEAdQ
C/LvC4otS9NT2Xvsf8BIWAPzctm/UXOT4Hr/MN2/8zo+5ID83YI9kjgig0kXBwM3
ChTm2z5o1GMS4Ddqnyq/LdoF35n6jNh6FIx91L9ClZEsr7UcF3SdwZRsLw+dC/iN
n074YCZekbkyoUGTkstf2wE4GiNlWjObZ+FSCl7e0rtu++4j3rlywFsyqooCxzII
pEFO2w+FNyh3aDDKNLt/LgZsHljgtN7BfVRnz8e6p5aj3Dz5iynvR+YB/DL2/wz+
ecOQMAnrqtnA1KSA8hPsFqsfZ8WyT8GmgeUHtbIIiObHv+rAhDcGfCkNVGoBtE0G
FT14GYG889F/QqQPHt2yp9LjiyK45USsBIXt+Xjvl2zFQzpw7qKzrciQSb1b1D0O
bB7mq10nsjZd55si319jphNVCwq4kW0s0PmJWMHqNZcaSFJa7qJ6/h7+GCUe/zFg
kyRlt5FN9T907Fvc8XEfy8dq0QXJ9rz4mo4M87a+xTHA8Yz9HTMLxjYyNL4ndpS9
L6x5NaEmRq/0bjEh5XEA79H9Yb53mmU2z7Xl5uvl51GioasXfWqbFxO2DnWzrdM0
aOBempER9UijLCzZlubNP8zvl8t3w0p9p0EpsexO3YrdeEFdcZugGjhgnYA5yl2e
ZGY8N3ZqX2uX5VQHfw31BJ3pests8PJQDEAppA8J8cJtL4ca08UlD2zU+mNqCbfZ
lWLlsINuY27+ogU0jisi78Ov8UwEe7737sgf5TW5lqg3q7UeYjf2CZCMetAA+m+B
LEHWti39iVdjLc1WQtj0T6NQ48A85kt1ADep6WoQLuDDKYz8YMvZA3H+3O6En7GU
8bOHI8XWvDeu/sHLqvQTzziIZZS+YYDOLrzrlZGx2r9a7gTTmwsFCAczf/nGUwwJ
Qp6Lgupim9rLsPzRJJ7QkipllIu12ylobEjGRBUICq+1GEFX40nFdOGS5aBNfkxT
oisW7danQDSz9yZPqKPzHM0I5uPzbm6ZtRzVlUnBx2nOHjhk6MfmyppfQG9/2am6
4BabwVmKoI+QGnpthcVV11IDV7WQtkmm3wgH/zWPAelIV+YD28boBrGsrcw7DQjb
KPMaPC9Hi6XGPhlTgQrOwYzl5FEa2vwPYEZNxx4H8cxqDNpRwMn9gY5BjQxeWinb
nz2nAyK3cb/+X9CKE8NerzDnFWrKAmccl/LrdNfoheE7brdEp0OhUVf0oSnA+aQv
45EAMA5XaCaAu3i/h4K1rXf7swg3gwjhtkEl48u7ujxAeNK0MXW+0enMwAJektt+
1G7ZJPB/TkGr4lKGvYaAtI6OtSX2CoggXkBmhjdd6CkEzdgy2Kp4SCgHkwdAKTKK
+qHCLfJ6n1fsIcGXmifLYcrxGrp4fiim8P/yXCR68ieG0iT+dF3NDx8MuxX0s8M4
fFlC1s/Nohjj4TKhO7qAue2AVFb0SJk2zneD5TAjOV3OANE9Pck693W4DJergOqr
GYsbc69fjocpcReC2r+LIalqxMloAbEUVtCrnlOLVngpS2wK6+XIfEU0iJpET/tf
T8T+T6Tc7B2aaZJ77F6iqw0r9Br2iwqaEEPoHLgUz9hvSrWmy+qDJWqCSI3Z+8zA
fTFdwsfZ31gZ/yBYmyJZAa5dWligRj/RaJqFQzlxl+gMBhkSuUSrcxzdlq6dVU1J
OfTk7G0UeMN/NfuayrnSiNvkLi5AqEcYynrcNZQZS9tYvPCJpOFjo0JWHjNG7S/M
2ukQMw+84g044ujaSh2uysIOD+4Yj5GrOr4tCd9QggU++j/HUl4JeqmaQCFZiAr5
/Xr5c4k3glJhiU0dmGKj0zgRnAj8P8ktoyaqmoOoc6YVcBtQopxxo1vvJidJKYOj
mqJRrNPpJEQiR0Xr/hRl3p9fbrvsyfREWZZQBYc1jmOePCNn40AyxjhDgB571ocV
tRsuawxzpQCRblRTPvvaULPzXV4QIsSMpzMJ3WuWaO9a6y6WAT/5wlW4s6JDGsNV
lPD6O0MpEZfcZq7MOYlQthSqTqkSlyJtD8nSGSv0QHjQUIAcdvlGAAdo2EoLeDd+
BURzbGwjJGRCb0DJi4YkIlCgzh9HmMEez6oEavNcuMeqINlZw790xyhW7GYbxbXz
B9JLg3CzoKgUGpJHW9LlcWTD+bb0J5bhbYwVDDVzM+aEI3gxCGpb6O3WRycINa96
ipkGzU8ta8BQzrh15tRqijI5d2z95tB2Pc6MrnA0baQLF0TpYT1cF803IK6KIQpm
rNNIS20+2dxJC6BTZvLbcaqaWN8wahSwHDW/C/9BrgSeKlRqaA2x+gKF07wCZNQl
DteK1keT57Yx70tSdWrjMH0ALErlXDnu7IPvo1vI+ROFf7PtqIe/Wnff3MoIOJPN
RxIKiK/fMckq1noIP7HwRiO+KLxt99q3uy0EQ6PN8GiNuitFE8lnZD7U4BxdEboD
/da+5lrC2t81mZNx0SNJlZWdA6li3jsWtq8GSYuKhj5nMHGWRvfeWyeL5ZKdv6Yd
itKZBYUcBjGzUoWmNd1olo474KvFWap4jzxJj7lleuxvkPzf48yAvyyfLkMO75mV
DKy6Tu/7aeYmotKRxdsu1C9SFN5iOwWxan4F0+MgiQMc+Q9ihdx9ZE6tzNupjEGY
CFVM5VrFDSBh8Pj/8nXLl+6Y3fsItUaVkskKpXiuJ+B0owex0eb/eKhmck6NHkq/
RUG9/IwQVJ6esHmSHyhVPVgZbxi3mDtdD5bO2mxUyFSylutNyYk0cZym1QQaKk2H
RG2CCJsN3yz18b1kVrrT4RGkIZu8JDLYgl65t7UbhbhDRo4ZiTHv3R2sy88wImYY
7tKl/Ilk6xP2BeMSyWJtP7Gilv0QP6h23tS9z7F2WYp979/7XhfooDP6jtpwIu44
do8zm3cD5hp+MTUjJrAduK+XagH0XR85qSpgjvoPH1Jr/powraJPiZCEArYbBd5R
yv3rFnhSq24fQAfQbT9lo3TURhlMngfsWoh6jR/uDxoIVTvBf+AkAfuj6flB5tyf
C6u9iqlLkqvO6tjTn0WZMnX7+QydiX5K0laUF2iBKaLMYJOxdyRSvGVVTW3ZkZHF
HIzt4hMDtLbMKBRm0ULZlE+vLi9Ak+ep6NjttEbQW+NkbA1M6N4gU8DyUzdw4aec
P8BeFrJ7z5wbHxmCsEFVtv2x2sKl5oqBEloR54TaMXYzlfKAFUcKY1X5JuhKempk
NgbffSj2h9ObOS5AoUXtQkcA+XdIuneUuvGT/2cfzkPUFpWb5ZrW8/YjuwZpAmoN
rTyiadZ/0lr0IByvVsZ/NrYe4v/wSE7BfZMkq7K7Seu3KQwdB8whkbDaJ0mksFXj
umv25HrVuV3ZMOcW2/XLgqGiBjbuw3BFi6CDVIf8DFvtQ4QMx1jrvAYbOpNdla75
dH/LuvnbXOwbDBkVu44oojdVWXsaYqIosGgYg/9YyF3UrmqCAl3NYPU1jd9kmhav
kXyGrHF0rmCA2Y4cHdGLL9hmx/M4WDajg+QhruGjyh31QcLxm3REon+xQzL/rLZH
1xZqQ5HjfT2PwoVrBykAMGxZPQ6Ga3sc+RkUJbUeJ7Ta8fwvgIx24+LmFJuQpcSU
k5JD163Tm3qh8I5dfM0OnrRDEiBc7E3at8K69yHqZ1UeulametlBDlwOf97Dya/K
OvhvDaqMOruKGGV+rm1dhr+WV3K0EXQakPBuJC3kfdKSHsz1PRjsDcEeyCYe7fBs
k3UGwAfsPJ+A4YCcw6bFXAwFjTwuipHEsAW/vW6+xd35bORgqMWCUrxwZmu5oOrR
m4afuOjRhv9LjIR/CgfIQ+XWIaMWzV0/mXBvypFyRGxcOF+z+Fhe/eFH3amKtcrd
1Un8bL+IInSA84jEGnK6kHIdam7TApopQKItzEBuLiVrTry3oaqqrHWHg/edO4yZ
1JRJfpc5klLS2S3S03ykifl9d/uqbwkc4b7P4b5jwiVHHMo2oQi4OxSGH3LFtJud
pweiayYftrXaaZ4iQK4FLV1oKhTbjj95TFJuwHOQ7b7hKJCnn9LzSxLQP4qRoM1P
T/RXXR30ViTQuy5hiC5B8AegBzY2aYxJfOznjkS4lCA3zTnAiS0jKAqOPn1DqbSF
TdB54uIIAQ9WTagjBZ+O0A==
`pragma protect end_protected
