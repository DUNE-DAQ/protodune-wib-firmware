// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LPFABXUbdP4ws9xNkxQLOaaRhNRUvrtGF8PQkfYSwN5HgLiOxYhvjyj2VQ3hoq5O
0Kq/W7cZ3Bjb+MlmEMvEXT9Ot2CgmIgUBbnC7UGclXnh5KTbGB31CbwBI5HSkjzz
yya27VJ5UHYufyVFsfYbgD9liwUpLWuGHnfXBgZIoiQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4704)
hxX+fE8b1IxFZXmeAiPB3g+zKAW+r1kcGCxny8L0gFxMQVpK5WwXAd47gLwMOFos
RL1kVv46tiC4d04Ivx4Sz99BkceIYqcFrXEYZ/8YzNwKVILNIwJZZu3FKY/NeSDb
dfZ3qFOMRnqTBezZ8ipa+pd1ONiZkr3ibc/CDiOZqyY9mxBRoJ5BdzWi1yjZ6/QS
oHOIJGvR0rKOYQ0uES+eIuoQj6iibELFE6DuSWQ1kAOYpO8kQ4WAOqMAK5Ed+AQX
kTYVThqXBA1TIr6P32M9BAjjlO80aMkgzB2Hbkd4iknOCDgiThYaeoq3fRRm1Jlw
Bo51a3zFpk3GnPeA8y8ViehJYNwYuldYYmi/QSZOqCczsEa2QqQMsKBLAkyD+ugx
noyZTrIZ7HV/VRUjmY/49VuEprdS/WkCm6V5XggS27MqQB9WU5ZlPyMwxYxoxP1W
1GTB3u7DsI5ZVO9KuSVMeG+80MVXbGsjVojCPPxnzK+0qUEJ13mVqfl6ju8CKdh5
NShFlFK93Nj3S62tGnw27qHP/iTozJfEz2B4ppam6xBEWp19WyNBhmELkuuobkpa
uUQgGir4jXcMZFSJXM/2eDXkn+bENhvnuG5qGaJaHLYa9eq4sFJzTIbZEJbdtGoh
muMl7UlJB1180VpdsLpFCL+RSJ/hlfcAW1T4sQ7giro3wzUlE+A3LYcTf8yRLwxS
xH0qL6vdZeJPC90RI3cwbbecq5gl3gpQ5qGTaxoISpvnTenUVH2tOq8ZF/WvpUoL
L4Nx5hLpws/LjsQLuQh+NLp9Xdct6Kn1keDCjfprzkggOSYsTKcafdB3XOo329nO
+Zt1USsliqpaod8WK9lIKgqA3kp5dDRMhVX8nrHO2853Gp0SFLRvSO6A2kCpUjwB
7878RgZStGb1RB+owPeMnxGNED+2UJqzoaSN1cFY6MbuWLxygQAjk4RqFgSphdFo
Zv1/8bMekU0bZCj/7oRHXhI1zh2ZtzjXiiNSgEqpJ2oNDSNEruB3TjnT4232EZdx
CY8wUwDDeId8QC9S5ZcNHVcE5dOsZ8DsiOzvqZhR+az1NkzLW7CCyOjedfQ84BtA
ilDaURG2gj1a+jWAnVN5KoE0hgDbkjvJIScrzVYQIIKYW8eP3cVsmdu0w+U+auvb
K4b18Ad2/DYPbsctLP42vIo93Eu58YqymiMmR80DGDDiHjZ3O5QR/51OGDM+K4E3
vAc/GWOcs5lrV2O6L+Y1aaPut9qK5yT0kYoOyYWWJ5tTBQuiWMy7JQu5J50Ecb6N
gfIBqBjYyTnXlTBEBXaPpp75+vwCS4mAxVLD2NiX1G2Ua82ZW5Ou0c67fZlpDbQV
nBe60bKUGsLQmR9lRUuaW1rngzdQ+xxN0BAtNTtNV9F/6CGKujTTti0soqGnrvOD
433dZ9kdExKXwSTjZtnS/e2YPvqcN/pXuCxkFkMkpgIw7/Fz2ypn+QcCCWv4awim
aInMdqrzhV0B+wa6B1s/9ao10UiaOmeouAXYtoDy6FlEHdHowbUy4y571mWeOdRA
uTYj148BiB1WpComBB+FMlr7foBic5VIsWKqq09FZ5+ulA01bLIJJz4WLCUabOBF
mX6IB9AlajVZXRDN73DJTzKU0Fhfzm6wPFCqzUaFxcxDJ2rKYaSX5JW9xBoVkCuz
a+Fx+yTjHq26GPG+dSgLgfu+xNqOxuMXQrunhfXqyN4FdclQCSfO3MT7PllMHi/Y
iFL/EP1tztw5coPsUJvQm1xsOlqC8fD0gdhQacN9VbJ6uXpQSo47wlh2jvQ7/goL
ndq1djkJ5oReEZYSQCruj1RmcB90Q5z1QQ9OYJSKeyZMz45eOw9qm2GFhI3nW+P7
trZ6w6HoWtOqblbKp2hGfoF1LqITTzXKG8tt9RBF+jN6iqIaSA5Q1m6jyboSqWsB
rqcuUf7s1ThLHZlFYlINVyM6z/iA2ZRJPKSbNL9MLJkDVzkGTErVqT7Qzg8IpF1Q
aoQIAjJKov44qOxq/g5a5XSMrlshMOudVj3GkEpiXIo9/bPqJrbZK3uQUv++w6db
AJ9C2a/sABOYwPA93lQDW2JLu1Y2lPDmpx30rwnk1OSrqpKIkywMJfPLjzRRa2hK
3sohLupIReCXjuANTMpM34y19WHIgNhLWeMaZ1AYDHQX4OLNNwmDJdypCMzAJl7o
zbtjh8P7P/Xectmy/i72zcfs2wOB6WFMyIvHtoXFqVuaDylju9DGhnYE7WklFNlq
eh/4nfwChAmkutb+eVYaQJnSkxVB6WbrZdrfMSP8xfMEGUhQdHUmMvMqgfjJBr54
idQxgLOLI4/25sgHuMP8pP7CG5qs86JJFYA7n9oT1ip8w4hinPPvFiAbcxCuqnlM
zPMCCMgYi8osg2T1x26+Adx5wOYMKWuxrbGqPIVX9MwXK+2hqbZM2mAKn2qU8BW5
4af++d1g+41kk8SnIZSHK4lIkWCYHmN+IkJxbynMybPPZaphruRdEZiFySy7kY0t
dzPJUGRSoQog4HhfY0d509TYHF++ehqZYbVYZoNGoLT8FOml9GQF/KomBKKnV4ML
O0y0OW6pENd80oenF6eVChkgxQeAn599Q5U1v22iaO+YzjOWUrZnkilDG2c1LVpa
Gc+YYGlzP6rZDS0Rooqw+kv+XZqerDAqIKl/qFY+GQXODLBWQ8kPJt2ThHfoPZIQ
a/BxaHD2opJCZgIkJfOxCQzfysHGl+ZutxqpcaM+wXZu8vhYqhqCOxXc9gGp1THX
bZSsdagjG+HsjgWONLbbpp5QnpAmakuJzYVrzAhQVh3lGvQ36kbYXIFQjKcA6Kuh
r88mw9uzywDVqffnw5/NG1A0NxqsjKyRBl0T4TS+H7RtLQLNXCv26ukkJDvhjkT3
6gEnKv1MYv0LVhZkK1v+3UsFoWcJsh7j06rtScJ8+JjNANG1Qkd1DmWfQnt0l4Xk
LWnUKGwXpTxRc2s2deEWXmh57sY6PVYGnIiUFzGGqIMSS/soBD/BdtN3IZJdRyQd
oNf2M68aqW3zwDEohCxXviWFGrLV9cNxqw5A4YiXG5pu/5skR0AxvLiVlptKXKnp
h/x1/WgNKEoEyYVxpCt0liVkrR65FcxhztqVhn2lC05xSxPn1/KHsAFE5wpnxQPf
kKhOe8sIzyrIpF12H9WQa39qSrPVnAqxbarnaj6iEpygksE16fbIOnIAtimKS93P
d8n/jbRF6HjS6KYzlHD2uMirx21Xw7VaghN6CSsKMFCyqJ6LnkZc3A5Foqk41HJI
uCoQxvsdXpNj3VUqL1QW/uDVssk0MuqI5Vcti8hTiwZpSgEPV0NbUbQIy9x2+JJh
cLLozIX673eyfujC4lifGOPzY8eLoUETCOF+W53Hyl8qcg5r4EviStzLtmfav+VC
sRF+RSNId0e5M9lPIpwnN3QEJYiG9Q5HuqVSY/LUcQ5H37B/j9cf7/B9LH4b+1wb
Noq/5h+mutv8+06lq9goj/k77hhetpBWe2DPwWdl4+KnxUg/P3ZRhlgvLH8UXNFx
J7+PYqQm8zSeYzMPCxLMW8cHw3afi8pBmM+ED4EDvBnB6tgLcbgbfcd5JxOVIwYj
nXeDgHfD948OfPxJo8XWI5AZOytL5jgyo31cvt5ZGqKP7nEBsE0PDklkGajq4VSg
je6xP83GZaMGNNUKWmYJpsOIfQ0yd1IgJbx8dqD1WF0T8Z7ETp60aMgiPZ7STZNM
WsKWyb/M23n3WIXILtHnYgfgHB1GkOTg855/7BMsjyS5bALKeJy+NynUWXdAgLQv
+FZR7gjgrArjTSlq1qpXoSP8nzKho8QgQys2K/wEGog8NP2nOden2Vchgx4Zveu5
dzV5zZi+5UpxM7AVzD6yuRHlZxr49MC4YpOSYpuCv/G1L2O7vrKhyIce+BivUbDI
H3jyVg1hIg5EvUoadUzowhDwAtLriwi3LAeRDeuzduazGAAVPRMcF+N9QOkvBNnT
Z6IqchqrlTi7mr6yrZufzHbwSmV0nJG/Vs+2w1Lxi0A10+oJi6GeWzNmhSTgajsU
OupWf+/n//Er7Sx9ZyIZ7R4JyTX6yjkYjdzkum7tNfYK9il6wFeNlgCly+VshHKx
7YBdCG3X2Y/39EXayY8cD6+3za5jLT6Fr3dN63DAACXPTawG51R8TNLzHMyv7yuI
f8DnlqY4gjTuE+dinwofG7+xBCdG2oeK4HYLbN9uVX4K+9Hjf7swSunYhqcJcpNB
SdI/HktoqbShA9sjtbaJfDh5rdohbDBzByFj56dNkzrE7FuApYuFeKKHFMjCFf3G
9g8vCcgxmB0S4aA7DokOTtOIrxCDJtmVvy83bdryy1nvbScgBTWcXVpQVGLezerP
gBXQ+crRxLvQgA4eNSrNcb0OqGS1Pat07bEh2nbOOJmyHekVyLTpcAuhgD/RChb8
Dlro0OP9Vy9H3gnpYRt3eGqb74TUSg2jsHn82f2raHDNZXiLJK3ByVObGV506YcL
Ced6gW6CfzjIohj8smUc+0wYZUoL1AvwH3rHKU5AKlOCI2LKTJubDv//wecB016g
91q/zpTEXvjgSyzeJDQmp7ZPLKkJV6yP4hbYvxHtxeCpaKk/BKaQqk122eNe2U5I
5H2x8Kwaud59DOiegzOujszGxlbU9jYv2ZdJzgXjvTpFnTO2Vfyv/ULaToigFwkx
DkOlt6iEr2Y57EMihOpxHc70q4D2bAKQFXcZEnQwbL2QZWydBqVSfpOqpiU2DEhV
4q1Bn5SZdM+Hv60tJDfr4BaOwe3fpAbB+73ETvRAkroqLv26rvszjlDWhksm0I/r
SFWoR3+RCWl8jbSV1Ycc9hOZ376gBvSGtPzvJqYKaeXb9MBNX4G4bf0r9fbAAQCb
tJ9HTZm7T/UAwtq3Z195bbrmx9m83qH2DI9LrhwSBCUwN64ZLEinRAasKFnLcF3O
EoB7u/g7J4KZZYbrPgK5BiyWbAlCDKjLvI9W/Ghd8Z1dAAauSnCrisS0JdOySutf
X5Oavr8wBTk2f910Hly+LbUcmEud4i+YFvz52xXo1sd5BHwATvZYOD1b/I2wvmFE
O78NIyfsw9Md7+BDxVhSaIhpLXy12uUnXHlDTLcTJPdUVe6itLqICLt1psCXta4I
K6dcgZIJfKyYYJMHItpeaY3SgasDF9zknBeFmHpc7KMnZmVj3/sEUw4FBtg0Nvvj
qubDTFVhS4S9UVD37QVrWHbQo9L/snWvb5DVe8ZWFlbsPjcr1Aj1+LKpJl+LIUWl
piT2RaMccw22wmS4A1qMQdIzDoDZl1YcyGqOcEbBW/GL6BuSfqeIkzWiA9Sedsne
kfBk+P/qvjAZuj2OZ2d3QnsxZXwq9CJPd67YL6NfPMr4mrTS6Zi8bIrLFgeusbYM
gpneUkP33GAYcW1yf6Mg6at/evWynH9JbpYIj1tnPXL3fIQwk9dBlQQwGR/TOk+K
26gAJLyeUIvfiOJa62wiG+5F/LrxBx5wT4GRb8QyML0amjlgvLq8x6KS936R+gEI
m2SC4YA+Gk0YN441ERSKqeqwtSxYJ0uSdJdXoocnYpyXLl+0SpPDQc4QFN2ggV6D
YhR9ycMbjtXIxqLz8LESy4AsMNtZkrCg1HXYOj5kYrESofz16GnmkD8nc0wBNLGo
6tbV0ds0tzowAXjjoxoLxksgyWAvLCqbHmgcss6GvhYPo62WOXk5xeUuy24gtoY+
kXumtwGQH/AeZYs4z63hvmEA2ZYQHdrH9ux2Yxtfo+Rkf6BLsqe8IdREcOygs7DQ
/W7ySW2O5IqcL/p4yhHXC7HJSdt18n6u1WDPN6Khn9s7BfLjs/zyq+syyFEn1WUJ
Dgt7hEI6PtC8AgYptobGOV7Akb0GK505qgAxZJdNnrIfGp/1Cg0EHQn5B3uBWvWA
Yt5t3/O6vGK6KWdLJ4gxs0/QG52PVjWuIzG7VinSfw38K+18Yt743bsDJgOrKg5+
qdFz7Y2HkKqby65tbmfUYarj8R02sDSZs4RdQQ3H/KWN9hdkvI9b3HI2zT7hvrYl
VcD9gkFYDAMwQp1zeHb5qvo2JNd9pDcdrjSVGvb216jYXasxlbk5nBVYzRSv07FJ
TqX9oUtuqjMewH5OG+cwckrdtLBjDoL0tLA4TDWqzmpjpjU8w9IwK1O8NeJnM6Rr
hn2NDrlAW9+HFxcX0dUXJ1nmz3lhwrWCUZpLj9P1B7a0lWuhXXWtF6fg2UQRrnSL
sk6RGZrpwltnVPNMPFQqShEKAdi3l8DwOqo+TxC1JsdreGZoTZSuPk+X5XUMShQR
`pragma protect end_protected
