// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R+r+CNm+3mZSYMoGPU8A8uDO0njS/JSWqUjZUBx/WXSdMiYKiSWW3C5Gm28g9Jq6
hnKkUm40A0AU8UgTIybOy5MG/8sPT6mH/lZy9tgLZSDnyi6ugDJ+b6VXSqqVGZDo
GxTzObIHUAWM6Zjnz3OaAbAz2+W9p4UfPTM/xzFqvAk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70016)
NHEH7zddXcwJjrYho7q/wHRhAoJGgTTT7bpVfN3tzLLKvvXszwO0hjoR6trF1lTu
h9K6WQvbCEHoUNJ8yv9wmDGe0RpSSdesqdYzj0ZU1WMI3jVLyTkFP4XgCW/mnz6b
DJVOqRVDFvZNQZUkX88NYZeuZH7i5G/poF94uTmjHTuRF+RcibDQV3Vx+1zO16YW
bDtqx7aoeFz4bld8SbfnVUA88QnY+UBgZ6PfV+1+Cka2+FICbnuaPBoO+yYSwN3l
gmFJnjzdCcuIOiLu33PGXdtRZIki7P5U7bcEuhJVDz7FG0L/x71p7ywV1lEztu/q
tUNfdfrlPp4FBu89fHhFP+gCjP0XHxm9Txrb0v2dYVuj5JE4ok/umc99ebgtey3b
eM17dykdyU2xmNC1n46ID1F2+mJjYgBYPfS1/EN7kgTDV1QrbKUuAyyy9S9Gx2H1
BZ+qswcMqy7vZ3No4hUunEFCoot15sk6GiiXjGN305Z4fkaK981+H772ZXoe61n/
or1XGv3WqU9ERPjZvQKlaoBSyQlqApYrdXmkJyx+pKt1gFZjojm3z5I3wEfDwQ5D
9tcbE3VB1lsCihOk15cCU6qmJeNGw/lRD4XuRFTGJKcFgvkujGr7zccxRLR7invG
yBTFZD5CXjlDz2RbdCr0Re6UlTgzUtv4P+g5C3CLqeIT+bjv8PtYmBNiSlwdI5ft
G7pcNDjCAkK5ZfcddDkjd32JpQpO7IrUrJDiJOvOrxFoEGxAdmA+R4lUAY70jByA
NTcDhg1TYvkNQxd77/6jRwJJXJPFiQag9mCKdLAiFArno50/MDmC7T89qpO21RiR
konSD01PqEURoqM+czZx7a1WJQD1CpTV/tDZEe4l8Am+Cp7GQ/K1M5x7bMSLDPPY
Om3JRJM9451JNRfSpBWoLN0Yk/vVbfZMjeFpzQoJsbTaCkUkO/VhqdAiApU4jrb9
Z4og4/MNnOnVai+mrRdnQkLKjr+XuoLz5rVoaoH0K83KA2zluQnspt2PUyhCbxV3
He19ZdGsgwDyCRl23wSltzfs6dwqdok5VSBJYE9iRMvMcZ6J6mpNS351E8R4uMRI
6Tjt4PpbUx5HeRAZ5qPKNzYirpUGhLnkR6GlpkFLe/l6SRqNMcZEuuqMYqt7EMeI
WhRnzihoZzTx197V8WTKh6V21XECqXgaBswfWmY7igikRqHf6DqaIdN/hLnZB/TA
zZEyMVavXsFIBjHd/9emmN5gtlBEYOYpjoAUOBB73sKYiH9Cl5suZLi7jJCJqgIN
zEqDuTunapg48avXKMvF3M0NfBpQeLmw3F+LwY/tcDI4XNqk0nP3E0FPiDr+yWsI
dFVYn42wLY+nWfOapkt9wmCuyyXMr/NK7Ec586Ufc2o6OSzqOv9WrT30D1TibMPD
dhmA8TKQ48UaHfOs4cUH1X+kPMp5PrQvKY0EMAyvaqyo0rSOqiHA6NrUMc8i6hYw
tJUJ9clzwaC+HIPSqWjal+dA4i1Ny49umdQje8gswvaPGDPT+bo9Ki1nimeNIFUI
LzWS3Be2BUWKSCGpcZEmqTjYdVhWud50DEzaF2VdTHlzxTfDULFfyRG4bNvn/yKq
AYhD/UAzEhoIs6bSfSdbz8pMMF7Sna6clBzI+eoz+8CbAuTb1dmvFWJQYUaMW9SM
hT3ohaVXFUfK7FcGJ7iYteQch0d/wJyKAEiPVlLonLVermmx1mxErhuENUdyCCWy
+5tutTXwAnlwZZWro2540nx00yQVJYSvL8upSwftuNSyBnPUd20q/K1SoIpZhrtH
vZQ7cj9l6RTXUvW1mka2ZV06my6M4iMJ/zdYCImvQe1STE4c3FzGqVrQFmhLgxsS
RG8bKq94WnlekuEmkxBiMY2YhKlltCwnY2qVsozWTLdgRRdn4Y7ht1wqgQ2RqViJ
Mu5YWSMhrtE9+wGm7xmRLS6z0q9Qb9R2NufE4XjLmFf788XTLtk89vGR86UbEGzf
KTSElCRn/0vPPWjeRzDkIhoBlLMAVXvosMGr7HASL5n2vmpmB3W3tyD2oVQWVczx
16TO33MTrOr3R1IDdWhEV0WLe4so7BWvzn2/BCVajSOps6YZ2Rn9cowat9m5feTI
DrsM9YT2XzWVCj9nvbWzctfP5fDwGbSkS6LDXws2Z6NqhKOkxTIdxLDMLuOsQW6h
6tjgwh72Jf1Xmm0YQ46CrTEEM2SuekYmlajPGAzVByx4616G8y83vVVxkfeCSnSu
Pwhd6UWPGTW+qKPt55JRcxOARi8svBZN+bWuwlquj/cyD3tX70g2esfklsA9BFAw
GwLoHQ8f2vBDiVuXzhEaX5RqwTpDvZb19cq+B3r+WWo/cg9AisGe79VuxM7mccRC
LBaar9GVRIdiXToi9H7uMD5noffe7mkj3RSUSdUojai/zc2dYxNpIrutYVlCdqFp
6TnTyvUxJQtwdgcwlXXuXkbwQW24Bazja7DI94Xb2MDPDrLa2bri4fQdnst2WvHq
K1SXxn1jEXZlNobCqfmlmOt93+gcMO51ZHBbqCZc9ZPBS5sA8HyhNjjn/XNKifZB
0jvdhOJhfRNZrLy7C7Iu36ngjBkK302Gc76muhResV/LLF28KDLi0QrDzSpVLYH6
JIuXRNXn8OcOA0JdN3kghBEpxhs4oKcwPM7gXIs2xMuixxOULZUM5w/0yzUcp8Qn
aWVyVopF0TrDWVTx2Kok0KjDJgBwAJoHdOuZSrRcVXoxBr8FKPlcjuNogMB2KJc+
o5sIOMYBWwK1SIGdTyeejwMwdORyZjothzMsIkHHKqW7GNV3b2+ZpwX+hs6d5Kr8
3a4M5Xy4Sj2o2FvAhlghZAQ8fr3X5pDXp9ERf1ujJ3roV7h5qlTCKvW/zxFQnEBm
2cjmBAuuuNvOXGr3JuolG04/79fPDd1lLckSPWTY3unO5llMcXn5ELKr8yYfhTfa
tEvNaUEuOpIpHc5HK2hB9qnnWBdzjJZ59afAm0GBGGVQ902bxjPsMMfOyGBGpHw2
0AMrGfeS9ajEl0Cs2+ay48Xi1L1sOikGiDrSQLsxTqwf9GrjqUKuLGyZ6v7grT6u
Iw80bWA9JWUG9z+UhxeGmeFVIkjAnWNiGjqBnp8EY0Ks2CQ9O0P/eJ8fjR4mjKOl
oIIWA+hbOztcIPImhEhqr49z6UwABKzCwz+UKLUjjSrQbeep+yGty4KH11fKcOMl
cZ+PrGUIJgDpFpazcsJttig1HHTsggsDI/61yM/irtEogfLZ0KIRHGCHNLEjgnnF
uFJdvW6lO//B6Ltsb5O7oJixoYRCiAf7OIlJHhq++M79YOJD0kiUPprWn9yM0mad
jNydYcmsbktakev1s6JccnSsYe4miszaVE4QFJk2wsISSJI3A5sBw4ji+iR4qwb9
vQy2OfLSvFXyZr2wELLs+qbBGo4wOd/aFDTHBvhkMwlXKR4/bqeACDH3WGP6P125
yAeMuKSlD+3DQAJ6b3xOxKjoqSKpGNiz25skmFCK+HuPpAaWuviii7tGkfDiR+99
SxJVpa1S27e0/l2iD83sNYyuPwOexNfA6oO7pd/cb/BK/SIyyv6DsAM0pZQPXVPn
9qv3fgJpZ1Qkec4nOdpAZE5tX042Jn7TTn2NnKKyPlwVyjefcXUWxvEuAlRRQt3d
79MBlURgsK4Loc4cKQvxZoGaEC7W3VNlVahawhzdrjDX9EzIv4MbZVINpqsk3ODd
I6+gUp/e/6xGUfTFXhsgIoEvwJMbTO+sqnQskjX0FkD015kfNzetlXBIXgRVtJ7c
AEIzMgcKkhIzlhTIIUL7qMs/YxMz9ofo2aTy1x0csIgshfOXOdoD3jNk8CH/93I9
WUWfAmpm9oh3yXMpYknRaX3DBie8u8yTzZTczzTbzeGeo9V2K+DIsXQAQ9iLIVdC
oQ5230AbRrh4g+OCz34iAH42W5biIO6L6b1uPuTjd1os9RcQFrR3HyEFWlrIfzkl
XDxJSPuR0k3ylPJV86Ov29UXr0c6iM0QybgEboUtDUQ6pybYPleQ/DqGXtWmlE3L
lOZoo4HcdZStwX+m9nUKhVZKmCdkkuM2a02HmdPmg8yfFaycB1SwdlXLIty7GEfA
PDbFJ8ngayVV69WLEDH1fuRdzQrhzxn8Z1KvtyX8ZkYNzMyupwfxLODt2T3YWhCV
ES5NmiBhdln0DI1fB6rhfksbNJSSpdet4Jl+ucph0NVBm3G6zN9l68DbS5AyvzhW
Z4mm9Q5/zprz2RyvdhqeNhpEKxu4Ok5QdWf9eDw0e6wOTsZ1E7TM2FdhX6uda0Xl
zwEVm3cHokbMS3vL50zA7Qh3ImpaAGv1tTKCq491Ew4Yz8SBEU492GeqapVKIMKB
MH6g5g2pLyYZQsRlPVxRtwj0w2Ir5zTSmDqv3R4HQ9sqgN3Hk/Hfg7JsHTeL0ZuN
uv7vtysR8cUjCz2R9pBLa3Efst/l7yOUn2h/hE31y0H3U3YgiXlTwMMxT/Bod57w
41CRQi/cl7WzqLXZKxHm0CsGD00dZuZeEwuwRP8p6VmEhhU+4fkjiKf0VB/+1h5/
LK73REB+M9QJlS4HB8FNe59QaMmvBp/FkamZD0wG9pcU6iUlcEfoGHkjIe4VNNc8
m6mUWII888QKqo14eFXr8/goz3vnnmKPsfcMgKTmQh0QkkAtOf+tQKz5fIrjM6Jc
oWlh5N0Nn/2NMafQA96dSUzyxCRK+frNd63bHnyxwfrh19NJd0j4WFiuOkRX7Sx/
OTAzLhSgbX6UxNmtwok5WxgCiatLqhGlBcFrOshUamcnTfreKRDqVj8P+JxqJVDk
+MCfgEhRiLZcAT1/BjfTl5I3d6MPnF+1pGwBqvP3khwrjSGEqtvz2RQf4+qTvKee
ERVIMB7y8qNf0kvskt/6GQFnPXbTtWMcTRTKZ9m5gauThBxbZ15Fv20BgN//I+jF
QDX9DqYZPvisAMu5VnuqtnxUlV1szUq8PJxSwRWdkMb5YWdK3hLfPpqHFEM0ZTBu
gP4Z8HoA4gfMqI8GCOSAN5++cBn+dMiT9LX9KARUpLIPvXoF770cmGM3J5/RhGes
1z4f+G6ufDg2cJHizbGXMaLVSrx0KZEKatzNm4bnkpLCZZ7t/WBtPdAZ3T6kectv
4vCykuAPRNy49BAf7ZiYqFf4KozDYPVfuNJW9z9d7qN9sFLIH/mXMjOj2nB5vp+3
A1s8rP78cPhAQLH65dkV/91t6QXctexyGllkdL/fNa4gHIDiwz/+6Y94OsQXjh8F
IDogBRfSTP898MVWPcmFqJiTJ+rk7fnnGtCCd1KA/kcrnNUp1QWwgl2cp4V2j4qv
w5K4Ny4PZ6BYJs6Otvdl8JayGZAwym4puMkBrkWItG9XTU53i3d6hJNINzDQFqZ1
ZEkM/UcvTaOZSPO5mv5nGEoGuctEE3sMBKMxcxYVq5ooDegUeQ9+/wtrRC+q+3Qw
ELRYtMhgZUB4JoFZMGV7mqyWfuVeNts16rtDYiVvFu9FI8fkm0XJTpervAq7XvuB
I5eWzydtTiEmeFNrBucXZo6utRzSuP4ggflqqjT4HSu40Xxxc5AMF5MpXYm/1Ctt
xSSKpNvVubWigxr6JW6xxxk3/F/ffoZXEENXaysBcrfaaeqnVLTOO679qMgm41G3
o76XI21tnyXry8AlOAKB6ryggWamr7ZCDAtvrtkz/CKdf5CW82T1G1EnCOOyneXx
i535QN3vUa8bga2j482hF61BBThmdu7f2YRK/fDlaLiXsyC37mKcUvbQrCssDys5
n9jXADfUcie45aMNFOiTN2gIsPEnPkEKk0WIDqk22sOp0v4/aG5Xa2xTyZT0JVIg
J+WkkZaRgftAiNFUd59x/efw+42FF1TeSKpNncnMA5BIQGmO14XNFkULBz7C/mLl
vKVswejdI6bfS6IPwgF8t4os+TKVPbcNig4VScoYGU4eV4nHjgAIuQ0rvqJW4ufD
pYS2lBoLj/yiOu3XVP+G9XrJyeWaDKvyWYX6AQxtHBfu5V8+JyZPhgJ2aEfucC+7
tSOIJ9THnmPk0KRNSsZHmw1/NhiXNLOYCcE9ElOnbA/0jlG7LSwHXpRFVrnfuGUn
ReuszkbPTQnw/1p6ICIo5K1oGkchZ8C4OWhJVDrOfs9MzbJhdObRyWVbyjBNEMwq
Fuf69xraX/aLnErXk/no2xY/LL8lrI7qxGaXNOnsfNCb8y5YnYh1QIAozZ1PIoYE
DBArgByU9gk0Fs5vUzVtUSrum/Aoc4kCLesmCnISPpXlgC9AHUOXSJGiimaiF88Z
UReDiIa2v7nvOkySCOK6OS8IPzoxLb9z2jS02g8LaxxNxg8hO33bAcsCdKqzB9Yj
j7DaY00OQVr/nkNX11ZdzewczkKLxwKIKzsaR0GFqSZZTlFzCWfwKpL14s+R/fGf
ZwzjiVsr3nWjcd8Laalx19byygG/Lre6rlENrDTV3mMHlVQT9y5Sl1KWUkaQn7mv
AXXzIf/uKDlf+kSxiYYMJYrAvIFkTWbcVvR+QFDCZDNhvbI8+pDOOAzKhIdJWzTz
RclRdliPbsUGMje8m3Yr9Q/YO0Dib7oddndNP7BbzJkv7JqVhTr9qhIQzmL6yTUI
mSeSb2n+SgFFiM3133t4G5VNSWnSiBT212xutgr5uX7erh9DPbQ9+RrLNXTp6J5a
wCrqGVRz7+VM89MV0eYbWa8EyUEBNWpWkKlSBChSZ3CGqCrETKH29w5/SYDWiSnQ
hiFmMlqP6MvaC2bpVosrNiclxoqHQatAFNYnLtkqDRwZ1FHEShN+eV25KrVh/mOb
b612RwYpYfvIMPu23J34LH5UqdPtARqWpz265FMTwh4i6PWPZomhjoy47y1EfPMq
QknzW3ZdSAXvlk442KvGpTISXT8exZNrHuKFAdmQB91BFCGfaMYiFASPgfq766Nf
LidQ0L4uCc/rvrD1u43wX7GUaAMq1wToY+ybzCiLLB5DfQOy4VoUe1ljDbJpIM67
/ftUJa2aHrnUtiD9t+nQU5AK7wvtYuYbIjLyvRnRA2yxr7+VGvxwn+up9Hc2b9PB
/v/HbltZiQr6SuS7ZShiVrjEv/bywXll7ggZoSAQWVxAzD3gsOB7qGzi+LZVZDrD
J3aTO1qZSFo2/+mId44Z7K5JuuG1fv+N8Fx7rYK6muXeG3eY8FmKHZGT47ZRO5ZV
owlUmZ1iIevt3AdsBCElhXfNpPQ4wLd0IIuwc7LCFrruXO4RDKcy7T1lMlTZwRPT
zzsWxQijX3FEnADeGcZJv6lrzM1zX7koNzNkE/bAMlW0Nr9OsUChC8ZlRys/7+4N
4eObqJza1SUsdKioy/tGHWE01gQ7ahSCwOWh56JAh5To7DZs31bLMNvNAeyWBvnK
NuuXQ5qu4d4Kl+UpRaUQ1G+FEP82arnPDh0l+LE0QZ9hpCzS+PBH4neI/JGy69oh
CsoGfh6XalHcP5q5289WQM0TZxmrMp1hk6jlcmAl0xZPhSCQD0gvVIihnBQ2bUAy
apaLajUWCGu/CrFnhvGmnZ91jicCqQupfYo6+okGKJCvhG9TANFmZ7oDcw24IfX8
7imBnYU+JB/1IWJGTYQ5AC/UgpnXKDfmZ8D0B7PgOpApWFbGlKtJ1ZOBtlQIG1Dx
B8h7z/XXRDFs1pioPCzQIeY4iG/DSw3gZNeKsb1SPB8hqANi0VyF00TT8IbABgZr
1unedeIbhfHMUT6PrQC44JaA5exLiBuHpS214yvV6MDKRNVQiJhKcnBjf6PBvO17
fBzXshuFIo0EJLRPGoqKl2wzraUdt05mSKW1JtdSaQV4FecMhzCxllaS3HnhjiXF
teblTkLEXqaEsILS2b7wA3JQprWKTHLodsEVx6A0cufoaZ92qXEVZldyBtcu9T8P
x6nJoPGMmwkD9EFeAcMnxEIaCAilfigRe73nQ9a6iLPTA2BMPyxKJgGjCqA7bHlR
r/jFBpaunf+geEaTPHeNB2TIreECv7VklVPcxF60ub5lpsfsYJWmIWtuZWuIaFBO
bUicJ8Kj2cEfK2Lg1Du/o94fsL/Ok/cb2LegFelNmkMjXgUrKL5MA24lofHqSnB2
YvJVkSEappuAVjmQgUgvOCUyRlKD4SBbn48aiDhP1p59Ht9yBUSma7GbZzBV5FKc
rDla9wBdwNSEWNP8iaxN+dMCvostOjfXz515m7lRhwrtbyi4qO8IePvxlDupbZoO
tXoAY3TMuywdLiPO7xzREp8uDpblW8b0/egSbNMDPx0Se68PZWJGl5YdjBUBefkU
jw6yeVMUVV62hlmnHaDyo4jjFEXVshh76UzKKzDHZNFdltaQXPFCn1e0hVFMHmNP
q4lr6otpDq2nkK2bYJZirj/9JkmmFUUgsBCFVIXiOdjVCAaH4XnBFEyCR9M5lVHR
cXVLBREVu8Heq6UoDzPsOGNrUgEGjHKjZwg3SCdHryGvkUJB9jPCuGJWWZzTom+U
PMQ4SNVeTxqUw4r4HiGyTt5S2zpNkYVLdXoIaRbJm7x9uPiqTBCXiaRj6qlzqQIo
L12bqaOdX9y/k5y8pW287v8gI71tYgZDGdil9P0zR0RvmLCakNMwAzkBejkclmMb
+d3z88Cz44grDzaLjwCCuI1CUMBKNfWxbnslGP/6tQ0wn9Rtg1XAg9QQHhfkhpPy
/im74SrfgEtwgAAtorBUJ4sATS/FAiijm1FrJJHEZvXcoU5/o47+5voBDa3KxcMe
g7zR7S4cMFWJU10FiICh02c+VV9HyNszmUd/mQEYddmIrDd3EJkELTePhVvjmSOV
6n8sdaohKciDL95QSQ9v+dE8MsropCf20tTe9FKJui77GvWduwqGnlEpS/pxv140
EjEU3FGKhcMnyqyvjjHzHBkql+2usxC/TZJlE5cqGXzHoTexPum1DpOLdN7igKkz
L/N/QL7zs62GoynElZZZc98fSh9f4O5zVC1Y+yjdkB9hyKYAVJ6vnu5WqwICISTj
+H8xRFwnmg8F3Ms++YRT92bZLJbX43NPCKiHz8bezUDxhQk+2tDKX30d7HXxUhoK
oV0tXL/X1sEL6oNT5P71N1hKJSHqt4OWVBDJPdU7shB4Gkuxv+waK+v4JfPokkWP
foKrd4eQzn0YJdJpZp69sXD4RkW91Vqcm7LoTM7ya91oGwDDHMCuyWtGUPtBxvXC
SG+3fdY+xPGoJI5HhylJ3OOOn24kFjOTNR05tzAkukvSktqWn/AbG0w47tvi6+Oj
MpW1UgWZoIVJExN5AxzBtvHDYgMekKB275X9hHiUttqMYGqpUIAmVITBrINRmtiv
QALfxPZxugjUaO24vmI0IDC5UoFrAKNowfj0zOK/baoZHL3sPBlK/r8DRRINnnfe
5p3/nZk2oRM9fURYcUPdejuGP5bZ7TBSzshTZ0Am6tSbMextjBaJgkhaKODQ2ivL
EIpmVMjO//DIrERE8eJN610KHUVRicTpa8fdKmrh1CU+8TFKOzuDI6cFsrPrtes9
sPyzcb20H8pPcZQapfuRz/JgaLdGjsoZuA9KhUJWwodxT5Qk7cw/tWtZtGqDXHgi
PcIaRhkLvB4JUYfPYjkQcPoI4Jy51+NHaUtzAPKIz6GJVIoFaNxSD3o2SKqDl55x
oiF6KUjPObFF6U8YY2v34F+D4oSA871M44PJ1qY3sZBCIXt687BGQCvqGbeqHFGA
B9CEzQseTTPfXJVSLze0V9St3qEu1VlZmL25/16VjSKLQoIe2S3wk87AGx4ovk/6
qgdtAJw3bWUHYey2aCUfb3j1dVuaF7MjD1LOM2hjZzzRHLiZgYQmJe8Y1j4RRkAk
a4gDCPKsDXV/SOh62K6fnOW/8tN6dg6FtDND5CkpKOXWod0Vhe5JL2onatbzjzJw
Qg9JB9AuXkkj2T8sRptVCIC45CTY9ik+LRLLq/KbHQmZB/jNowzSaLrTaAkWeHql
zb+xmu/G3y5vsZrx0ufSjUoEbbGstcgpSZOazgrhF8+eigR4VaVYykjk+1j4hLFm
TNFz7Dxxqk9QVv0Z9HR0rgisNUQwalLoP0u30dgvcSamR4mE8bojQ8UXZ7QKEcz4
F+c0dZasfBwYVWsU5eJZyhXoLhRl+1OOK7ZEauOf+3Fhp2BDgda0Tkb7XysiDfIy
+uKwZp3svLqV5z+oLdy/0xVfB+hoknCkA4mmmgotblfqrm3L4u9/U1Y8p2FqgZBo
D0x3M/sIV92zjDrEpQbAzqFXtp1P8nrpDeO+LP/ocLRmqUEnaNsTynROoK4qk9d8
OubEJuf0gyEUx8YpioDiAsUaHi0+BHlgMnnPaCssGM5tq+jJbSBYnGClh3mxXnLm
I5eA5bIZoNwGcPNO7JbMYOJZtxVtR7b1uCOnvm4VezUVm/KdJS1k8+0qERBbCz3h
AC2RrpqCGpWgTYt1odtLxiv8lDv+4FGR60UGNVzP/6XV90CvrNhuptLPTwuDX3Rr
PAOPjVF2IKmuNLNKY2qrhFK5U+x5cBa0LrBDgBWDKR0jSZKQjq26MbYqSh/OoWwP
c/RkyrcSUxZ21hPDrqJY9M7cLVYkuK4wKsiYiQ79cuUw+nQZR9qwqBxXo4SveFRl
FnA2hpdcktyYz/5astroVj982M4htx4zbcBpiGhChkEiDtLS9XjIWEoWvAJLUrIL
yKouiMnK3Xhykm6w21m/WpAjNw1FB49zbq3Iv6LpYC7y6tbu3cRWjEDAcKhcr/Sl
24amiyZKXtG5+RJ4fT29G+CE1S9dLozyTZ62A7x3vpUZKbZzemgOgaNhi3/IONAT
NOvmv/eOXu9p9SUyYZ+h9RRbdhoticXmt+O27c2EvMLfXYcfGORNatVOxzSmnfze
M/mZ8BqanhyMQusmC/rcz+Hl+QspdhuExX/g85Wt8E7O+QO9g8q2Twf+NT4NoxRC
jz5UzKbSkbJxw2fCZr1dRho3mfhFbhtlr9su4qLF9D7W+ay2In3f10rgxnnkFnpE
b4cTOruHik7IV/D65cyn/LBvyovcReFX48Ac1Lnv2Mjukct2K//nbdMvkuEqUa/6
j5C3/2dR/nobL/OFk5+qI/badqsjqz4XtnmYUXmX1UpbM/YMcT53uQM5gyGV0JUo
3Df0Zi3+VelW+yDX7Od3lkUz2ThO8nbbSKMbT7ND1wn0E90usKRsSbhaxMrO0QlA
o2YaOvGARSHwnLVpZ0FPp5w0dZCDNGcufbJWVi6xIB/QhQVdSR1WLfdQ1UiBmUrQ
QnmXfOY43T9btA8BfFxg4UgIe9PJ8xbju1KSMXSN0RBz0KJbjZS/5OtO+XFXK0Ra
0fcJiSS1L2OteCyVlkjxwXHaOXy8qMj7IWeJrh0RiHspGYMR7X7pJKolguKDkZ0Q
itKOwLgi+hf7/8L6T2O+Q3IkZWvi5nyfBdKn+MDpZ1hXxOWQd2f3/rybbrSXnnWY
I2g3OM2G2NqABVMwH1Ifkm5+9NxMahiVNOU55v84sQWwYm6iVKrkxI/pacEA8bN+
OC0L8u7JCv8gczcd7jIv7izEt77sJ0IOuk+wFY6TaUSnrpbjaFcGAC2JEYNMiRv9
Cb0ck5Ppl/vyvEL4z110+GqWvDUEDvdYjqUAN6HIyi4VjcWhDAw/8sve3jbwj3Q8
XW4v27lcmOPuOEOgdlg1EauGHLX0D7QTlYhpWkxO9UzbkKBipNZj1IVot53uKG5d
8qw5t7Sh9uq0eCZG2trISD2oEI8KPcvzTptBxe22Thb94Q6DANAsneXJC/ccodWR
qqYYo0ZkXbJ9OzfEcgdTv6t31O4W6lQtszi3O2Wzgm0GdpAkU6e7tIaZVPY8PeG3
UqfcePpCtxjtCqiX3XKQl7Ln9RNfMkICJyMFhwa+v/kE6TGRkuuBbRl3xQRW6Aoy
cFkTFY5O3s7akSbtKMSZ8C29qjCTXlt/WhDeHzcnb4zeAdJkfAFiYms1vy+KdQDk
2UDbxUaC8Y7j6+KcSAyLpS0Ql3A4VWkOdlEryGpuCqfMlgBgJz0KaaZQRO3LtpIf
JdsboeTMk71gp8vFsfjijbi6/qvffu7S58QGQ6KcGZzvvKiChVACGRUDlz3hlDlC
kUeXH5OlsCNn7yg9Gca+zMZCvBcE90bRcZUsH4vz9LPgLdjWTWix/yt+Ob3ikbxg
rORYdCMo8AL9fMJ2IypBsmON723eKR7zs/aLg6tVIt5uuNoy5Gk489Zov6c855pq
GLonbjnPipqBRAm3IKZJ3QMcpislpvo/Tk+xMhxYhfrNu8fvX00qt29r12zxk1gE
R8HWHhx8fBTmxOOC1j+pFFYru6Blfwxn5pgHONxP9SQx/TMxhI/tOj9RI+Wqub1x
5sAOjPPWsFI/U3igFKvABWg+AssL+9tK6+V6xgSPSwzur9usShIlZ0XnPWBvSNBG
TDfE/AeR/wco9OmFLaYLxGQutaGvuTad4DxO2wQRkKT+qlhTmnYlQW6wE4UtZPkW
3qZ/harD+6+3fMs9dmRPN0nEiXWPL5b0j+xa5/WPGhzmrrgcDB31FV6xPb7W1Y/h
ihMtJf6x6lOFokR/gV1WeEb7m0Ma/l8lLgp7YzevAYFlZKT4zel74UjtvddfASUa
MFIEWWOTfp0V7kva61ko9De5IA1vof58iuw0wmJrCEaGqLV8hheXBvmGWFHEihGq
t5wgO+UEyyiPiDm8j5SsWBIac3d4Gxxb9HY90bNuqAnUMU3q2oj++ufvRwI8lb31
gGLNI12h0td4PLZ4y8eFuP7C1EfTJNV3bllN3Ed9eSJTaT/hGdyY5iGsSDB3xfx2
8cFNny203tkHO/XmlitbusLYnZFKsydKgE+zHcV8xgTxclQW82GOS4x6cA1YDV5N
kzo1B2l2/h7pjvJrp5Gdfanrx228SiafvobZ5BtIJ1nudhSr7APC+9OoUV4aBTJv
7pSELsKp0NBq7msZB96UAMUreuCjkD91RfqC5/bBGDFkeDRAq4wB8aH7/OKqhYlI
AORGCTH6cKA0vdWB4b2ScGMbcXRVUkcYjrBwpg5TZg4PBPhp9BfvJJt2JwUQnR0/
9hCEhgHe3McummXnaJIRUSb4CpP+b3czNREBhNn6GfdqUj+fEcqJ/0uOhf+EbCnj
iG4v8pE9VIvxh2v4J6NNX2s9DeMAnoJ+LdxsVO+kCJqNqKrEM73pwQ468gDxotON
Zu2Rx1uRSau+1Bi6d6BbfPOV0XAMgHauUpc6Gsdy5nf43+/7eDK2hCq05UrTKOD6
ZTOfAc0Jn6HIo98oG5KWIjtLgDPHA/J2tL3+VbLmvNTk8tnXanmt2gY7eI0ngwLZ
5gIgS6EvpKbb5n1HN7uV135OOfXPIzGyqKHCskjqihKdcUS5+BbQeRuA5S3JILlj
3hGvNm6Co+5UpHr90zxkdrvd+qmu++RiWmdj1BOzdjzw1BIN9uSKPDTfgSfB9cJx
dx/HBw5NUS5xFv9mcqoHu8mnvJetmioYLtU4SdMRTlESgOz/2S/D6lX+Z01FnPNN
zWv5500LqPPIaniqyQ3bGYQyWtaVBZojt4J1BLmOy+Xrv02kXHO9R4+J0uXfBGkD
speauOK48xpUzAdWGymTSrtJdLZ00gekOPpZgBxS7e/YVALz3Bfoc0JsieDhNc8e
F4F2ef2u693GgD5KSH9Gtfb4zQC1nQbDOqKdGjxyLc/PmXzjlot69Y2/PMVx2f3k
ORld531laafHLKHcjl377JoP9LabM0dFtuoMGcfW3wTGOLukxnGKWwFHweNiy6IT
NoMn2dgIEMLIBTMrkbg0NBG6/Ib+zywn5gbQ+B/WV8foTuFMJsvk9/b9mzPjlyJ9
rUp6+L8zTv/SqB6mC0HaAwU4cl/zVQhTUjJOReE7itLNZQw/9/GzxZqXhf0AMbHx
i81wynJp68cJvGggln3gwrWYaa79/lXnp8Hczjik9bHwWnys0ZJ/5AP4F7Fb4/7k
BYE7Xa9Lvndlv0Kpu5L4Ti23O08CUWcN9R+nfCXmNk3quaiWxIqCBHAtJMisbhbE
h99Ls0Tfzpsqj+po8+AEsbxUpwzeUE3gdui3/O5gi4pUSzZw0nAwS9gjQYId5ruM
5rxtHnEO/frKLkxCLHkXf+Bi928vODC+9nx+ufedi6zDqvLpl5Pi0id90s/oeAqA
TGApMDxAcBLREGN0qarq+UHztAZfvusq3gVM85+SznpkfE8C43BxdFirUR7JhwxX
7i7LVwJ5fLMODnEeV20kxykrBXen6wAl3tT9TCXVPxzYEPXlcKpqAhe5e9uzDKFY
x1g735cdKaHqN2r0rKlFGbN7la7/6s89F4CljRMe5gXFsagnyw8/CyERvaeCsGMu
/iXZ+Navif98Yz2Lmt1y1gb7OTaBP9mCbCJXRhkKknkD/MURqJWo4JD9iyoeKR/Z
Fw0K5hk7Hx1q2P4frCfbR5BiNj+7t+mMVZw7eUmbrbJRGgpw1xOggzpMHTmtqJMc
k05Mk/uJr6NC2ZSTMerHPqkBEG7egf3rMOXK2gsQdv1bhaY7LV5iZgBfMAsUXk3Q
xnzfAikB9YDB9Gw/16CxBKNd/RytKza6qv+bLmtGdOVpYqUM4c2M6DnkWsJ1B/Xh
Vxd9mTgf55SIQxvy8zVQXgmnVjdeZU2I/z6QmQwZymircDfXnjzU9zV+deo1KcOX
pkbFngvpfF+fknbFmXAlzyL+aTg0IVED6KMNOxHh1QNIKRWUiZSf4DnNYxnNPMKX
7tq+rNVo6vq23MqsBfp+wLIlIhhPDaCl/77nOSODEFXM31bfRKAl0k3v5lCebx1+
aXj9hL7oBGXvCIC5iYTVsr9Vz7+YX5U7ngsPERjZ0oM8Qxm6u3GgzwK/L7AbXClH
FxYKcxYV5ORAvDF5ipxPGYFsoiCSqZqYW8FFb/bNo6w/llZ/4tYpwT8z8gB2hw9G
UZPGjwUnVD1W3XxMaQphRrUsqMt4XK226r65HE2Jd+8aJQJCYUQ2uHvZDa+ndV7R
PYzBeyVJH/tQUbJwjYZfLziC0PNjgDg3G/LkTq48HaU+VLNsv/TiXTaciwwK1gfg
E/YLwvBqirK5Rd6WweQJZW6isUM6xt2tX0QIsc2T/Qs4feyBN9CWc+P71kY/rCjH
j1d/xckcnintBr/u2UvYEcpoSxLEak/o2dL5uZ/jXk4wihxqcRdsVKGChMjqKsvh
Z8A0NZMa4ULh0m4Qyq/7I54Dh4wImYwUI0UwFP4FYQQ34eotEc+WDnZigr22yQCQ
J1/e/J2oSKdeEnQN+/LCv6q+NlToXMpp8sIeV8vXpdeXimBnWgOeMYvUn6UsDTkm
gy60hdcIryxJ6jc7tyYG/SgS+GF46Iz6nLVgisv4xcpwln6/X9FqpZLoJ7SgqB5R
69alAhR3xJXqWpTFUsfGn/KRlr/5qahj7y8Hno3U1GfTiwNw1U8DxAmKgNjFM6rO
qWbQDH4eOYRHJ+9rRYIl7uCsMeORmpyw27p76Q/raCq/kXlEnv8nEE2PnKgL7Ba3
Wqc5ab51VU8zB0NtDDOApH2w5gGaSi9tvBqZhmEOSXZf0h6FDSrHCDqhop/k6dQl
/gO0+SLdat3hYX5GWofTT0GJlVnpZv+oRsfidaXQx8l+4UTvHejl/Qbf9HDuXOy6
CyqvWczYN5LnojEU5KlImgDPN5s1mwKH8S1urCjhg1e9orq8k7MfzZJIu7ftUBko
S4EHxlTAt8BQHtXuYK8GeHgT9QZ+aIpsKEu37JZSWdyNYotVbcn+yVD6+Nlw65En
BoK5Nj+nl2+cIBYe+133t14BEsFXgxD2ujByRXRza0cwuLQvHCU6N2XahD1GCbvV
GC5c3jzGFS2We67TIw7NK+WOXubfL1GFu1JUxHGP5wEstqxxNZ81SPoeW+f65ylu
AIwnVNWC5cyFmGQK2R3rtlgph1I6vitXKlEiK7PXQGXZhKrWpZ8NvrtXQ44GQWzE
y/xGBOC57oUhTVPVu0Yw4g+myjbSglFnA2xlYKpGLa37TuDRdUHLSveVZFDChD6T
ySl53e1d8Bz7It8ZS4iOF1qm7O1TSmLg9q2+QSveqfMpNRsBSgd5lJMdKw335JE7
RGyoGoFTWYoKHgT+ze/zSccDIlQly+5p5XHqqLiIncA+EWK8uP+7FdEJVPKjZDGK
mv9vRnEdFUpix5o23i3X10VjmhPvnMvW/akJXMHIDoQ7kqaoc2U4R1gAMBZLQ5v8
1w15IGb6gXWDC2POvcb4g1gvAIWts6E2YnKqdf1SGyD4EeJjizS8b87w3PYAmz/m
5dLi4YeA22mcovlrPXZ90AxH18PnQ1u1kfPjTW4pQrC2+b0v2mzxg1y40mRc1jSd
QOnKeVsU0oLjUTHqX79z+6g1EDzEHhuJs86vIejalNdjvfdPKzfWSJm3it5rwncR
T4dIXhdwGsbo+fnkHx8mz1SQZsjFeejiFk5QmUBslUligAzcN0I27KyNXYCreTRq
tB9RrR4ErWDEwCrJexk+TLUl/NyItpZFu7WSFxXWSnBlPsJsyNn5cczU2mxkhYEL
Xhv3mqNaW9k/6JLctpHjJaqd4XDi+O69uFmi27SprgQMRCL2Ev4mjifgpq7xGuzT
YNM9oG/0sS85YFmE8V3lmh+Q6yH7orPuhdzbUFhdB4vBwIdVNp+vi9IdENSGsuQ/
DPWzZW6mI8AAlfVPLPIf9eg81L8wfXgJt+fSHJrECeAmnTI6Z4PtbMbD8TofLhBm
IQA0T4TLriCcbnwaXDbsyUA2pZ7kOBIug9W7rEH8JLCOYkILOCSc7nlNdI+OTurY
dNHZ5U4ND2aTH5XU4zAw1sQokuLpfyjcRSbfB/As/nDXBktrQmWGZbHLgiA17MjP
ifWXU1wdmTNaJ7asIWs7iTgLcLN9YLxuIeew3JPOaitfTHDk2YlFB3gn9L7ShCL2
cZngX3NJ0OkaioHfSlLwoL4lQXj+IvaJ8tVsvooPAWCSzdIaLhU8giWrYSUevXvg
IR9UENp4czPwT7WlsyNiK9+E40ibvVGKBXfGZqOEswSw3TGEBbJtW95utrkt6sB3
omc4tfVfF8ufhLD5YRWPzwugHSoowCUqP2zqHe1FCUkqUPjHUVqa6mjtiELOWvGL
Pz7v+z4R6+J0QvU6BwUkBfsSfPqq3yHg6BzoF8vRu4YrdZ4TwBBj5fk36SZ3Rndp
XQEI1rowGkuxqj/1WhdRAkFQtAX3vqlAz9ZDg/XoPzchoSD6R5F57WAUSKJ07Tim
CgwPi/vbvlcVESWxRaaYFC+kyNN3J4cgx/gdV2ksnV89lqfgKjLMUkKULVKexL0q
INWx2JG2cXKYVJgcPFDNmTx1lhHWhJsMessnIuxjX7LJRPrzWvwDp48px5ckqRRw
96p04EpWPKONRwM3TESwFzJwGlofOSsxLw3vyxRZ46VU249u2eCCZcd1DVYcwSLy
h79OanLxeNJVVwvMsarqBX3ugrBvB87SPHlGCktSZxN7qdVnM9dQmSjRYGJiAGuF
Mu9snBqwnBFliI1aTWf7fZesJ1DBVsiTBSieEpyUcujDcGn0AKyXzHMRdVxiJrJW
Q6irr5gHbP3U7tovajG8NUy/NaF6a3sNUilNISV9u0hR7pXVX7/EHYQKQGDAq+mJ
Mu/+r0p9g/UAy3Co5c8IK+XDk76Vj0UJQMeFRROUILaw9gD5P1YQ47FZP0Y1Kw7H
EZLEmEI62ep3yFcUF6dbv+QUOi5WuzqSb3l8iwvKb+YulNLHQ5HIW6+zkvhk3/Ul
SpRpLc2krF+E+egvS2uvvt3twYDD2Xvx8TX771HJC3I+7/4C/g/xFepTZwoWy0BO
mpB+7cFhRWlc/KwBi11Re1llvRt1+uaH6k71x+5zcuCHcn36sLFSLtjv322ihFRI
Xnvj3nLM3qOp9C1A7JGP2hWIkNkULghukXvkd2KowQutx/xghcISN7KcCeQtoymu
pOdevNKLNvZs+CNXItwrtDe32D0VRYaCg1EdV9qY0ayEkhAkQEuBdMf+8X9vqKs+
/XgYcYelTa8YgwtpxeujwCITETQcwOsJBul2nvB13FfAMaFEeeoNzau84W0IY3eN
x65HOR/9h6T7r/HInGJ5sWeI3WaiicY5t5LHSWPcMtVHWtf4cTlUWiU6T5Golehk
gMOZgdfjtLZAg/c23yDAem7ZaM4S82n5Tm8AfQQndcFTIqnVpwBbeMhnfVp1ifju
4ymqZ+bXcEdOkz1ODeconIcjTth6ZdKdG3vBijIg+H+9zwVmNnDDMoIeQVP3tbRD
VeqNXLFWYNe69bRF8rmLFXyUBEtg3KLlegMzAAdcIlcZMiuvSJ5laZmvlTLNQz+O
FVTbT2uPkaJeUieVeBVwezJmWhqAqaUqa8DtauXTEnhNJOf1SrP5xhmBv7vJhVTV
I6pSRmJakcHkQSTS4FtHVH3+Xf1fQaiyALgQE7Y5h92MhqyK/WjJuAH1pXKULOzl
KLrY1wZECVhKn6wcjZnyOOv3b4ghSF9n3KNB+LECJr5sMiLkml5DYqPOQybG/7nj
KFnig6WCCoDbpfot1od5pkxMjPYBRCAzuyu1bdv1vPIzIx9ue2LDcwvjuJqNNbj4
rIgwBNB0drygpeFGi8qVf3ch2uPsHuq+W0SyGRj3uTzO1JCGExDJWCVsbvT7lhVz
HXHNdoPNEM5DyBSh231tEET5/t2SfvW6fA9gCEI2O5qKvb1r8VJP0qGYMhpQ2SNL
sbt2Q9WNNmrC8A8lg+f3yp8bbDIan4T0Jrr0NPD6rijopxsS4rSfACyZs45v0EAR
FzBfvi9+2UcxjT/sHPXxEHR0Df7zorBOogiHvZIQNJaIAdHROSCn54o6WRAotekr
XC5BOpWhjJBox/EAn55dAtFiOcoC/jPflKHi2oVDTgMxuo2Ip9om9F58/5+PdWu8
vz3QSc9cScl/SDpifklGtE4QIInTovXLF+OZSbM9FLy6jcOTfExoFlRLdpA4FPdR
EvCsIC2m/VlDnPWuoDvD+ngf3pG/T8iUzjp+YpNI+QOToOuDrVsS6kpDjgkUvnYY
XyKyWVuWUbUE/2Rgse4sC3hD/YOIRJxEIH19lo4cUdRpqGv7FDrFuGhskN76bLuG
smiwAaeIitu/jDpezOjzPaiJtWZp6V050xwWhSp+xn3qgPFKVCjfb+cpUnEoTmb+
QuCL5We535nQpfnT7QAerxSXKKvEAGw9FKdOga+DGA2ph1NnPRfSh9epmWzdVWac
xIpTHIJ2lt2oypU+RPDWBafjetg0YCdaE3BZHdz4yBRnjF+JQ/Xdqh11mtQ1IQUa
RU9TqInCNHNGgIke7kQuPqVV7X015yokRKj6hyu9t8EhdbhdW1+T+YcmapzLOPPW
yXm3U03u7jWTU/yTEbDUzJf4NdMgeJPu28lqqzgwpRdyMragK5wiZwUHzG35ICV0
DlgeFdibGSNey3Ai77bIoYPXFksp9FV4e7bodXTPIBQ5TaoH5TLzHNPy/YMLeYDI
7xBKzUHtJvcLuKoAL9oNmryvrEH837bhzJ+gC6AYlz9aEf9tAW1pbCQXJhWOfWR7
RJCVuKneXLkAEqW8InSOIS+bSj29ywpIyvaaHvBZaA1VPsIKVv4koN6M62aq/zmY
tstgHUc9NmWxgPBO5pdvO/2edUPfhbzsXK/5uEnEOn68zGU0vMzIW4jmWeMYR+Og
SJ8se4jZtP3q5mV+HxrMlspSxvhdGVrzACK7MizmQOnxg0p9hl5J1ss8wY80fUVa
KhcIWdMqS5WIsQ6Vx9aa4lOlrmJSv4a9LRCAsih4iw15PeqVQfsd0aV5hMJl2cnl
bXr97KnvIe/Y+FWvkyePBJQtQV11Ba8mRs0IgbNzv+6hmetutndwQHxYHCB3CLd+
FGhS8l/ER6lU+wpg6A67GSkDAM4+aiDs6DZCXQuOUrp8LMpXYkRHVigqakOO9aVh
A/Ks2XC+wg2tAl5lojTO38GHEygAgpddnCRYTus01Amqv3c0yozd2uNJIC3/aWRD
UcT88h/Rz2wPjt0P/Yojtcua7KswGA/TaX9wWVjR3bAw1wzzOlDvEG+O2wkdP/Om
cvVpGb29BBvhjPUNMJsudFBUgPl12sn2KKQnxcMSo+xxnHHsrXpIradUjtC23yd+
vFrx4l2RKyUn0gtNfVHRHQC6M7IdxVEWiT0o5/gF0F+vf225jHgW/dcaUjmxMAU+
N4ei95nA1RarIbppz3uwH2V3lz3iH0r3Q67LHCgtXmTsUP+qLmlq8yBIQhkw7GlA
RzSQXPGdUpi1XkAAtNfzFrS+uazQpmEOaAWH0LyMmxTpoy5iScIABi2oWb9pieme
GRozRzu5bWC4UVtqwrOnLZepHXl1fi0/eM6miizegxvzAQmvaAvRKMOKCCCMk1zP
Kxladk/W0zZyriOcifz67YxRwhb0YBuAy5oDU+L4+V5ZAKN958tbwGYcfbSVgEiv
NTdJ3xVvdGKhr8igFae/bf/xU25ZnL8upRPEPtNY2gdLktrfr8DrlsEYHFvPiLji
pwkiGTUimNO7xUrXkltPu9YUV4vtOlVaZtJaUm1G3QuQ/wtPK8hDetEQYw7Epujx
pGRMhX5jDx3p2DQu5dKQlLBxN2XK9Hjhro/CLoyC59A8v1/b7NXzN8UrSCsTrzie
bR4O5fFRt5CHGrhm5WA/UH3ML5W/iJUuEvxCJvVbrSIomQtIFjcWdA58uYlJSqn/
jcfUPExTdLwO4e3glzYJqzSj86Im/Rfti77urybvfwcQKUJta4zKaVyplLZszgWZ
wXHiml229k7DXkwP2gaKIOHCHZk7+rSsHGUyFs77a5DkQD/Na067+YcDfCguj9ED
5fFT4N/A3u80E1siqKJ/QYmVUUaBy5ex825yLV4OB3WyPx6PKOfx9CraNIE4BQPq
RxrT+2ioKojbWes7xstBz5evJhSbZ+rJzbBlyb2PjtnYQBTp7y2kouQqKEPZB5fl
gonz503Xng+p4rCrTxNjeFMMh0QnLwrQsC93h0Ow4DTdB/RpBMJjUOejpTWCgLS5
0Aq3/H608HD87V59K0+KJfYRIekfd4lOY8HWyuZJS8wpe2EQZOtDhG27ElN7TbEG
FA+6KmO0UcYT/mPapHTqsqFHYnHy4xtfpQGbNkzaKSfRnCrkWOgA1txnRZXuAMff
Jl0W0OKQslS+sHu6Q5xTSicluAEBas5H6OqhdtrhM35+h8jP5G2yWfBqD3qpGVgj
36knb4XAZ62N4E9N7NUZolUGY7UmyMb6EhOHQmgxlbmFOeSuMac+qxfJ+d61PqGN
T7/t69/CKGuE6CeYEZmQIpyRkYXu0FaoNOHOl072FpFx1VTJ8i7Vr7CS5rLIaauJ
pHS1tzM6jzC9lnHuWM2kLEq4v2pvLdolntdn3ZGMHGkvDhe38+++GJB5a7PdU2Ko
CUaDgNAAHZRXUh+RNLoXyvWBR76g79aJMGmAku2+FqVuq9NiQJozP4B5c/IwPG4W
+t6TbdxbNWcSFUfFQ9WRUGx9MiQUp3rfvSi30vz724AdjLzt8O7kSd+UyZQ1L6Fk
58qDEh9KD4eDGsxKhcU5bD5Aa5o/CMDgp1JWlCA9NpjY2YfTO++wuxAwSCbc7Tzf
cjInMZXd9yGy3z1yW8u1soFqWCtJu7nOmTlge4NPX86lOsH4sm5ELO9idoFY/x5Z
AzEPwwYu7lXwg+2tdk0NJnixPdyV5sWd62fT0/8vW0AbLJSSRbhfv9h4NvxeM9wD
FW+CYgvkC/zxpy5qRDi6GcyzKZAnOeXm4DdUUCTDBa/xhvtz70ZvgiINBr0w4JBm
Sfgdn1QANiDTQJqJtKbTAJLDte5j8xgWGyWCVD1y2HE5Bqx65BQJ19Cx++Trl5OL
BlIs0oJUUA6ymOI/QsGttT2qLlQ0jdzvAEU3QoLCDLilfwu7RPKRuhO/ai4dWLNi
YzkYM5gmVk61W87pouXyfgr5CQuFQwlDZyjawFdLO/TK+C+NLcOvx2KgyFyinhIt
IrReyqjJMVF4Bv+uG7Vj9K6yyZY0Z7xIAtRbfZtO1GdVnmQgJSI1jx04SbTnI+sQ
/ie61UJpEfthpmznJmN18+WvMWs+UIGJuFDB9Fh5bj7Wea/F3FYX653EQC8TyIDQ
Q8IZxRE5aMnkkkn1E0m3VA07zZBsK4B8x79FMc6r5J+HZQPJzWS6iI1Ily7TFTbJ
3JqhAmLrzA3qFo8MOHkHZO8vB6KGixyTgrTFOCsWdPqQoPU1rYTR/dKnyTkufKY9
MoTVpqTXuAIT89lkA3bgdaa36lql9lvhFgBv/Z5ENssUY5CVKSOxrC7/vZl3vUjS
rdqumrrdqcnjJcvYDKw12QDq3wWjL9dUb2oGy/r+usJxUfLbCGyDV2vaPSyyExin
Yvlf08wpPt9rMKRbpZPZZXa6d5ldAyROyvBunBT8LL2fPEiwzW+XcEQyu4SPt+pn
2cwM90RJFqUu5O+ZuRlUD+azKusBOG5sIOkldVcJWKpARK8iqxi+VT5WSQPAC+ro
K4RKAY9kZYLZV1PUR+hMlNnVXRLFP4wPo9UkWvv25C0+FtAikd5Z+ZNbbjaKRUf2
TFZqoLSjLJH/DXFWcq9gJ8qBGBgRg8RDIS8M2+U7YAQmwluwiwOoeLMhZHvZfyz8
ZANLGP5BMObqfMrbtZdpopzYq7DyLxRR2VteGN3+ofR70dq173VEqqi51YSeW4QQ
1GZDCVbVrQ4Ru5ZH6rxLuDqth0SQX24sJIlJ/sgmIB+kW4R4VQlHDihAY3ARgt/T
Ip58cVLmey8Ndm49gSSsX9LmV4r9eD1Y7q3ACw80whKxj1tbZ+UPhMXMDLdYvE3l
xsd6okgyrqJ755+W/zEG1n9OOyo7/k5bofD4kfEJ8A7nVIVCOjBcmjc2CsgKZtam
Xolma3EjOzactm47HbwBmrRS9z+5ecQF8NM1YvlRDLa2Noh1d2Ht+LEDJh/3PaYF
p+EZ68vKpRXjN2h8XGFRR33SxjkeQ3RsKGlVmc7/kAwm9AmSFgaMrLhK4jTgoKDU
kN4L7ldwZNWFx6DbsLK0rcaZ07d0noPLuXt5e9u5lQOAES2/5Llx8Pu4I4PlnuGX
VndwaLS/iRJpLRGLnV+1AiFoWFKnS6PKRLWJek43mDO3V+o/T2rtyHxq+jpSDZbc
wTdJs3xtwcFGlU048fIERmby1LQK2s9Fj1XHPibmXJpwdHBq2ZAdOz0oYvUKfqtK
xU3IgUn0Dph48C7CcsnoJ8/0huYzzYVo8MW2cCTlhX+qCG2Qcogvf9cXqoA0NIAL
Lxa6WoQr5OiLcXSRkKcfadPk0zdzY1tUTXcXtjf/cxowKM8GW4RB1tK4s2ck2kxY
QzHPUEl0lLKwtuG2a7uPuM6BA0Up4G8nr5IN4oISTzJ+4fqNC8Ndx9CsHb5N6aZB
eEqMHda1w3YzNHu88vZN7SqETmwFquPXzeCipPPgUzWfLN0RSTOGDy5tVJOQyvKk
G2Y72dZHCIi/CUbyUNSWNvThWPQfX6wGiOgVFiJkbfbCzKok/NzLPUA8thkhT1Vw
P4xYKi12r9ReoDbHJrTnQkhCvqbfq/Qmo+kscOYqlWfYCVO/lFNu0rhKW9LXa9QT
n8+W1VFRyDvVfVTEKZXEZjsKPFcQLoOf15GWgOi7KgZMnQmYusCRxkq/DJAZtGh3
GnKsrQ//FHPVKDnotLf9LoLVrJkaW/amD2Om0WDvyiqM9nanib4GlA60yM6AwqlH
kYxdcCMhm2zUvfRx7K8S326oW7ZOantH83RFnJmtsSx/AMduQCRGvveo8LsnqFON
Q3msybFaCFQ11md2WXjAKm38+Ty2ISsBaLTc0bdx11ZoW6wEXiERS521eNrycmo2
6+96bwnbpTr2KKTTAHr3WQgQGmC1t6G19MnQBwHMfWuc86RUBpE71nsOM/2k7EFB
WvkZg8B8PhfZ1WNJCr5t8gmRKBdIp8C/eBcxT5Scz5FDWZypg3VjAWo1rUwXPPMo
4qvhF9RyWsAMXMp1a2i1og+b7FT48FzOHaRbGdlGdy9bK2ZDCGUnuj7B37Ql6ny8
EsAXAu2Xh3Fy0qf51wjKhLcsCSc26DLGFRE70NKO+v2+N9ARbKDFJApp/l1wrdpy
qQyqy6AgzBnQ5CbdoASV0pECjcYSgiQ3V1hmNfbF6yRVJy5RRGa3+s5kn4bEiIFK
Cylz+/1x+U0ekX7yWNV1V9gmoNqTTqXYhckwFMtK/1Q88fP+va2p8Krm+TOz7EUU
JGPkhgzbSFeel8ecEiaYgmtakAGYWmqaHoKnNxrgv9X7WXE/OjQ5lIHIpr6PWWfC
MpIBW1Z0cPLKPnt0HtMf2kp4OVxPrJ5PYC7bsgl1I7UwpYG2nuH2nhWtxCGFpvbM
iEmR7vIxbcIrEKsDxPqiBR4C2rYnK8wqUmiMBvjhxtPOAL2XuTyeVzpXEEl/sWC4
sGHgHz2XszuPEyt2kuxM2e6lVNWXCxjYx06tsGWxUap5D2SPw+3MD38lw7pjqdcW
ur3tGdyoM27N29S5oJHP9yi3q96CwYzpWW96AHu6zqajZmh7CvwNPAk+hFIVEYLk
MadLaYBYwwkuamhawnWslAtr8jZmv71qdAgusL/2FsiX+HG46Qf+UiEmu7eG0Uvi
E1zAQhOpEQ97bz3yQqXlJXK0aH4bgLQAietpynWvTOBYbdR0P4lAxkK5Mue5K3G5
EwstsU+EoLIo2eib1pOHR+DuxquyWF6kpK/VN28syKq9VrJHLJSADxZgj/YpI38l
n9+dQl+kbYxpMJ2t4sWi2WSWG9Bx8tlXq+RkB48wk67qdj55WM4c3C8w0v4Dq0Qs
zA5B+/ZNUvhCdAdkc62qV7khwVWlm3Cwc7lnwFf77Zqngl90ntj6WY+ihXaQgbP2
5Ic0oe/J1+thd0rEGODbcM/YMI9T07Qeu2dbpCqGyO0yX9po6vfyv/VmWdUUYtbW
KS1tuScRXmdMeNvIt2TsbvOYdcukIWH0lL2egD5yZkFLBa2YwIxjvCpNRCk937sv
EJB6rmVFmFuMakJP+Lu5BtqSMumgrzPq9TongyWTKmqOoMTu0sdjebqSYNfQGnU1
4eV1EXaRJJJgCyLitQJJMkjgj+X0e7wsO9AmdhNPJqQoXxJsppZ4Py5IiLcfENsd
ip57V1cXg+QrN7WrJP2fcEhSDofKpynGwcTxf1xTWTO241Wso3Gr2jllf2pnqhYD
HJfMQ2pmcvcph64jxzgJPHeO/qchuWH1fI/aZZ3Cj1jCKnFwlV01GFzgkfn1f9IM
9A4Gt3o7pJED3aSfA4FtUtCWbPQzllJ6aK0xz5Q1aJ2pm/lqTZwCMCfUpR9eA+FZ
wOzlqgszMJVznl4TMH4HA/NwUi1J/+tiXYMMuH5seOVnj/qXdtEdfA2B75pGTScT
Z0rVQe8ehK4rbw0gv0R+WsLH+uEj4u729UQLvqalJuIWxaAOs05yJu2tEd2R+gDR
d3BpZonKx/wU9DUv2XX9S1Ha320JXPUVorAVckvymWWdl3ztf3mqTeA+k7726Shz
En8M3LdCMaAgLSh6z7x/3Ri1/AKq4rJt0i93nJ1S+OjxM7hK8sAEgNHHPcr6JIM4
sckqdzwpJ8InejELYp2/FAUP3F6+w+z4gYDJoxU0N4GZMwH0sYNmcZpuX77vxJk5
8EsBflzkEPxwXBzlyIdFkWjoztNebdKIJEu2J8DinUF0nM01kYmk+w6GxO+uhF3Q
QxOL8odcDefCmwUK6K38EtmdqS0wdxc8XoOTnthPI8227bcS9lk35zSWDPnspRIH
WNOjz3/g6KuQyyxeeBFc8roPFmys0YAT6tYUQEUK9DMBH0W8BTxWWbzWy+lMfRSj
JUppKZbgrIiCgjlgSJ5g5pvgQ1zZoWz/J1D90yo5xw3X98OOGH3PEtRfch/QNLie
jI5SXyhFowlBMsAeFzsVoX5EXzyIqyvmz2Us7hiyAiabJqmaAr1k+rdesv6vOEBU
bMcBiw0e/sgPLdeWgPgidEOE2KgNqb5bBzzuQNC867ZqwWjV4DRmUncC0I4MV+y8
XLun8UZoumrKgbWbYn7PSAwzbpO0Ucpm06V0KAYgvhqhwhiLEgt8yll7gUk5VN/I
bdVvB8IrpVSS7ileSOaCxXI0ImcHZ6hOMh4FuiKoUl0kFTG1yDQM2BT/t8gXfRtU
qWj6efxk5WGUV2eq8+4eg9d1afKWY/W3sTEV+6F2mZ+3YOFEoY7zYt4NXxSMuc7E
v73lvX3oxinVwG1rXQFrh8NpUxcxMEN6fYhwL3cdlq6KFina1B3LIwMGEouP4zzx
qdHOilhCNoMR+0AmsvLQ+crluPb6iWjmyGFEAfDQFWobEGrk1AAIKtUSbZUyhR3J
lCtE894dewhdauu0TW3Okr54wA9NO0k2v6pwPrW7I9MD69XTXMMmKARnL/gmZjeF
9NTPmlApow6TmXAhwUeHymQe2PpOe5BA8RG3uukXDNB/SCgRBB1dz0G4+CF61i+0
qET8mF8eS+Kux+C55mS1w3cvgTa7IJgDS9orPaNg+jU8tdx/XWxjhWhbPNRBV/vS
aRkKN8kBvLX7ZYq7dLsM8pXEHfuliAV8PturrVE9/kHeo/0lR4yfthMv/amm0OXx
xHPqBsahZtEErX+m0+HT6Q+4o9Cyloeh5zhPbEv6MWl0Vye4djRQipbExQ4jncgR
V9zr6yMe81Uft9/21NYfNxTKwOnhtN8yf0UPpRmeBsx3gd20Wiizx+EOQ7R4LX8s
3iFzJzuR5nSeEeM7s1EtAOwaLWcmA8kI7e6Wdxm4UeGtmHwVEKv3JKXHf4r6wStV
jptx3j8Y0TY8wIW453P72j1xWs6xE91wyc2NGh2C87eU7JrJcdbFaldWH16Hr/fA
FInOiBFFMjeSntR6MGbugVoTj7/Z02NDGDfK62tuWnJUM9rWx519M2TVLSV11dQf
0B0JN2/wCTkfPShvnKhxW1T+NAQ1G5/8jYx5e+pOCD+2M/UN0UbzvXqBemOs9kcK
7GcDgANDAre2Yp/b357l+YAoz79/UijbFfEGlkQBhqX6avI0Ynw3Ju6cjfX0xDlf
8/H787wVn4PeLSr8CIDwSMUywgmp8aAPmKQcHhGD9B2dJc/wLAdrqmLOFExDidCg
Yh6DrYKXGyvr9QSRGTEACCkRbms/CdXoVELm/pIDa/6TLDEGpYF4XSKUGVUxwqV2
GWIl/fVXmH1vHGWMXu7kRSIfn+aZqsFfVwhsULFWXO+VsAhj5v5DYW2kVWk/epQe
Cl8je7raE5d96T7MBf5IDbAErzIoMriWciVwifeYNLsx18IJT42/kQg9XupqfT6o
MomQ+5HMMOB90n81HT7toEUFjr5EWaL/hE1mEtVZC4med0imA8Kqm4RHv36Ogcfe
gZYzWCZltSmxy9jTd8kl6sm2z93+2pXC7f4vDuU96/qdLl6KLW6Xi3PEuQWpC4EQ
c5ye4Zs+MW8aN7W23iq7yLhQwHj7+RWlD9YFgX1NGOW5By9/sT6yB6eTv1mYYk5H
L+uGmmL+ttc+kZxGmywUce4gFYwCwTDAptP9ZAYcUHif8zca6Vsa8AQEQfQnCzB7
846M6ae3J0sOzZSJgwz4Z9rsLKcHJLyr0GZhFNYyrJip7VckMJZWZJrrRL7DO16k
iuU6NpvwbFbO5XvIzKkawqDZmO/Z9f0IEv/CVuDRUiyc2Z0BlSb9R7ya3E8UJoDo
7Er8RmlXsgifbirMkhoWgtS8wk4q7nAYxoPG/JJa4cUiz0NJueti8Fv1DrH7q41n
nYO72S9zzmUAa0p3FfFH8PwFzHhKh6BurPlN53lNIqe6uXSdUkOmBk976dD4kLwi
U+/8949+EbDJ1fIjB2m4vRqDE96prv15Jk9DEiNx0du17wQL1u5TjlcrJsq1/yc+
NFRI2Uot90te/+3MWq9GqZLGAjSS/C/iVnJgnt9WrK2vAqlYYy4nm2BZae2EMBqZ
pvb1Ang3uxTek5BKC3r2+UyUKNyp65oZXaNfI9R0ogpV6YAhe0vzfoJonj9xc8UV
3jLmKdlLwEro7M8xmMWj0d7nHbmju46/cVEr6xfmh2i5T4uZfe/vrphK/680lHQO
GBJ4R1W4m5qUjPct9yYVUh7kXJvmWuSfhCmUTJqsVcvCzJqehJhhjPEGbAGyf6cg
S/LR6VYYjAGrCQJK26SwLUpNdbV2tbwDwJzwyRhB4uMB0dvHon10mO4rwfjVHpmN
h4DJzwpAb+kePVlz0gFRZRjmkVHQx/7+FWlw8gTqHCHeK3stDXDlv4+duaTUAvRT
67dIKYW0iej2RWOpiAltS8dgod3ETbBIkfDXWya9T7XW6fwLMGWz3mRsMnFIKcK1
UB8ws9wTQt6sxYF/mwxCw9Biy2Kz4c5U6JjWdMU24hvGR5bmoACLx62ptcRVGTjt
bUMKXnknEKxG5PAiEz2wR8WD/AJrOSdFLi5iMRwoInFb56MDHZ0ulNeZMG8z1WxY
oST8qs6k2Rs2e3uw6Hvl0mZm+HKmzubiAnPGvGV6le7iDttvkbZ+ChaFPaESaTfS
YRlTqabez7zXlVTKo9DN0be0cKRQVm+DeLkjKwX/GRIWGCqdfM4Tl54iMKDKVLk1
ZY2u/rCYk3HREx8sIuFR2i2dONVGjDwMOUpVvgsW+EqfkLq4n39AK3M6AvO1ua0E
bm8OKgpwPXLFrlNWwZjPOLkMmVF23oi3kqKdA2heqrWwmGzy4qsOYrsuBtTYU04i
QSnMmLGUbVwF9+sSi7Wu7E6UVJ4+whfJVE4SHmdKVs9xKo+uiHXD3Ea9pDzqRtZu
Ri1AwudibO8TKvu2MG7aKj/PukbXdNS+S4d/Wf37T2WLbLThnHt0UpG157ZSrm5Y
fgP+yECSxoBktYcbmmxIYAPdnudzCF95VPv1miWrmE6zbjI2+RwUEkPIZjiQcjMh
eK1S1fBab9+x0aSLTpLdX4eeVZUO0VkgzFJyxFcuo7uNi6mMdxGfY8b7Bxd4QBXp
VLjp6YmpjGESNVNOtFb0QwcyM/VpHWE/ACN6zo9BiKRhFGYPaNG7joP47oWivHkQ
GWOMsPBzvrT9WASgMCG7SovuYe1y7+grQOLSjmFR0w/XKJIvKymI74/RFuNEHvdr
Yb229hx22RXHXzbiOPG4I+9TSaPOpHcUv5Ew2QFEEmy/awK9HZgrQpPABXxj9/Ek
8iGo/Q03wLohfPb1lKyBlrUHH5kY0Fjh01VopO0jJ4R3QD3toRhBC/qvRlqfc+sj
A9T6we6Qg6vbGuwC+n1aOjZGNGNBw0PuaybQeqAlc+bAB3Wk5hJr5owlA88uz/GN
IWNqrRntmZBokMPaU4uX2eFDUinrj/cT4yQaA5ThXYN7mc1i72Ops+lLEEIjAimx
PIJCkivWKv/UOQP8JPTMfgqd0b4rn+AWsjQ6A5jplV20ZddAYv3vDgcValK18Dqe
JpXfZJeC4JqT3wLTwoEdCJ9TVm0ImbxSjzI2hu1FSj+XenOV0EDWzpfyiPRfkqxj
7v8YVEgFKZXVdYUCQqUX28NUQ7ejdxD2rvR0jmm9KXZwn+riTXB1VSgGljj51h+X
3PzHKtaBQJGezyokaqz+0wf7fwflRCf7aiENHCU16tYPzX96WPDk56RcnsLRz+pT
N2J1CEZGifW/jGFO5B8IBspHkg1HxeKXRASEpiCJzceBeeJ6I0pe/6N+3I+r++0O
LwmYFN2ZI/FBIOvJBP6HWHwhYiSDgMHCnqxGHe1ShCs1zfHNM0ZLkeR8n2e+91gB
KUyPIEEHn9GhpEVt93PF+DcD8FpM18OJ7VLb2FVH7hI6D1rlT55xvirQWcWS083j
kblNY1//nQE0O4NuBS7QHUBx5Z3JSHk5PV4SDaqTadQRqaS5Tccwwi4cLCRhTaMQ
+aZZwWN8NvX4CKMxNgQfD53hLXRR+qymOfuKWw8v5n/H6XZXqBwJUhaKkN5RktVK
etveMdKr6a7OKr8gYLFWFKFA78zHWgQOCV5lkxMIDg4kfBNl+Q2LjGFpkgTK0qHH
659KNZG9bCA5x0dMaO40r7/hVjcWk8nREhvf/4WHd/MpvwjVQcjRgL+tzICRWCht
bPm+mK3EHBXjzlMU/4woB4PPJ3rldrVywsbEaC1cwDuxd3q3zOk7K5IrvwZ3O66m
sWdWBirJ9OdPLjvuUB/ytT1y8Es6+uleJJaKA9zIWqsyFI1+HWw2huYvsja5jC1x
TgRvUqJB0aQnEpmZal60wsWqkUU9xk7P7nkCJprZoFPK7Kn7e82Stn+C+AtF31r5
r361uh/6iNckYCxMDWmdz/l8+piyZ9hKHlJcaEc8Txq/buytKi/HrIqUTEFmVPzr
KR3/RqCjvLoXbGgvK/ENRvbpPfBtIwDFANM9iP9NKIEhWJ2NEGROB/T3Suwqeb/x
rduUhQKhQ5whhPfsPiQEq6XYRIe6B1z3DDRvyuXtng48GelcL6FOtqqi6H559p60
9NmtxUHHx4jMTmwCUgHJaAgaHz2yGH624TbI1L94jx84yIwmxd6IGujtGolD3SpU
4dnDLaVGifsT42wWibxFWlwCnPpCyDbEjFp86ef5Jc53J4uAtDlYs1lxtHbLBb9d
h2Vrs3NO2kz5VC156saFC5CkQK2ajOpmyfNLrO0QEp19O3lVKhdcxILDR1j5ziKn
+dfxTdxUKT8F/CQ2PJ69nlQbI9hSwxwCJNiTPG8BT46R7/VavbePfYrRXj2Ef3iF
qBZvEAxiKxNg3l9G85siyHf+wmwavsff9uwDm+uZUz6j7uixlzXUsYIVbjWK8j3D
iWYC/JT2uroLzApksI/1zefF7sts94ZG2Eoe5St4k/kiWnkv6iOA8wGkWZFhH+N/
uOvUP4LGJelSy7eHN2Jra3QlQdYrR1Jv+izM10t9/pWeJmeNCZgaQ05+2+RxW/Op
B5UYMKdHv3EAvhv4jJyaWMFCf+TWVtn85noH66hip+87EuZT2eMWON1bHtOsIpq2
bva/h5NRgTJZoWgJQgLc7jvKEwG/DflgWU+kXO5dqXYNfSkSUUbz+nR9p6ZqWf/w
iSCoYwfcdhbXT2NwdnRpqxwbQOxmy/UhsvBdIrfRjlVclHH2VeNOiHIljo8rbXV2
vnDCzY483tzz2ggxBbDAjoKYY2gcr87CIbfFf+tGDBcPa8XltljPCOsJ49zppztS
L/D4fKi6D6Vl4i/yI8ehDWa/CJ2IXdh8zH7yKarOA3FuoL9ERa+QyugsTRqJveIO
K6vOMBP7L+jH1Y86NjdT4DAKDYTHG/4vvJP5mforF9e/Q5jGq9ISbnsw6Hv1LZLH
gW/ir0a/BCchOpVph+jW0U7+YjGGj7kyvyrO+TZwnhQsxBU2M/cvqKHU/hqE8o1B
6qLruw2S0Wrk26Jt0NqgEqMFrNiwU56mpBZbNl0R8UK8NvvHhs1IQBXQFD5e69B5
rEx86CQb7J1u4ovUHS/pNqOJVFRdzgf/Yl0lIgkglhryNt77KK20+eiiQwHqTda7
QBqesiWTUDur097mGCnMMG9avDlfBM0dUVZV8z75TkunEgPDer51Mv1N/ALRUiNm
xgiXCDqBKcRuMbC3zxT4+0K3x/QSCV4iISvQ2oAdF2qq15u/tU6ui3GvjxhE9h0C
o9jsEn3L86kYaOkYvdiDf3oaPum8Run90GTuJXpkwRZozUge2V8Z20P6NWtkls0x
taxlx8+3PaMWKV5dW6vukEboXk8Jd20o859GdZNlIJB7V8xkZD1ervxosObnTbS9
TQywCfLt9vhhPDh+AB4Ya9uOgrwiVgnJEfqhqrqxgb4j0Hg74TRmTe6oXDP1xYFv
nfhqGR8VAjwiB7FNspS9uVVMQsbhrq/pvQFbcp2Noe21iylN2I37Tw034qi63uBX
CMe8JmuKKDt/7mWbhfKENzRiJx00ZGMrdj68xmPGepxA5NP8IYigFbURB98aSZNs
ZHHF3SUOH0BgxnxGJXgS5+04zqzyu5Xa7WcR5O+5MZgHBkKeRgD53YE9I3vJXRUA
7wOk5ZkliM/kiy+hUDUJv7zFFAo5U1epaVOoi+EMF/dbHBXR+Ycsns91XaCrhgEn
BjMHydrIW+uv7pJMqqYCMRJ0AVzBcDPWq/iYh7Zc32Wz51l/igb6GgE1cbphBBT/
lavXveM4NKajnuWMou004C7iJFOaUBZXi62CnoHIp9giMhy5s1mCyxS3HDRSgMv+
cjrzlCeId7tEn1hjOKvFov9d8oKmbcVRFgX4XmibU6wqyIdo+G26FzzktNXa6Tej
kqD9LRUSV61gq6fpDERiM0enWYcm6wjjK+CJDiSjdXx8rCvdUZrjfgTdu1p4ejuS
PcpinjPE4Nn85X4voG79tax9r1jsT6x8QUGCNPyiC3Sf324PWEaiZTDtWyJB01Nu
MGxqkEckpczKZTZQDUHgsltNYE/vwCypvOvaeg1tSsfapxSRK8HOtbCmORXqDl9x
+CY4jG8SbFcvHF4C16+m184wBEgELPJO97NlKN6lUSX2+0ECevaNLKoFdPJOiXyV
Z84fqBOpoLOOcVpoL6AXMhQORWcbAO/khybncflrv5MrJDisr+MLRp1M9V2w67We
STwJlvCOID9baYY8b6mID4e9Vh/12Fpkr6h7WDtRpClXHrTAk0qTR0wTHuCHqPO8
A9Zuhai7twQHbwhmsnjqTxmDpZiuxaSoGVJJacsKFNUvflRZzc7C9PmM5iUqD5dD
AWHKWyX+MIujDqzygnekpiWgLRF6sxjN6RC8bZFsxqJmz3s/Bl7UAfsMqEnmydfq
15VMbg9BsyorsRCXa/FPkgUp2YVkbLz/0zR7o3XR7z7RZDzkBDdsmCdr7U5r6Xxc
oTm0mJQSiidx9uztfHBGuFLuWK8Xx9I8pXx5660/79dzbnmx7uG0MPDZOxHuDQ5k
SODWa0HTvncX1yds0Q0Li4bZcwSkH94ym9Y1cTUri4ntZBMPMDaD91JS6xO3Cnsm
3yJWP7Urlo2DuFeoDsrNCkBE57XmkgsJsSAF05HXiv7LaeQeToy//3HJddk/BQY6
3t7g/YCpc0bM0kXuTnBSS6LWcNte052/+8GiM2VpkBUZo5N+sCMX4z9zwQ7ECQSP
Wy1BeB9yJCdxWaeUZqCQdL/Pd26TkJt/qgY84B8eqxJgIHr0PU9GylGbSehfQ7ni
FjcYEJmCXJ3Dx7qsF0khKVuxUaQvx9y7W6kHnRwlm0TRTQjlq+CDY3MjsRNmOig9
hOBxExPSfexIwvM1xQGaRM0nwoigZLxfhf+Mem27HwhEc1nPLqgmEGlCGBCcjsk3
1hRuIPXzb4YOvlYVbIlfBXqkLSTDw0OKSIEYNv8S8w0GYLJSAsc3gXUTFHLCO62U
LcWc56l5+a64b3uebzHl+WX3qZKHJOtDY7amkbDKUzV7FTQa4I+mE3z2iER6tp5Y
i8SE3tP68Bsa5Z5l7hfK0qS1M3CLQ2A9u0EOFTnMhghjWRQ+8taAnRfMz3auT0lN
/ef6LZg/EbWKTGuTYJFA13MguEn3TxBREihFdrzazkqLDsF0HU0iNv0KkeHw6ih6
stVTXbtmkOyfoclkl1AiwpOnylYc6ZMmkClsQtGtmreuhhV7kWTGdJ/OxpeWriYa
aBWEjWKlbjERRr/14WsPxwDSpMFBHQU9lVfN6Z66kxgMQmrnYoBGjmSHU+fhzz85
XlixZlyDM9IPMeiYGwJTxQhT2nuUc9kGVJ/mRiFCDAi7KB6iJdjVVWEYoRjYxGt3
ZpyrUtMt+Mz6X81ILEP1FoWE3IzCr/FWqvgsK5xWaZqzwLEezEJLtXU97VToICxh
KJ/kltgtkPg9bKvWNJGWeiqnYyooDVmSV65/My2b+lREXlT3qLXpfc/xnB6D0O26
PvlVwgIDDNOvZJGOpvX3yJh1Q2qKSJBSFKnNMnRvzLjWO3p2yD8sSHaZgAIuuPzf
jhbju9hyO/jKHOgSBiBkUQbFJrcsCjC+7DfcHFkrR85ra7PxqtiWiPaTjzEuNZht
w7K9UGwFDvq98S4bVw0ZOeOp4shFJhSZsoLPRlNsGUFEd6GWNVhalNKBMVP8Lv6O
VReatGCno8NlE7a/oDeB3cSlq0CalgyvU35BqbAyS4d5TJkmAlgnu/g/AySQk4xe
8cWqn0+QvajTvbtxOjLBWnpYbYvUHDtXOPOmbbeB8IRi/zHKnGALdGErM2bdLvFL
Qi/Kir1frNKfn0wDxFdqDzeLhKzhB457HoC0vDeohkHDXufgdDdSq7YDMDN3C//P
+3yAfx4pGsNHVJtUIbKlFHpyv610BwwdtdAuPQYoR3+lMA12Lv6DkGpL32warXMI
cYa7T93IrvySr0NDcVEU46R8YZVOKeXJDBMeH0A5tkPwXEjnew7g+92a0Xt670gZ
Dwl9fCGvbhJl9K/KZkAadUcYoBZ3qWF0APbDuAX4GjXx2QSm3HdN43B5SB2DMSwj
9+wvU148ieGkVlEgQeof+iODF/DxeL9cKckLIk+qFIz+Vpa7/QWG6sLlhEqBHyAl
M3WclHrblu7qC3Zrou98BOZDF3ohIoaFTFamHbNY1NgSpmsdO87ChZQvqtgXC5PH
0JTtbHeWkHTa3P3adgOymTeFTcYnLTRQJfpHigf7Hsj78jwaoyGjm8gPFMjk9u0H
9mc1iic6rSRI97UTiTLV02dworiI2PGOd8WKL10SLYPOt4MEiadOb69feM5FLxop
2ZQjZa1jjyFO4eZkxGWQ+Sy/8nqY1ua9d6xqWyFdylZuS8Lhv9RGOwUeHiovxq+D
QNkuC1hw3fP69lV7iBifncBoAehotqMQ7BG7Nr9HKuP4Gp/MkMMTnQyYIrk04qvh
Rl9hgYGgXboMBkFo60s0e83lsRlW3NvwTmjBhf5tf3BzMM5LVB7nYV8ghKp4yORV
LsLluA6ixIU5+4rmUoTYhEfLr4SC0HsC7M+541u11bWNM7r746Qq0KRy9X/OcnWm
SPZsuP0g+Vh3PJL02+2nR+Sb9ILPk8ItSxCqNL0uqavWCV4qndS/pZFmc1GwCgXU
nVgj9xZWsutIqndwLqLaaylnRdamQyvRBkgssa4gT/1EqVsiClNQUc4mCT2I/L/u
PwYi8QqK5LhRvtXOHTVztEAHw2G1VCYXdwz6hNmSeV/1RoKMRJSon6fJcU/5aDTQ
kj4cacwLh0WlBxCN04/d8FbNEFfPyPGFCyu0CX9bXjnHGhhyuzNr+aBWrTGvxTYG
HfvmCP9edYA41b/JnNuXCrACJUK4e8EDWwgMA8wffuDLZBFQLBbBGTAck89yyk4H
i7E2O/JRrLBbwzTRN0EZcv0j17hYGuYBy6hf/GtRvcRJtztxB83Y/zjBbovzbktc
QZWSmkygTJwP/RHtZgK4p5UKxkVsGvuvxBVmvcQ3PYPxjVzwHh9IIv+Y8zTKaU0m
T5EKElwjCRk098ARz67EwqlR8UTDI7fk/LBNwxVEixsgPsgn9xGXSjR0VSpHgXzA
0bjIszCduc+RGsQho6lfED1ydJMl/8zyHFvGakUchhEcEf4UQ1X9klwMicERrSLY
zEWJpYyW4YQ8+/+gOVixf27J4p9Z/M1GBV+W6ueanNEpZUzx+SFiQY/zUDe/EgTi
LjApghRZiPo8boT5QnK/66j037ZbsDarMgvULfOYF5ORseeWaxGEDO2T2ocA+Gu3
gyusZNzeGEUnPrBElhMXxK4dU++oiTvU1tVFWtzEI7hUPsJZ5Ulibkhl1TC3OsXw
AIbOa1ERyS87oXKt6rNuUy/SerY/WnrUByfAImhHN23tGak8nJEmG7XsZtQm5mGK
s5fADknwf2Zw1pYJRfyxiJaitwNzIxDIrMocHFh925b6M9wHH8Uu/Izx6fZZnjcn
64wHveq5zVWrdzxHzHToukNiGr4EaD5/fLnT5ZAv5Gm+e1vZ3p2nBTeewkgrfiR+
U+3MfsXHOWC10q6XA+DCIV6ODTWqwdamINn1uQNiM5prgQB+QISioABv8PdKC4Jb
jksgb/gsGyVMBCXuqPExj7VXWdq7f1TRiLaie+qpjQYoOdcE4FB9tcZPbspzbLnD
7sHSW0kTNWutwBc6I7gwppnaGLYdp+M9v3VkNY5kEKlr6jxzJOXh78xHxGtc2P4W
FyyslIcwoMlFbB+OZpysP4b8nod4p5YB3zPzCTcimP73bGPdvv/aq62iKjF6xzx3
98c8Cc+oLVnNwn7dg6adsQMVqPg7Ut/G6rHLoa5Y3o2hn8bFvhhSUuxNeZS9yQ4V
H6VqzOvWt15veJrGZMPl3sQW0LeYLoZ8kgUlFd5LUkqemGMXRsEs2h0yTbOWIHqS
v+J5G5lF8m72/gYcXhD1sIC0/vGcFSq2pQGQYfKMxTn4jpN0SURkesWXLsAxwscR
u5ApXHDtZPVunF8RJ5oDnsydZ6rdaR8SKfwQShEFC5a4LzU79FR99UDOp+oOSogw
xglZDy+h3rJnIok5S40B9NdCsolLLDBDEu1zBtjFkguxx/mAE1BNPgtc96VGd4II
cxc9jNcg28G1/LjXTP+vIu9EKU3/APY+fbGcf0I6dkeiHXM4gf0oCqZygpoNqppb
vbiDyhjSt9i1W6CaCrD+VEXZfrqrCXTTdUmtXFpaSEs+KlsGNIZxDm7CrxtAbhjH
D2eb5GiPkrW17/zii6edZp/p8dD1xxOJ+72hyU0MKnz4bz76krJruv1CxZ9BE/7L
8YcfPuuW6wCyiLgPUQBEbETWhkFCJyUaUAe6Iiczccw+HCkL+MzYeEwe4OCuTNi/
o43Vk2oqLqFm84C7K3UIiKuB0gl41xWfn039Mve5UDuqdDw2mafVvZMaK3ZcpXoI
BatR3HszzSbMv7IonymxtpozWInmS6UweXZpIHNJwG34JZO/+Ox15CApKr41Yo6j
ot2TuZb/yCjfzsHf2Vt2eyqbSU0K8AkjJhom0UMdXt8Py0RzZcdNuKaoQRklSh1B
Hh1SyOB+hXFOsqDU8MqDqLfc1Ix0OnzA03N61gVJsp84K8KGn8KbceVkEkWuMSb0
iWciVwMTsGUI2qhsKGGYal1Em/vbORAFmeyetEv2acjmiX+BO+RMmreM+qs7C5rj
OPTDnStIJdK1WoSXiZBu4sWqlzef4+Pu8uotdPAy8PCarJmRBpgxkVwN8bcsQBnI
KV+PiBPdlyWEwj9Gj/nj9sYBJOPzU9XFBnT4gOdu6lbvW56jk/QRdQ4Hd3koVtDA
7GRyeRkEhmkRFdy3ukfDpeIPjmOOpc7OJm0yADnEzXhTwAVr+JD1pi8eyhsGbzh3
TiWCt8th48PUO8jEpoKqT0xRq/DPovcOeN/T4ropvcIU2gmsogX8DnFViT7Cro7m
JUGRd6a6H+CCozPvcHBU4PuWCwqJpSmA7KfySL2AxLWaPWCHC//hdBHNsLUHi5cM
f0n9UJkeaVH4okJzToCMO0djbojniGKYroIKI+AU87x+N6sOeBo2mv/rnOdU+mHV
2agSupEi2YF0FJ1/D9YoB1Uh82VHNOpGBi/dc7k9GDnp9stNmwK9/M4lOOE9pD8F
c9eG/zkJ/J+v0AIAfNNoUAbgtUklyq71ex8vGPZRtEGj6+Oew+WLKM9SiQyZmGE/
PD6PRWp6btRH00oManAEakaNHsgBr+WrTwLXTFwNyuU0qotKLWfuF7S6tDgncq1X
4phTbmgeSO9XvG62IoWusjlNSNlgPrQKPg/nwJcE61LHH4lxPO0QNog2vYBrO6b1
KgMFzA3dYGxEoboXwMryBlyhRtEeLCeDwaxwDMk9QUdTVT0gbvUhTnzMxF2nMHln
cQyeyX4dZfrJVPT0xGN0sW2Q2DOWJ9NENGu/Xik3R4Gw5Pa9khQ2O9RTmjEPn62t
UhUfWn2wdJ4xmGBLTwdr8UQ3IKaemjuUZdHIrnTqg2K6WvUI/3M0cCVYbhRkGRQ5
RCtcNLnVwUT8cXtRSB22uwq0VYF7bUwsFb1t/cRNcrU+l5Dw2z5AHH5Oz13+3hUz
paB3zevlwa6tEuUVQhzp4n+PpFLZshZfQ/2WljGc8C4QORiIdYIHAWFrrBDiT9nc
lUwAwY2Y8lUlgyA8ISmBUUicJAOnabBQJ/ahcSOzb/0e7R1ojqHTSBrmRyyeocdj
B+hRijUEEh4IuRT1eXSqg4J464O6dfOorTyZfTR7CQdahvnFyj9hCO8uptetqqFh
Xvr7gHfsWSOVJ/r4sQpiKa8e+QFV8p7pRCAu3UIjeAgXMxMDAz4HFdC6/RzFeWHy
eTGqs8upmEsI+soGKcp2s7uLCbwb8cpjhWtmlT0pCMv+44Zd5KT/+1mHS7jBAnNb
7v2iHxnyID0odgQQApzULibOyj00eNHNZQC+SVIAiKnCp9+NGnSmIET/6ucqNwBi
Br48oFINTFaJ1ORCXnalFBGE11Yse/Vqxv2QMx9aFYEppQFCkZ31vtU0/jvpUd2X
gpMIjVU7cBx5nG7qoXkLHyXE2OQmHnxVBdut+97cYvxX35VXOL9wxvk++pXkyysj
98iCtkDRHdGuCwEN2xGoyFKmAlbo/W/P9ADWLXoruoNnwFcawq404g5OCgFKLt7U
OFfjG+WcrTeEQUuK86FX2mqOp8mwsr5bjrv9bLx++MorX/jiNo6TLt/gz/wHCj3/
j4KbDDY5C0fQHoEpv67VRbzGms2BTwOla1ImNCANJVDunu6Tdjnet2eEWS0MfYDs
9TqHWk7koZKjVx8m401ViIMfRgRLGJVrhna6d+KWWsk35Kodtm1Wn8ehpUQmcC1p
Q3hpbyU7gqGWuRqOUAqclPcWybBXR7hqKc05JVfh6um0VzG4aZSsKko0RFE3sbpV
EVXXrju2WJ0rUMMq2OtWkrzbbv42reRgb4jTKA7QlilNfZuDTZQu6vzwReNURzj5
QPkmWnWzGUi9ExHvcucDEy8r26m1nMBabnqr3MEwDf7E9xAzvcguCIzx3wNgm2Kj
M/kjszNjRcU3lHlglHKtSXSZcaEQQuRo10bIPeyUTiUb4hNVcIq04AqCBokx0Ur1
h9Kqyaib/2bUN2Fe7qb+R3w6nMrmbSfTYsHNMgEfeZxCZOBxtttJwLK8eO9MGLub
IFmMxHAlCmxfe+sXa9JQvjQeuWARGGQM9Qd66CfkmkJYDZK3W+rZr/FXBPzk142Y
017EEcGpbTFoQMQbgbebC74HjpkUwlHmD5gbyEst4YTMbnD/jex0HcK2OO4GgnoV
PGk0GY6yEhnLRCBrw7DBPV6fxdLKaDfUpgV+Wx9luAXfoKdmkCFlg9H0H7bfnFlm
Qo3KJG3jEdmtktCZ/PVwh1XrP3pEeXIu1PtcCnQ7S9VQEVZ5CIAvEdhdvu3uJrpT
gpLc2IJ1qU96VdZQqFhjbvfHqEOuN5um+C3raWhfMMg5IqKPxEt6aj0BTs8NrnY4
m2cqBTOw5dfl5+3AiRAnGqAjqA/vjvTBLKICMtgH62/XJ7dK7/Cq8yNZU0ZQmDuJ
8YCrC4kgKT2xekGvjhlh1LmMaFM+ualEoWxZyV2AZPfLt1Scc2LVz4GUHVe2wmcs
bhandLbmDBKBS2Es0FA2ATUnFgg/CCxNEUrFy72mYc3J0lwzwJGrZ0yRzS+DgC16
O4M6C2cwmFm38JGp8gAukJkSbo0II7KiOoukk4g+s4wcdeahaEzL8Kb1uDpPj9KB
Qji7eEZH1qUY2fDSCyHpPGrsfLsjFUKCsoIg9WXXvEDlshr1Pwu9egsG0EWkw6mZ
HeE3z/hHqz+NTOoSBacmYlHuHTGf0df5FqeGip5SRRoS1lJE6h1AxEE2S06ydgWM
i6lW+y6C7A05dUCInGUBZ88R8bgHvUUmCqyuFm9NLKFnMHQkewS91yym7yYKMmu6
DukHGDZAofxxeQGzSw3zx5voKmX7YG6gIMJH3aL4+s/eCdXe1WGuLqe26vHMYUaA
dzjSX1hlVlX2Ytj+nopogoaE9jZdJb5TscGj6jSpErHcV1DnRZkGUtFLbOXX98Zy
wqKrk/we4qHG/5zCTY0BQMJNwBUd+SKtThn0WMQCTNSUiEKDxwgMmHS/B8M+/VtW
vazM913KLy1kRGbPhWKnzgXUtUJcD/SWxZRWLqRqPlxrOWXE8t48GAk4roOiCOm8
YlZwnxdAZVvXL4GnK8cP4mrAjpRjCEFRk+xWbPM+QQ4YN4bJP4t5oj61N0BexnDD
zsGP4UUeg2iGaXvz/vA7VZ2gbBK5PPOL9P/gj7W9Kw4Z4yuxJoXDQnk7QJuAzC1h
FP2LRnS/xys7KKMdOGvqBZo5HJ46wMXV4T9iFDaEa1W+8eHyIrjOU8dG5sYJUblN
vIWXArKdayAkjOz+X4hh5ZXHv+Yfeay97dUTXtrJVMOSIgHCfaF3tK0sIXfuwNJI
M4+dAEjQO5fnmYzZ6Vog57/p969LlWxBajvHMS7IMiCDiLJ7a8fIEqWx/XrqN1h6
6QnytMRc3q8lUYtezTz73rcr8w028DYRHtNL3AscEGEQfstNDpibT7wNq0M5lReF
ER/0HReCJZ5lzCQZAT6kElaAwG6xf/7UjDZTHWRNn6zi837eEP1ObHgWu+cyDE9n
YbVY2oNZcqnkNH1iQie3VdyHIi9dT6XPTm0OTKR5xHJTQt8lClJI2e9rTqOlAiN8
0GylPrHKPj+9W8FXjdRAFELEgDry65sXdkiF5f9ZEDWunClY+4FM4hyBSYt+uX8a
sGaSEaz4qK57GkBAUmPq1RFf+wxsVgGxOTJGqqfnpGY+nLf4hjzD1UyfyWatTCnE
4UNrYnl2VanKmaN13qbdTfHT3397Xv2uXeV7j2/gbNeiogAx6P+yRafJd59tfai4
6VS2QFPHFtNwRRNqoYOEnqI0TUjPccdeqnv2BpMkpkKM2vakMu2XmyiMyaQpTn0y
//ixSMlJCmi9X4InYwlbWPY6f/X82YXJV6jkoI92mC5Hsh4LVE46jzT4/MJ3/QTY
2Uh6p04Ew+1B+Jdv2PTYmXeJaI4oadzgtuGQM7uakhKVmKvpnkC5SFLKnnXXcGv9
5HfZAWtgz607lQIiCoEaPUCQA3mQWIb1YPSZJPrFBdENvR0+JtcL4G9XwQ27YT1B
y/RXa0o/6deqF1MUhdk5Tdo+AdmKCbUI5pmV+AC2rsOZCjHZK/06c36QWhmySJS1
fvG6UvbTbozsSiV9IIUf8eaRfymoBHo97szQ5zG3a6H2jPF+N/G7DKijp1XdAhWy
6qY7EEgYbAt1NIB8y5kQSqmTJrsYK0wSJpUleUs4W/iKd0yqEpZZVEle2qk/w/be
hxRmwjMyaJem9uqlAkYh4vjDD85Jn2pdRCra9QDW6hpag76lB9yD6fL8k3bj24qt
Px3o11LlIWiOzB4rw0YCck2wZ1O9qtd5lbInDW8NYGF6FerZHyRd6h+9pWuYJVlG
49YTEtl6T5SOGlEmykTPlZ6aqddb+1T90PjM+rhVi0FRUYjAXGn4RYGHJ0x89NkN
wnm637oZIfU+4+xra8zDBfHT998kGJW9i9MdWmcfi0Yrpkju+XPnKKaFjbsq6kqb
DvZAyQhnDXklSL2kn+xzYrBF6ylJ6Onq4BvKGedaWQ6FTFYzYHJVY8yg5B3xGO7v
G2rvFhXC4SXQPcQfhS30rPcZEqP3uLH5sKxxOiu5jMp1T9Ejq9kFjpUHI6G91OLx
8ZYusNNVTnImPRBZOUyrNVaDE/a5fBuENu4KPFj+n0Eb2+VNw0tX0pbbFMUbeVxt
ryhL8/eYJk0uzIbDPLOe9u7QOPV+IcQjv5vjhuYoENZxrBn+DQfAzH3HF/HVEE6C
ogXWyLZ+eqVFZyffrW+bnwC5hRsIWdAuyjUYSABRo1d+Fyd39wjU5l5Hqhhc7OEB
5QqvBwUeNzIeCSyvzyyRckCMg53sLYYANAomq4NcNkya15AiceKxiTYuLfAukuJ6
njsLMtgO+fcvWkTb3Xd6D0ku2saga541p7F5MDx5Yg8dlCdOFPMEk2WQ9mZ7ZOva
xTGu1uVSDcYekxuPH6VxC1bPvtmrWVXC0nruknbcmZsYT2Fw7NZ+6baI7w02JY2Z
Ag9CeaHKe3xkUEVq1OjQP+iixVmkDsa4D4PI1G9pHqq4BrfALwo9Yi/xC2vbcVl2
b7+ET0GJr7QUTF/tc0AoQGiKnCcSfPdA6NSZBOlEDsPGTx6w3iYSq2NaDSAoMVDn
ZSbJ85ViDRBFj+4F+wJaNdK3Cjx3kGDaJxlPhCXLlQnhG5o0fiMb1tpeLjAqYncf
UkuU18UvpX/nPJ5PBXQutDrdCAhM7UHsb2xaDe/GZc1jhcT+9ZXYLftS+GAC2ivl
7Rsud8OFLGjuxzjhyk1SZZN6/+1b2n6StKIs0F3lBUtpyWKbRiC3iFRQ67q+e4jS
mBhQt7kkih3NZh6AjYOHYBmNtfySItKcJL57WcZfqcYEHGoTRAhhkeWQC+Ybkq41
efxDkej3VFGZtuAHgw9eyDYxtU0l2Wn0VIFd/eXRcdGRLU48F67NwD6a2FJHKKb7
iwYof1mrtSTwMnZVxogy5a1FMa+jsPc60IYP/pANP5qQlG4xhDlfX/Tl3jVfEWFN
4s9lrzZuYYL7XVEj5/jyAu4vmDlIhzbECV7bSxIdw/zueoYnlsaR2oGEXoDLbXCc
fZbuCPtevKanuKhUhJl78wFCG0NoaBTJ8FoXWJmgDsucUn91zyjy0rofkQtmasYm
KEP30XQGEFBK6ZRmlZQnYrUQB6baQv6SrTYlm1jIDZBMI8U+aD+U1QwjFBIN3YNJ
oS3FesyZ+sQ5pniUCyURdjFQccMLo0U+J8YlawfgvlvC7YEObJfUcuIavA2akxHh
BLyf+SoYOMwtcyQLaA8wyGaLsOtXrRrNKVYEvJC0wIuY0k38dZd/022k0M6D6Lre
+zo4mzw88qpnqVqUDtdxLwr1phzCmX2bKXfYZ+VYLM/IVEgmz8tA8NYLIboCXm20
qQssCtnFfAzKbEDjkJQEDRBnO8IUPo4U+VaYD6/Mc7s3EnQTPSY3+ewfwWwlMpe1
wdm9vr/zVnnPWSUxIpxL8ysUGFsiADJgCt2NNqP67wER4JjtCsScQ5Ekfi6Nqdkm
N69hb65JePDlqOIhHmjjYU4oItkM5iDkNh2D+2aqXpqpBpe4VDkS6P4q5jw60CCT
oVulVFOsn1UDZj7AjvoFmbXOfdCgpeKmEtT3iSm7PPy++WpJG1avacTaKf31tuRF
jWfgdPsG3U69PiUm0mbEiTXwF6PFma9NXISetkvCS4GZZrSyydoY1oOYNa+uTq6y
ePRllfTUnJco4kOaxez+dvV1HOLP8ywBtgbqX7gxm+wHV3WZSOYxRNQNUMEkNyC3
zgIt0LguJyvZ/3NtL0/2NnENc6Yoltiiqu8gddRe4MP9wgLAhyuYOf5XlqImXfho
Z4B2FSZN1vpu9bHqLz/5kayyXNtZ+MHYroLVz3ethizBZt3KI8AQ/3vcMhgziia8
YEqmKmRBXuWmiyzZP+q4nBKKLVzoCzolu895tS94TZQsBwYdJ8SQC4ipk8lDHl4w
AzcwRn6cqMGGmMrQeYLS8NedpHSqYsZnNBS0GCf61N3da0pvWA34VyUvHIYOolhU
PZMyMVgvrvT5bAr8X8c7ZLjb0m4R3X1+yuZE3l1lYI3AS6+BhzQfdvK7jNJZdOyf
jhAp73dO10bdDDu10DYlMxO4Xa/UcjlDEZ940hHv0rRDljACLqRenRdsPWj454/J
Snz0jgPXX1uH5rtuEc4LwSTBsbyORWjnA7rxlZ3U1bx4t281DA+n9tt3RshdjhOu
t1huC4twPicPxrC0xksmi9xgvPtUKU0j+ank4K0nF8Ajt86LYBht+dwImup3gjgm
+VU3uCVDj1N8JTUjmOALSH1bZuBROVp5azNHw5ztMPb/oS6TU0nsY2ILvWaEp/V6
bV/izclkDlSuQVBsdmjDABvH96wQ7RPrU1t5JNudXV2A7w4bFLXWcuYZcM+UAaie
MSMhsySZKvqWK6oEY2fLY4UH+pSMhYLA4YRgXfgAzErxysyuQ+VAu6FKSFgjIN5X
sioC+mwQvwAJe4H6OvUTudiXjt6ep5HHVAJjQdr9n/M+weXK7k6uY+TmrqrjBVsl
DlbJ1/+bYjWLqohd3dkPv0BAbjx0Wj8uCIYRjSwc32UFlfcAS6OolY3G0CGrTZIS
VTMJYY7Ng6Dry7kX2o9T5L8wULrz63iO3Pq4RcW68u9gaJokpIDuF0cH6XCl0bSy
PnqVzTOiIlaznUSsSMrnpkYjf+JG22s8h6yQi/G3Lhvjr5nbDfSt/8IYCAQKmpPW
9r/uS+jH4eglOruELUdY7rHnZgk0ha0E6vgw66LP4idylyI+Oi/41KOtymBPsoWz
/I979RRSJeP7Ja15FeLGbxQowbnAMyJqabtydD57ZDklPOykXdrv4ZWjqBTShrCe
Hl/PJMTaEsvP/0QLMZirvQKyyHSEQRWOShyqvdEdHq0F5B3lJ1Xd0t3lPL54nvlB
5LF2ovW4yocOqLRoRwN7OtISXKAai/NKaAs3nDZxDNPto3skPtN0ECJE/1ljl7Wn
WvWFgSuhn6Q9KwYXhUwCtHWBbv3I3XcrGOrXyJQjNu/52p0wh6/KSe8ThtaZ2ym4
5nyJD4PAgmFHs/It+ZaUZGhULMWX1kFh4goiFpO1plo4R9SXToJ6wNfJN1fln6Ah
6upR+O9p0k/iDLDZVrX6ppQ+1ZEjMrAhVisZ7HMcGdEcru4zv4q89Fzz+xAM+NwB
YrrCgrpLJ7jUhP0QQu6k2cQNRITgncjzO0xN9zawGH7r/hGPHQLCSvmnOPB/ZEO5
Y9B53fdxl9DlSbLDPpRT98GwAolC6HKf74azbRki/EEFYCEqtzre8zpHakoLeYkE
Y3ybQKQ50ilTbl110u+/27VEqMWvw1UFE02vzn8HxRhngzMnrNolx8R0Dm3cJVAO
xRLXUQHS5MrJSpVGvvQtL3vJf7KctSf3/K3esFh9ClzyzVTNtkcocoh4yQ2kqEgE
HjW2LCQbsV2fMR54kdU48eVifPZdT0+yzYcqtmSXiKZBIQ7j42KxvINaOjaOFXOn
PQ4CdxOJemqkvbye9t7Xj+Zqc/QYLhNxGflTsKn/sG67Grrn8M7vvvxWqxYO0IhB
WJvgf60fPkrO90s25T4e5+noYPL4eDOfhpLduF4gUFSekdxd1VECMCGXs37lK+aS
bi2PdEBTvAnc1IGUj+jh1pwETop3h5Vdd+yTs4SvzPw3M8/4qh9FXUXiYpHoiUUK
XHJBHGkot1UTUJW0+h3tlrh/voAK0B8D4OqySG4gZ84kf6nOgl6fTiMAKHeaEjGl
0Z0C2eHb7lI0CIWC+vW/6hhYmbNYtdHsgpG/Lntaq55K5poEFXxu7ek8C6Fn/GdY
ajKSmYkQmeD11CDTq846SRrJ7rBiKdz4H/GTrAmIZztrnWaByYX7xhV0MzZ0Ggxk
9QapqQFg4p/Wa3M6t+uEv/2aiOXzbbKdHNoEb0zQ87lvaJXzMklbYUctMPQIfv+H
L87l27tlILx+pDwH7FUfHcZUtKbAuLCD92wpvJtzzgGUzvD6B/lJLaPsGDzbS21K
Q45PF+4nZP/u5uDQMIXBAl/dmpHC9LOdX57CwNv9u5paIQHc+y6j1szK386NjoVH
mli217aRzkw12xZ3uVVJ9LN65H4KtYWHc5QdtCNYOhlco7YwCt4hwwk1i1hV9hfc
CIdySSPGvRxcng+wrB7te7u1BYg5anjASvQrcQHjUV1ljQu2+X5nShfvCyAtRsRd
14sqDI94xVfqAa4RBTc3Zr/6qJi1ZBk1GOrC/9v8jwdzgZ9ZxrBbQVoCHUIwr16h
xiVaNgRwwdO3BQN8U10afoQDsNhjxPDcU99oM+ieNpFhkUz5LurGyFnYqzliNxja
mXyJT5Ak6sR21VaOnOUDhYkbZe5TX0szvYfTrnRJVe003+VALyE1BeBHn7jXnfTk
IvuwxvoPhINCjvcMezqjvkmUw1MA3h7IfnYcW3EW0LEMliFiIlqsWtfsExgdDX0v
ogviMEXYTnl2LCghdeiQ0GYVQMRk8fC8KCIVOUqb8FIgCBRcojFR9t9Xk3wt0ZdK
8yDlQRq2RgdsIOMlzOl6hWnNWArkvWnPseMb1JH+n13TL7WVfsXRONJXMMcENyGz
or7z2RWfE1f+Lrx8MRRv6VjRiKnUlRJqTbmFt1nFKWMct7w5OC8YEjo4GfWPbf22
XATcUiNXsKCqtGbd5coQ3iTlNiLhEvgenhLXiRQEmtimB3/pySozNI/cWzpi/pQE
qo/H80rF3hkgZuNhZVRCaT+duGuunAZGKfJ/bJdp+NyX8GR8Mwq1VGgJCqDFtNO8
sZLO7IQW6tcTkfoSK5Rr3sr54AFn8r5uW+l9b0AZuDCDsELHSxiU1Ag2Pz3wFpks
JcW2M4US4k3PqkaNgjB15e8jhVubqBmEUg5ciUWsGWF7Ko7INDvmdvLIsaWxgw/x
11INl7YQVgnjYmgpnPtkf6RjnEiwQgxDYIY8u1A70GQlR+mPqfJX832rQW/dot8/
2lZqRW3/sG5/mp6ze1Ee8uXXD6eZVgnLyUwINatkO6CYpJtkoocQIGA/HDiXBynq
6Ldkg/1wEEYsKvwtWVUKYgNut4+uLKN22f39Z4RzeYWLbPZzxb0ETQTBCWf2Pfrx
QtaenZDW5gPGhEnEyXCXI4G4zyRk1ZfdcIqpJuLc5tec/KCgbPVSllPsb+jSHr3v
hgPnmMdItqK0YPCFQO2DO7Yz7cOmo315vTtM0S9xKd+eOl/fjZXmuWlKQsojWeue
PqNv7iSFLSbYGt2agNXFZSBerSKcB4iZU95qBbKlXkSNLlfUTKt5k5w+c0cZDW8A
72PKpL5/O53Blakls3XCtBVeQ+1UGU7IMLSQ6mnN3svuEdtiHGQ6pTBO3aa49H2i
0IGo6hdId2f1/ubEbHphYh5kNWpK/ne7uvk1YRq+eui+hwf/++rHpeRX9Hla48zE
FGOY2fcJG1BowX171n70gN2tWa17IuROPhNs/xVPJLiTExSqbjWX9I6o7YmtMDOD
R3KHRkQTKmOTxa9mJJqJFf36hAjGo2/kGW3n4aPuc7Tpr+WNeolsrJvyddSdgJE8
+dNvkHtC5EQnu6iGXZFZP/Hn2B/WwW9pjyXN5BFY4pZ+H317h7AmPGAiR/G/zqYY
SwOQZWBmEsPfj6s7mNYFQfJXOo88DIhVdP/PWZxLt5Ca7xLKgooha3owKji9qaan
XsZ/WJqiU56wlWaOx6f5hP4vdIJjBzd4iTMxX9RwToAw9HUONAlKoTqPQxnVNMQf
vtB6pp0FebXCzQLK/x0Cqvjn4T6pye/AXUohHI4GemQ72MZ2TC1ik30eDDDDM4tF
7j8dcw5KnJpd5nwzH7Emmc2mjyLMnkE6BFmiBjiwxAaums+UfqwVWOUQFjDILGe8
klXB32qwf/W+V9YSKrWK3MzAfp1DFUZ45ccTVQaGE0EB+I/l5gQuWnErcalIBGsI
Eyb5XCCdNxUzEQVnnnKvHH93itZMXsSXc2RxuvJ+V5Oo8RpW6P+5dcB47Sv1vWEq
VMGBMp81nrxWTk6jCPK7B+/aUm2r7FmnExqzzJhv6a+x+8/ngg7LTUZS5K9+FkpY
L7Mcb4QXvuq8ATa3QZZXWppxZTjPsOTNTHNWUGQNrElbMUeVmqYGYguAA7ioaVFf
Ilg/bfrhwZWFugV1xjBm8up0NSiWOzclU2hlk7LmayIEtaR8KJ7+uixbnsffzLcC
9dPRPu/X9jL2mZYGpVURCWvC2c1AZDjydiGWyXCLUgkSZuuKBqFfItmNbwxOgN+a
4mCt4FJSG/RGn44pTFuhQYwwmTjFgY01fhPJxisKHMb1kMXr9UFqR8sxGjbfbNpB
mK5HtKSjR/WBt/fjuWXRz5ESF51riQ2IxP9pmgBLvv7JA/0NYtRTGLbTn8E11I1V
9ZkdGVb5HjOJQJMSxDfO1B6TpKoqR5d26sWkIcO8Zo9jXPxnWil/WJcFgH2HtDYu
wciPLriRT7wUmjHwlcRfld4o/xtA1JcM9i1c/S7QSuAct0wzDstcmpW042XW6rVv
o6sMl181bN666I0+mDKF2JzfwOlc1dm1QULwlrUJL8l7SAScPjJO//iO29G1acTI
BFP5K2ukuo3SKEsWT6aKSAZrELIt1dkwHb0vSZWtH1FGf2HlQwPkXBbHYdZQtFV8
Ql78RqiWDH8+PF9QYAwTMZceOriAkQP6teGPyLTdwe8EzBfJzKU6+dwPWU5UdiYV
renshULrnNKoEMAMJyl47xGVgERwzT4Aw4imUrR9Ke4OMxwGpvjPBFM+SVrNW1Sh
Vc5y0Z+jhJvsecJzhdJi4Eet7bdUZmVOXJlDQ2dGCA+kW4TiD+wbrRNLN6DuMtcK
LyC2e1B3CyXKmT+cuaDCwS5B9bHe9q2vpyOS856GbnwQiiqxZH1wD3Rohdw+a6jV
GbXtkOEVWGnEN6gN3mRH7UMmkm3UqjOWPQ7snY6om6rSAxhytcwl5BJWHzEZFNr+
lM+2k6KzWLeLJSmMDNv8+ySkFfAWVEwyIKOtiSh/AqwglbWhlW0Raj/T2yeFUcLz
QyLUUYXkXH8T4JT1EjrIi16+cgtqkBl8DihkVbgQtxzC5VjBSxwKLJX5LWbN4DuL
4QquMkYMU2sp9CyTEnasch7bKVgF/NpnyURhmUFx/YkC66alUgUlAkT6uIE9owMP
JH9vHRsSQlCHCCn9DzqgaQAv+sVy1P2MRnRZ93Rbi5rEh0fyfeuUdLYDhi/pK48z
OLNqbF0NfoZW59MBHDhljXZlCA+vopjpACcGbVXU+Pnhq615um2ssAFnudRs2mTB
6PrXHLvDfdlmIZXNQ0pXbzzotCsqfTg6N2rNq8p4rUQOIPrHh8kwthsG6LDSDCuf
K65qk0dThuFr5iOIM2GW9AAuurWFX5cRC+6280/gsMhZDI4p5eiaDy8JB8RJ3F9e
tIXo+20i+lxkw2yugZPomcdwg+C4xxgMaE12PicxF5uTD9gTwmIhZRcB0770CtTJ
jfrAX1ZBe9LDBL0StJEe8rT90KP23WGuaRLwgyx45GTnPPD1iRaQvA7jzT0NZa+z
7fz6OC3r05HgiG9WHJ421oWalQLjRzjBGZNrMKKQoEnSOoP2sSJgFV0Zlpsf2W/4
4KSu+9sLAGM7fydAzuiH26SLIUR4F7EuWvGERZMKY06KLTVXRRJ22royqsNnmTq6
i+QwYYEaBU10X/AE2AnjKdFTD4OG8tfS2pgnNdfC8PXxRJkT1GeVqFAd2MJeEzJ4
TPJGU34QYoXWxGXsjostzZ2c4OFT9VN6jBi0TJTUmMR4rMG1BCB5AL+hModx+pKy
/kEakljwGf5axBTTLL122XV9gVuuelTK2Yl7+mJVscg7bnT2o5ECz/Mpkev8LRtb
g7k5BUVXWzMFkiq2YLXn7SJ0yzirSfXVkgJDYAsasZWJmVJvkSk1nzCKInFtrAkR
ceBjm3uhW+96JO8BgueXDuNNXncYoJjAbey3Jl2aDLjk2SC3Wd/x1poBq7+wRilm
QF93BF5sDutS+fGQipHsms1ZXwbWkc3mKCph6VD6px37bjMLrsnUT4k5lz0QF5tC
w/w6IrX689wYR4QOeNN85NV4G+hbF+DfJXwJffFlw9023fFWcw4PH62SQyU5IwyR
DHHM6AKulebxEY9C0j90ELWva5YcD6+xPLr+NMywkg4cBGzii/46ow/jBTbD3Xk7
9+AdzRhV1Ofjg814nLfuCxW1mokVzqb+t1NCU0Qtnp51Z5RNTaGglGh7LUaizVQX
KByDUUmMCkc9NLhYmdj3w4KZBHawWQS5D5sQK+2mCii3F2A5A7fm+14uRHlp1P8b
FA+g5lxNNp9DwD6eGvKg+d7xNss40BymMKQrHtaBuoFDsOWkgnpxxArHtjnNvH7S
k3ZQDnawCjdDNNo3DEQP0CQEeMm53SW56EvjS3KiJbUnpp375Ud7RXW8BJpPlf+2
pi6XpodbLe7L5W7j1xNQVGnVlmMcT4o5xLpiRIpP5OJup5U9hyPkigmIzLQkNzW3
/ns+5MU2h5J68Jyat6a7Iou8gMC0ZCuniBVvXAo2MtnMMWopRsLW5/Eh9/OSlZCq
3DothlpMPy/XVtmO6d+n+ExuZdJUOAHzsdg2EL1rrAmF5p2vPw2ymsRZObMFY4F7
YJt+6VQMh0/gzffbKjIeIo/P1uOslTc/+GVifkB2f7SFOepksIQNtBp2JVTdSa1J
zfpKUoeermQmCe0FV99e8dn6e8Wf1dLMt9SwxtXmEtqqsE5aQxGxtLCD3oN6XQgb
iUgOiamIBRtNhxQU7MFeCUD0omvJu8pIWmVT1GyFN2fn16oKAnTDGukd2wl8FQx6
Mzr4HlG5fAxCuGbPmXEAEN5qF0o5UOIbFcDREEl91Oc9DPIX8Q+JHiVw7gK2SeAn
q9mc0aEPRKC7dVn5LcXw21Q/4IyEBRwdgg/kBZR6aUeiX9JJultpGBq8O9VBBvqp
uHh4K7cKsdiH69kyfcuIQLqdAa0S+cgWFRB2IGVTbo2UZ242GAV9Hd8Myh0UMzRg
rPbBGfpF3rw3Gp/oHdzIkcHPDneSnb3h4H9oCNCG6GUDxrmxzCrVlyd6ei/jxxMP
2+nu9GOOmhUiHCxregemfENQBb8rVegeo4Ki1yISF9/AZWO3eGguAPxTyBu8XCwW
zae2qSS7m8+ez6hMKgaN7rHDdw6NDee7hBU2aw1bhalXEzXmEIazLjn5xfxd/vnP
G4kniqacYv0xi6dKCLFznszm5OhGfMaB5nmuxfT184xoHvrPPPRKlfTjz1GZtpUl
Q2iAqBZ2V84VgYuIFxDpAu8qoCLEZCCVoqBiIP41y4yEPLMlZyxlJ/6C5ke2NZv5
5jdFBhPLP3JvHC5YlTI5mEh4qDiGHL1AVxNinbZ/arqbCv/VYPafgF/1sc7Sa61L
JfiszKfQGAwk9asqug/SYAeHo37dGVkuPgUqhQpVst1AkrT9XriOUyIxYfcvQWn3
qQiyJ/ma6cpsTFSJ3/q1k/p4bjpPZFcANnkBV0sGSbHSulgSBfUv3wFWdZmuqa5x
gDsN+aNgERqJDgFU6sVBN0oLrQZ5FAk7IHpNYOMojUWsMxZddcYYWgahcPRH7mCh
Q9slmc3QJc1Iw4QJgFai39iOPQruXnDhQ6L11hRNR0zxVlGFGwQfWHaQ2m/BrZWj
f5TFdvahZEbZmQjsJT9u81GJgzHjWJ4jNMsvWU+DS+siCyw8mNVEFfZPav3TxILn
izhrrCosZroEuemLSxA7G++Qx68J+eagh/HNzYCveA8GQ+DBPHLzNpQ/i8jGmPLT
/Lu6aG1oEdIN5J8v779bslnM+YA9cI7YRTkJ0wfBlBQiSV/0dFP4XFeOC3dZx45o
wtkj3fD5l9gFG+XStjwGhWUg5+Ya32AGttshymlpxoO9iCGni7UjTDJO+iGHQzpH
GpoxSHuAUNegp0ZTbGZW2CULGKGjvpQzABEHCIsdwBFXVwjGqkdh9MhNiDErg3Ej
UFFrYbLRQw20K7XoO2vwjEiDgsG10y2+0jVBJhv1cHxX+Ui5gdqGvTh9WFqfMqAy
pMiTwERjiLRWCKv0L3jxxr/J4uIViIObaEk1MKZ47kLNZIp9QhfjGtyy5UEZyDvu
UHK4FM0i53YVdRpkTgU7XcREtE4dGWWuyj0SiPHzYdsG6HWebI+vmbjznvj+FqAe
I54h7GUfaCqsalWdJKJyMqEWEIB892xCsN7NWsg18NXe7eDX3rUOUybpaEMjTI3x
7GULKHmOmSGOE/WDcXLUZtprcX7jIC1h+K9GrcIwbc227CJH9fBQSVYKeJzP0N51
U0glIFvRVjTjRMpnhDHArO1okeg9MjWUsBHynymd13CzFYyAr9Hl6RWNi6Qwfiag
STqoDpM8tzcXDwGBZeC37UetCpNZPK/isepe8RPYTIELpdMvrSdZPdgRWi2xLso+
Drh+SLaoleh12CFdZk90tleotVawiF6bgTW0oVnZQRCFU6o3uRmMWtaK1UXoiV7R
w2uV6fUKbYi06L/T4HUA0YdfpUlwzDehbWACSF3HLSJ/CgjbuA+ivEk7/Dkt2URj
w7VC5ezA2v6CplpyhqmZ/pj5nWPauP616myB9i/+3LmXViE9Vbc2qVGYgE2cc/35
HFh2p8Ope++8WOXM48yDreGfqWztT4scQjz44pXrPHPis5TicZtXj2Qg0kyRKWz+
geRp8X0MCuJILetmH3qSI11CMR4b00/CWRe4bmy6eLwi/sLPMPrcuofjuGTQcjJc
ofW0z/zBJshMFaDhCGC5Xn0Cmk9wouLAZllbAlQOdJZqENf41p2OX7qEHWnjR9Hq
XGm3Oj6D8nj+T+h/niFrZmW7V2swdGlbyEAeq2MzwwU16IHoKvGlq7MNiJK6SWHL
Ibzs+fa5r7uuVK8g1orEOj9Yag2kDHiJmbWrbfYaMw6hISBgS+kxTZNc4pwXxenB
svauSEZlWM0OwndHe8U+DCribp1kmLO5lW+wYw4zYJMIDQfrG+R3cVZo6pNBsvtc
Hn3scC9F3kNLTVH9K2CxHBRL35+4rP6u0T0jPGuREOQwFwzDzihP+T2aXhv2/hyz
UqjX/5qxfTBjP7jLsblLefVI/AewJNE6drPeckv5VbLVahREWcX3RE0XVcVw63Gt
Wgx66+6BHVSzJwxd7D/wBbn9+TA7IR5/rzTYg6bHh1P6a6UjjYRGwv1aspV3wN4O
8XyOaKHqmJvH6PeZXEPXSBNJzsdCJD72XWH2Y85rL0/3Jj7NgIuxkz28HcmGvt5K
6PdJXwqxAVErRZkU0QJNBmNXr7sj0IyJ/a95lf5TODosxph/WcmlnxmX+dw91VYJ
6EToXYnJT6eP0WA8dgcIWBOLl8uVN3EoxWg+luKHpBLcpSBSs7B7RnqniufsAlDI
7gLTT+4szlOZl2PRxWTgO0aRH7OKv4131RTqWhLXPRtqqqc6MV1AIh/+ZDeQM3Ok
gWfuq2tSR/35iu2Ax/jIOqwojShNO2Pv97RlbNa1G9K8ghJqxKqXckNJsa9bLDpP
uQPMZkYcHkyIUqn0TQBMOwsulsGNjetPIfy9YrpfiRdGh6ONhq2RTNLJ6esaF/21
W8jH21BUA+emrpTY/zwSATYT/LbA3USSFDipz456/jh9AuXZUA5gXwgOnyvaGyeO
W8fKXEZ72UJD7nTWiEEWeJ5W63uzQOt201G9dfX8NnmQlIs9MHy6Keb7GAbj5oac
C+zQ9RFudKnpUfZ2TRyyHupsVTiwRGsp+pEvyqHf004a4WHB6Bv6IaAPy55Zvu7+
49nPfGUEHbgsFtzHJEULmazMfxEUxLdcSWKgcOM0nE924zkOeJ+0fTPamD4lls27
QClhboLHS8aseNEgAGt27epXl5Imn03tuXi70YjfizbbESqu+6o2QFgGjyRJxiXC
3Ozp5e/ay9mB6ry2iLn8nLYiv65C+Tm61BjmTMhee0uTmkMAJrAYwi21Skq0Ufx5
x7XxlaljKm4q9sNspHpoQTDABgMAWcnS6ehTeApUa0HN7I2nHIrzxJUD7+M9RopE
HvwhTLHcqI2DiF0Oz6EmXZJAej5vg0MPW597sLkL2gWlNsfB/zdhbv0VtAgS+lKa
E3vJFvdg+1oldVQAPd+ufDfBQkC1V66aqI/vidV0re200dqtuN9yt5mDP65IYjzl
cpvXGRU0ieCvquaZDAY6o43eXgqcZQlzOCbplDc9nkcqMEGdlMuEnQJN3XAA/8lL
zjzBFTMGGfgHBHyD5Y2B+NeVh2VMuT3sLwFnBouPjRi6zWqfij5EgIT/atPSKBtE
8H5aJ6ynXg4OraqelPScVrGlCQMgTIYfZyx3d2Cwcy7IelGbbam8wolSNGCpyc47
Kze+AEGEgWeFXnB9n6xAGxWTI5yWfg9QXyBrEjpOmDEDeO+Gl2zlNLikvPinHclJ
x3qWZqp4a5Ghm8E5GAvO00DcyMJNID4ygTWgoFHNIWnT/JeV+XgRKDeOPoLyAFLp
B6BICxcPzyrm80iQyIeW4jDDciHknYzBU9b5fNsZvrul2JuEB33oiFh6/R6i8JJx
WXAkWCJZPi7TZw7rrOl0w3ZdnGIQYgIYUDocDW30vzqAbQBbTpEXcKZ3vUT/YXgP
cZ1Bv+6tt4i3zzCSr2OQ+9UdezAWdLITcCdkSqZhwd0QKKnKarG8mEjnh23lCJcd
6xda4oSIm3ZRXMBKWdCjg8npYEtq8ZPDWH9QFsnc2WTcHFdGdRNQ50/PN3MY2CGM
knsBRxQFMVek4/3HGw/0yzaoV/5OwKVIYA706p8i0uEOuKoeswmJIeolYMpFDk7g
k2MtWauSsLvi2NDUdgsH1S9RtKV+M8R7BA7wj/JGsrNvgJFA1OBiZe89mN6i1Aw3
bAAyAa3ld2vP+L8L7lszVYM99RPthQCkvxTTnvqC34xTOjJ72hJ9feuBRGtpO8h0
ICkzWf5N5cKtV/IW4jCjFnw/X9e4yuVRw7/JKI8DshajwAlkLO/cMRFs3VK16mQl
JiMrXYuJcwkuWu0OQYVvH80g3GQ3fv+ce+AvH5P0QCEe0qbvajy0AZO8iy0Muhor
vTku2pgeC5js1qTAd3iLruyVVBHqeGLHpLiiHyVz6sw2+AnPfjN7t9XFJMqL92NO
4F1s1eiGnWGYsgoJkkHNSXywQsXsZXdhvN3Mqv9H7myIUa9RMPKKDO3daNBPoaCX
dyoQPNNgUWyTYxBd3pF6MiWdLtdL9l0mwax78bQ6U3yOXNGlhkDzgl/Aki+bhTre
PmVKqpKcYS87OStcyfaz46o9rH75a0c5NPrsKeweEOcSJO76HMnkeWcJ9gPX6cux
qHfKCfVCvBt2iBTbOy99l3MQX14hTJOE40lMLedGpgtxld+9xBWWLX8ONtec7rfH
rxhxMeq45FlHL6EWqzZ6PUqmT/4czXTbTt8OA+k4AzDXsgjOi09FN56yXy7nRWB8
WR5ewlZYzk7eJYR/S86yPXVaWXDxPekVdyvjbFiTw4oL+wQA4q+jLEc3sACt5FZ3
BMPEqoLWmuYlnVgjvmkQJk7K29CjYSWTnDwozT5tL4btngANXW/vyBfKA2nbxk71
gvwvR1gDgqI6RsLw907kg+qwFwgjpeW6zNX7QcVbi/9Tfq3ckTFz+9vwuLIgHiqq
sesQj6RWj++ceHKQbuO6LGyY6pRPCIIF0BR2byNPLSJe0hG1LEFES5+Nz8uZqgVk
CAqDmN5K/WY9RGkej4mFv2bivwCHtOAzEaH+1RsaF3iOgNkRlluCvgIiOM9Ce6Dd
jUU8+BF/58eQE1wo2Gf4FqF/6N1NyQ2dq3VjK+UfDYlQMWKh/Tdw8HXzOxZnGJ4/
g9iTHthi24UUgMeU4mXnNc8SSRP64MuRHW1b3tfbL+FtbBix3uEDoi8ePXe5nOV8
rbm1zPTVhqTehJw2ZOruwIBLyOOIjdWqDfZvwgw48OddJsdYXBmPLkNCpb/id7Ac
vT6pxXosotqwgRDMplwaHtMCZ3NV+919IyCn7m3Ab5GOrZKZVz8M5xHHd7+U98hN
D8KgZt7cbvMQYABfzSRWi2NDpxn0J/OpTz4e3GbLuN+DKEzsSmOy96oz1OE86s0w
VjoInH8iIZAu6FMQ8ULKFpMReM3roYRJfYYpTPKOhZyaRyBbP2p0x594YeApgOlZ
EgTpdk1vOJeYtRbP57mlk6cBPXDXsnX7GbQRAYpAEbLr8xYSGuH2j1z3A5+WqVHb
7hQzZsCTuWHQWLko5+5b+udLQV652G8G1cA5nLOo6WfQjtju290NLxMn4fhD6pn3
+NON9DZXLHAnOIM0mC/uulHFxuEMNrHMHqqgK22yU64MHR8vLgD/rg75r3Wu7Bgk
HYgDOG5UJpzkdLUYBO4CNu7Fkgq8aefBJ0eBpl5SPTT2UVu+Ncc+SexrX+0IQeNG
GcELoqq6Ephlqg6w6R8cjdabli/Vfu2IWcoaw8ZuOiDIggMfZD0uSO5atrXnByal
D3LKlVrVrIzBHocVfJhqKkNdAMfl+py1801L8ePDJquS+rLrWS5janTJJ+bNnfz/
d9YV2Ns3ri7QMTLxDTWbVJG9gCSoLmOqSTEsJtej50WtbnuBlCP55EnolbOP9xCb
xA3QtGH2j7WaTFlQIXEuOqb+/MA4KllN5dQiOVkGId8dgS5Zn8Yy3ocYwb6Tx5Fd
a8dkjs7CQ6Vz4nMOkPm6QTCA6CLBvbCyVmgkLPLvjZPz5WEiswlr+rfG+gjg59aj
0tVwvXh3LRvdptxuP/bWfbtHa2xSJbB5Fzlj04wdI0T0EdYCK7nwTPnkSr9IXuh2
kqnrFoxVmRuMpiU9pJU0gUjtmfvg4OccPj0M0bXxFTRJI1fHZV7O2TYVdw+5yUYA
Tb0jRcJooY+u9tSAltNDPSDEG6UNTP9Ycpu76DiqpByMEiKiPxLQaYDa/9yulZdZ
RmyCC791sw7yVHppu5jqZk8pa+qRDyYJz0trztSVv9vxrCD3kVHlxJ4YaAPV51Zy
4IogMGTu1oLW43xOoBBOVStsLwHOT9l8UfIoLvPCPGICKMbMKcDBhQCEzNXpbH9j
KUV/3odPUu4taW1qO93wrhbYJ9NTFOKGm4/9a/67wrBa4Lrhz7n6HdMEN7XkXskz
Lyf3Ebr9EzgaGvzTKBwpyHj1B72IeqwIfMBGXCddMaT9+47+MXWS1JrcwsNN+CKC
N3y9WLNI7rVj7G/L/C8kwkjEJ63srZdEN8Op5QLy1GRVbn0uBQWUblPsrcbLtDyl
hRZFzRkh1ToEka9axrgTVgrCmXKoJIxZ9hANCVvvaxT5wJm/TRndgAPfcvUMyQ+Y
AXjnxzcJFUYASzQjG9S8aYFyYsorcURL30wtuMcXYETp6FGtuUsqrAHFuIa+3YJZ
JKWBlwSGhvvzWNx0PpRq77zfmOIdNMQdh+DxlNIGo+MARiiP2JVzU2Pn9Af8ySGX
xIR1VOSuzDakpha4qGO7WD5hR0L2ncp9+9K5eJCHSu08NVy2j18mlY9VTV8tt96z
fXtAaLCqyMI7WOsBlrsM+s4gWn4u3AgkWHR2NIQR8tAATfHtQsazYAbX8mlSPlO/
dR2aLXgDvYqywk1F4W39VGgL5XQFp4WvC00yWINhd/WnCVFFrBILsVIVtkpsq5Ch
+0V5PgfBmnaG09diW2WgKd/7N5GNcg9CXjGfdG0eUPe6qHwn3+03NET4WslqEu/v
oohoaDBF6PMUcSM8LGZ8DmAG7dQxLU5aUkv3s1qDhJOVCVuJEdukRiOtxhO7cql/
/gUN1fqvbu1Dm4wmjs7aEu2jRVj5pok3xtujBMMtbox97PJWdB9t7U2oBdx5WjyI
RDQ19S5c7luod00Dy02hNswv6vwrIcp4SCmxPG94+f015s3B7y0v6ANN6Am9gsK5
PGlcxu4GK+SRgjlti89tY/6QU6XJ3X4bRmRkjvzMlFp5k56cSYIBv+5/S8htDx+8
3PAp6qSYAeTUqBQV25hSTcXXbz08ESecjRSCDS+H6BsYBOEjRjAWLTPMURzvIxuz
Lu1l/0kvWlafYs8sLgel64oMan4m0+gmsJDvnY3wqW1FWkMoqOVZEzRDaQ4A7aCC
D8YJpUOZnJLd0qD+9x/bWeHzc2O3HCSp5qrhvrUID3qSYiBwBTJu9iw6E8R/0gjq
mQ7/ixDcnlTGyRz6u6SOL41WGaQBGPmlLfMBcnE6enqzx0vgV52dvz/VChtINnX4
nFBauVwI/fASNYJb++5BL04nGr+PIWEpIGYZHgX3Yi10pOwTwKxZ/3TogvST1rAG
J0zaEqrZxGHxMjwq+uljom+GrADje1LggV+ZpzjmWQ75eN3nQpObOK2+nTRLP6v7
JUdt3nfHuQQw5z86oStq2R5NTy5rY3EZ4HLR4vI+JKquoxa1CdGURJ92c9tctmF3
XPRGJeyZutGkBE/7snu1bRh/WKZziTDm+t6lfmTA+sU8o3ugco32V4xxUMkG45Vx
Db685nFcnjNeLT+t/RybY6y2j8BUU8gWwd0J6VF3E3kEAhz7NGLjGLEAyglmQbf5
z06AjGTSpjAPWFPI5jq9VvIcFlGWNei688w7Z7FSXpEOpVVJYCZJmHQvnd3rDYpu
LNAdpOPTRQBVxtTkl1pxeDxYtHl5WXEOGIXH0hMUWeEw79y8jTowD1wphqNB0/CK
YcwckdA9GmgnUgviWJsyrurgwRc2ZjsHXtW+6Y2CIKhGfikHfYrXzymIsvS4UmzY
D5jLZVEDidRjlV4iwdlmriNnqLvfHGK0BbcZl+OLKR4lKBl62fNW+5bntZEpNzWo
8zSouTVIrz0jqz++2F9QGEAz4pEiiKiDsWdrgN9T10+DuMHl1IUxMTOoqEHhENPW
bF2EHLpW/EcMk9QnXGTCEE8nNIAmMEvV2kdgr8nbnkqp6exbwmKLzUKFtoEKPziZ
VtxHPveq4XTcfySvBUhYvI76OADXQh3qXV0AjXUBy6rPfBw4pVt5pYZdyo6jnRs8
FZj+8qzY904Nk7UeivSyd0tv8eTWSv3FdiKgUA/hGhVT6CJdnHPc88aWzkrlDsH7
62WjyZEvFBSZJzD51CX6bwkMvell0RgWFBq3yddWbygMQfzANen1Q+2nLJgQsLNl
Cs3uwr43mNC2wC5c2d0rHGYK04tNp8NjOS9zo56nFeI39bG8GBjaQKWqZmBAXx3M
xuDQXJEz+C2rpU0pTZGx3NPmfhO2KxDg+XdS+eXmppZzVc9EMXVDTCUvqbgwYv+N
fiGzsoyy5rYKtX+LnWiAP4c09mgFuo2HU+2MaiwuTuPWn/iAh7xL7rD3X4NQoSpR
tyZBam4Ks4RSaBypX2ru60PRIcDBpw2aZUCdAScRYZZAcpSLlytOwJQ287Y/nVI+
Mx0Z5n1s9Ou116OlmMVlHOPGrlTdZuZWyw9BEL0eAOiGG8zS5T5nhMWSUVX1ZyZz
Jja1bJy3+EwxjkjH+/kYg+5yYvMAbklkoKLRqsTS/NEKZQ/BP4JHR2npOO7uM8vp
UvvHeqsBcZeVq/P3EQ4tK3rrpDQVfQcstPOKrvRxICHE/QBHYFkNR8wUOOPokJEd
2Fkt59yFysTvldWNhK6Lb52kh4b3s+mV4nsOigJ2HPzvESzEyoA1oDQLaGLH+Svz
nnzFHhltmaHWPiJQpvgV48lI0z7x1APF32XFYIQYehez0hlmJGWPwlplZ5Sfe7ak
YrAqH/JEROwoLn/QDNCyaO8MpncSqOtotBc8t9cXefIsJ4K4ymQNWfmHVMsOCQCf
vcUrx4eqPqX2JdCocfxCSgVfnqYxSXjUZBZcTuKPaADS+RXdXYL7I/4pZ0+z/NoY
7k1EQmy9Kc4BosXW00Uuov+7syEx5Z1cjzFzDiZTOt3nSNqomW9qtlh2NUmxwvAq
+Eb6kGmpZ5FhxK9ATBB4BrPhEXbjW2EmEq29ypqZrNqzHvn4LcGYpxxE58evKYWd
+2QugTx6kYrqNpsg4FCHMhbfLm6Oprq4EmAbHfNIxuIS96fOcUrMj83cvNU3X8yF
zB3BRQiEAS4B3sNoEY9WLzlSh5+llh9ge2GjRUtaRR7TC8Z5H2C2UQvIUQZ8EgCV
coKLTQwnghaD1OyIvC7dYiqEVSgr+vQuQQ1rdziWvjAurWedKmPfEktRJFx39b/T
LIl6uq8sDgyZSkkbIIiK2jD25LsRB6gsWYSH3tw5nYghR6e8qW4rrLLAG8aB/oed
CpdVkCP/FpjRc3N24vuz7JH7an4a3EdvF9xP226hN78RKvL7JzBrs2CL6Fet5xRf
shelHSCoJkaHjj4K/5BVxMyUi7LUoQrSHQ2QrDyeHGw93VVCGH0VlCNAkpzaxOUW
ycdA0uWudQywlCnZZdZ/EQklx/BTYFHRI/tEw/WlJBcS7XsV1p6jfjz42oeL6jkP
uwUPLdSQWZq5Th++he73L1prKgbMb/8xb/wUXsv8QuQtN47v9YushRMtQ6XMCZwu
6lLUNf2HraOTtnAjVyrqsqgRA7LgzEMjDnjRIXLYzFwd6/1s0jNGMUdpqI7FOnOQ
qf2MNg76tMScPH4orsTE3pC4W5qxZodNtJ5cFrc2fES4TUYba+66JmOUhZ173+Ln
18LnoCbICBdaAcyyKsopktuGxikgl880WlF3rz+X0sG1NLIqsmqyo8Er2bhB2BNJ
lsdp4TnVzIu2KC/awbWW9QzRGAi3szFr8V89/anISMcxivi1Kq/ZELyrt6RPo+lY
ALetPRvcHydZtmrMMjizsaWd8zEW0FFzhq8wIydfyK6BDZJv8UOiQVn7dXnLTrXR
m5ntYnwhG51xieFIfkEHAoNAykShPBPOiN8dKH/MfHMEvGB85nOhSP84jLwEnk57
khH4jVzSB4sSP74EdmtOyM/G8iGklztRWETYm8+6lGj+U9TXb4sX4dlQ1hYUDtTN
UqQL666UecQnVsGxTOhHb6PVgn+H0CO8Nqv/CHsJO3oPMfKjpvbJp64qLksfD+nh
pLwjieLRqoCVFhjlw5jluA02rCMUjUTe8ij7STe8KGUvS7OiDrid66U102qyGGaH
HvEq6VcUPU0SUySSIgHWYpalV2PNExVz+X3Ieidn3hTYabUG5ERPSFR4/Awi584Q
Rwnz/+IxJX0tPxsGhtMewqrMBfFjV0DZhk0jBcIk4V9TMZmH7sbe8kRTu2cZ8HDG
SPB2YfK3u889sVl8p30IX2+xCFQNOQOfMobtO6lCzTRooxkGHpup5sW5+jERTL8P
CUp+p1kwlqTdbXO4i5tMT2L2e4p6z8i0X+ojsOBnHIE/DifVHAqDLvhl3IAkGVZX
Qf7LSqlDTUmZAWLFuIwDS5n/fTlxeGDICHcVuwU1ldLXqRS38MaZpoEdX/BTLXYk
YJ0UeKsb4psfD8riTnLxevvVrpy1pA3z5p0uKeBOKpRDbR9e3h93DIqRo3B80PM5
6k5NvWXX5agVFUQ6GaFExNYxkkAOA6hMOoRk978KFTOnsLaEP47chHwy3D5UWr7+
J19acSZpVfP8ThLTdiubfXHQ+sk3wT4xrAZYzjKH0eT4GR0ozl2O3mUZQYLAt08o
wWockxmQeAthX3iPJN18ED3qq1RFeH6iP0iCnnf6m6LI3pZBda5fJZg8S34WIRTt
col7WAJ5vcrH6XPQZwj+c8yO6FIrV1MLYH+aouRhyviFokBQ5sPxUerIZD/IF3et
0hqbpuvnW1TEfuHeMZZHGjo7IMEKiTpDdD8MvkY4X54oo6n9gqaRZAvG98WAWGgk
fgYlLh4xG5mOcJmbu3W/SRqSp220q+O0mn8lt5NDnEEtEzGZfON4mKqY8elvJa/f
oAT3IJPJ9/zV1rMmtvUdg8a76RocJsbz16762veV2APEVbsr9hWv1/OkksqGwGaO
4YEgwod7+Zm3hwti2eRxp7q12QB7DMtKSipVNXWgQ/zZbfp5mi2TGtLkpp0R666l
jel8PLznOP07x211moBCUqsmyTdXeIGYg4GUhpLV4ieOHnYBiQmVMnZgCLmpzMQH
O0X9tW5ZaRABtdxLRXHYq0/sov4cQlhhPVJs8WHdekRPMYgOnLLy0b7rmL9rEGUz
UrAhs7nl5qjI6SpwKl9JnnOHjKR8VGK4fO0Q5tf/jO+aGPBRGwQE0s8iYQvXylVK
8rZuC4iMaeFSiT/Qjb4RDDpiXdMZ7i/W+9gYsc8UkFq7JCxGQwGQQafl32ZF4Xwy
VYD7kBMQUKM6INQ+4WCUanf9D3S6qgHqfYcAChYvBwKQ6MZLsWtuWgMErVBaYbLW
hLCv59kTfGn3zVpEiONZcUW4JEYOlFVfbhzZVvP4PP+TvxHbJTt6vvwHpdP+Da6I
qwSr6Mq3xmwBO7iA5mlLx9AV0PMLcn1rE+fm0iRrdMlSoWySInTclH/f2X+CaeAG
gX7jkDlI5NHY8JSspfvsKludURmroY8qtzThNk+COH4moLPXWtbVgkZCt+R6xafi
MU0EAGK+HSn5DEWwHlSFiWrz4wrS0RW/PDW+4pewlpzOy+qrTP+aA2y10U5KZqyQ
3L8cGayoMOEMtDSmZQg/VdK/ctfIXJjns1wwktH+Hv+cwLAwNq2aLyeMcG5dYXu/
FpEr7t42gcW1sFcST1xOzhXsitPdupEFz4AZXil7UKG/X+2C7ciXiFtW2cnpz439
PVixyMCS02MhgHlSfLWpLf07O4cynVA3eddtnL61EEzMGJoJm8b8+09QKF/I/AI0
hcslvWG/WsCwPLiUPae8LXOzSqfmN4165cgQLzWLLlaQ4zmiSaXg1KwMDDb4O2ct
uixK5Auu/pFZaIHY9g6ZcjAe3BhkI/ZtUMkowjCo6jnryCO4Nd2WgntWm39T+jlY
wZZNUAK0e0N3RcPEEo9vROgtcnBG//h+IWv+oKO19SPbK58E6kGLDoU2GcslGfBo
l1zaMBcFLIzxuV4br/OUpwl9lcWtXx9gaeXWygbmbknLumoxHr/IhxC4mzentfpJ
j6yOJxQMfIwsLePe1lte0p/lyHoOjBgfsvosMbW/q0fhlV3fNsjZnNju35nPtbD1
0qJbWcBgT6TGIYAyQ+xPNuohAnQmFEz+JzZ30Ow7ElK7K5L9IDRlVSBM/cO+Q7+w
Iai/AZwBV8dOMY5mC/hnfhn7EIDqqq2kYGCyJXNUJMIMcsF6oeQ4Oo0UMjmxHheC
EGxNnmc0NqWS8FR3a9hgN9755zcQdRHjUsZXtXohGpocxCUqN35o3fh6lJELGwIh
pqCvQolzcNlWqtJA06ZYzekpVJwJw1+Ki2xqOFf4eRZv5+t6CI6D9XZiwxvyAoS+
HkwqOP3F9jin6Va2GgtQE04obVf/4mvecffvRLXaPKZRszHyHP6/XPY5e0vdX3kW
/+LP2jBcT2DeC7A/H7U543C/E8fQGVqtZu+E80EVDt6L7QqmQ2u+/wJO8CsKAhrs
ZZ/yUg/N2hMg3FurBN3gBnvHrlC+mnNpn2/SamM7lGf7EO9ug9VeL2nPE7pWFb3q
rRmDG3klp5b09UHm1OEjVNTEsmvm73rs30SI4L3BDNXWvvxpsG2y2RxGsr1sBYsl
4cvcjIJOSQxxNNdxpiwl1nAVeLpr1G2bhFLmMFUL8m5u7mIz4OnTx2NUOD/oauyd
Fo+F9A/T49N9WY3YyWkLGPNfeeR1m+f60AQD7iJ538MJ+9AkN8FPjvFutTB46TEW
igexvbQiD1PvvG5YYKBxwVO6Boffz3qzTIJ26VK6xg7qwXrEZ3HcTAK/G9R2nXok
r+As+IRErmiKlgTwKrdFZfFuNrai7JeFGN4YgPR8TfVRfeIr70RQmlSEYFRmHNoY
3SKqMCBCqu5sIkv/D8ky4f3IclCGyzduGYXRetLtANuePpGZfOnXedxwUCR3AApg
0hCeAmpMNr+tbVctXcqEKHSum4t5H79ijSZWJ23hFL2pAxM8lEDUUUwGr2B45Gft
nmxTlGwx7xBw1M/ozkcggcaShLnWNWUH4j2oDDzUMrn9s6yc0An/zGKIeCbbgQuE
Pkol0QgD00+dXaqBRFPsgnFzZAaTn+pqtnhSXGRG5NxGA4lgC6QRL1aIKDfzLxW2
MoBc++hJk7HcctUrDEBDFeyrCGKQsV5XMqKafeoRFFiQ+CIDtq+3IoF6oNTEb2Fg
B4Lqe1ub7ww5g80YRX8Ur3ThYnSDwm3ixZDhzsZMrFi668eK4EHGV8evTU1TocN5
YZHef/8DzpC2v3pGwCaKzBgU3uaXWODTlg9HIiHnKgTOBMZan6m9331SiS1OL7y8
veh2KuxmdINK64DummO1ditXwaiT5qA9gb7W/QOSViSO0Mj6NknBFMEIQxMnjLh+
QEpnFpbwS4inwXRsDtMubsikzjk0UeICOm+jFvT2nkFEz7cWBtmko3V06vasjqB1
Cp1aM0FSObTtw92XjGCdx5rXvc+8Q43Y1BCL57HIQAp07pq2lM5DEg/wjv5B1NX6
zkCD+jd8H4aEfNELYE7/70zAH744NIML8Ofac2FOxYkyFl7ndo9w+pRpRWKtnQlE
4Kb5Q3Du1ARmMdcH4rQbVqCyU2Uh+OJZKF3jRSdxGe3jf5kTZTlbXzalWdHd+jC1
OnkM5I8iCsPJUinXxnWgzl+FQpCQC4wyivpagK80VMP6q/n5uAtpjZzbrC+N25Tg
WpcX3Fy1R4ID8GRi6ylKx+cuME5KOJuyDMUB9RDZPe0RAjdTerNPYyAFrPwX4/7m
9tGVYcS6zpr34qhSV3u1Kutbr8c1sjajQ4U14RonXk/NaFBcHMnwy1ejSClCEici
8KGqASZ+18h0UOQQpdCAc5vjzWvQ2G9N0SNKYOKtAK6Mvk0HOQaKseRxDzUVlf+E
eKvM1gHjaSDS5CvyxmKUixp8ahMayNLjjQWSRyNxbaYsnkJUiYoUSSQl+mXGtRA6
79osqos+t6uuDy6nmtnNdfolokdfw4/ZjyRY0yPWItxrWQK+LRvJSu5n6ALcLDbb
TzbHw7wFTBEFG9/mtsZU5cUaKyCf36X/fUbnSQIXl/gQBwcOnjEFamALglYO5VOp
/qOrRcyjcIOCSGBh/9AoCOnjoq3k2xZMxfAOCA0AgscaRbhFx7kf8tc1+A/fcCO3
xI3r9riGS6jAGak1QAeDrOj9Sivb9WHztrB+gMmdJy09XkhkDqRv9fzjxSekL7Ao
t3cEf7sCy0NoNhGlvIv8j4SrG0RaSY3ObpalV90+abqHQhG5tXoXZSYS7H3AxcJ+
sN9Z3Qwm2MrVsWuxSLfx1MeEgW2C58TrM/6CPW9jbLYH5fp3Z9BXksoB3dkWvAPM
06oWdnoqQL9dpkDzH2rphjGgv8Q2Mx9WBoGKqJqGblUqeVENtuFmKwJFSCczzDkX
TeVQnYoPea9RgmBv+uETiRJ2rjTC4AnkrSGnI9EG9poAUeRXXFEfS6UJYpeAEp6A
jsllA6lkA+zXvI3wGuJN/2aI1gkd6/w7YyhT/2IGfiJksQEepVSTIv04hAmymeVg
+M48jUE0Gw+we5PqgtDydysriYWP8ORkWte2DLnQPXcpK2FPAPpTl4rYkMnqo9Bx
T29BON+Ysv4iZ2dhFpPWUw+itffT3q/QZwwFsXGNrJv2lBJ5aupI74b/i4vjspaY
ADWnpZdGZYrnVzRcrDg3ZTWtMu7SbGuCsLhtQvE1bRJAJHNCGU8CFOE64muqdgV3
aJf8Tty1iFfQsc+pqd1wpkrcHNIZNCeX5VLTx4qJ0vPJbHs+zi9QjYzXg+QD4Ds4
bKINjBg8HeYpP3ryVP1918/JU24VwJGquLy+DvGp62/njrQbuMKd1yyGb3KW2pRa
6Im+w37ght56jzVtOTmKt08zESFbGz54c0ugWAw/YvUB2CDSAlAC1gS8EeDUWKXV
x+/VLJvtAdUtpldSkw7aaFy8/SiDRlUEk9KIbHZNEivtRdposa2vNYi1bpKpLeRN
sl7upeFXyfMw7WC1cmHU5KaGY4+mn7v2lsV+/UDXKuDHH9qzmqnajQzA0L+z8yCw
Qu0MsCt70VPwcSVpL2o4o8/z/QESrRAlfCIOXPRPC7vj+l7chCBfm60Wgpq2EuLm
I7kdRMT2tHTqj/deI9QVQu417hFUi1nxl4ZwRcPwZ+v03HZXkjfq7zz3sG1ggfxA
U69emfv/WYpwa1DL6cvs3NinLmHEGNZQ8LEtc1MgFmzXCpMCiJ1pw7OhGMBsy7di
FJtRj9uubEd18FAbQYRgQL74QOXGHSpPcq3indKt9O28ONeLtVXSn63cHF9lwJTR
g356krhnxmwsZ3AnYiP+j5L3xys4HuOA1qdYQ1jxYRSCAgWS5yK3P7cMznwlTJOS
RaXlUzN5YsbdFnLjIQEIR4g5ldVnj55C8sqA4UsWKFzZ27tuTB/S0Ea/2S71nnw5
cvlbQ18+AC2QkKR/aBg7xmWgV5b/QMWnWR5quGn4RNgc1/Wf9FSwqgrrOKMW9zUb
lFXvTvdFyQpem8+NgP9tEKi9FvS5QMzKWWqWwTheubxMW8bXDMIWRu+PvcSFT9VW
U3NajS1c0PnHc8MmhINGCtRjL+Sukad5R3Z078OD4Qv+r/EMQu9PNXUbO4R21Vr4
36b7cxdy9zUE1ZIbxD3DQI6ieuK16ktRxYZ3X17vcXHLGZAuDnGsm6oLfq9aLjBN
7WpSh/wCVhL/nq/SPix0rK894whj3Ke3q7HmouEDdicpwkYXDNW55FDmTRnjHeMv
WrCZW4/DyvQcl4+IksqpYRDkVk2RjT5cU4+dJ0yKnxQTkjX+D1RnvcUIBBasZU4e
7NZviismRkvehQGRYyL7tYvOAMCCgKiziz9BKKBX6u5lEDiy6Cd316LLlpdtjC16
JCPP8kLXUwNN0s/y0oGcGWIm33H2fUxtum//ixO79gprcAoYvCsDClt50yWClcAL
5lA9ObtRfdPWinALeV9nU72gdpQDCU/oZjpOX6G1I6wQgrRfUR/RBff212ANAUB+
FikucXfWn3JAQ9wMY9SVB0w8B1rAQtW3/ZtjwPBW5si3zj6LNlm8wN7Vx2W1+6r+
w8JPSwG9kDMkcQAbn+zOC7dlKRAqwAfL0Qexlym1XBswPsI6nHW8qf5/pNm8rAg2
e8eqww49rZEuHa6dcou+ogxEENUjtfMASThzRqQ6rlE0yRK3jbHQEac0UWS94O/I
O7jwcKEs5wwxZzVWI/vkdCjgwwAVh1XluJB2hPgkHoSArhu/q+8b7ODEla2edmLk
tGF4h6feTB32u+7g55hjEPsMDNBM18FbwOHueH15rn6GMXXnXnxZSgZds3GXpRjZ
wfD1PACWMCk4T3Mmf+a75ZyqCXBGWFxM8+B4pPIQcmVV9pWRXg5w/EnrSjcwCbNm
6Iphe7lWax+A/uVF73IkJXt0RfXClwKSfVBU0iiHO73inULxk9q5AXuxtkabfafC
Ea7rG9Gv1YcoMGfYDN7eqvdDMg+1SzCAqSXBYZB/T+Lpl6/TPCPsdwaVa+HasdY9
XYC15SAcvPUhbHS2Erq4vSRiu7x0NJqT8RhrIJ4zqtN3oOxDl2aGeSySwyELY71B
ECayKNc4S+jwG9tdQ5DhUbxQNRLX6xb/20txtrPcGPyTOlbpeY13kbYVWI+N0BPx
R5FPNXcchw+757l8KcXLAYabRTgs65C+chWw0B5Lx3E3srDKlVMxiw+DGAFUKEUW
B+cZF9hF2Gfc0WBcJasy7PzQg+LQv0xz+tHFnqOZAFturq+1cygkelyD4b4TVA/S
n/4ImOzoCdMEoqn4LhXjBcbpg932TzP0hpvXp2qniUqf9mUdf52WF6tJjnTJXyMP
CunYHUqUpQPGrsbiAdB2e4y8FrHu2sXi9iUXvVlyeCAaljg757YdDA+WWnAikv9r
8r/tY0iDrt3t4/mbUOaqwR5YlVthBqPPo5sJkkscN1LVHkaYJ5zFZNHOITXDq4x1
xsC0W+/Nb+WqhqmtLEFXMAQ1mXbpFzuVNRPZctBLrrtbPtOnCUpX0NLVzt4E8lDX
b3hBY9+pQ2WFohveZM3iEvNaI4Kg5MvhjsuHM3uQtHjjhjLSe4bjQNFaLyVYCtK5
6445SdVvCzK8QG5P0gPLcp+5a1i89eMN/8iuQUEsTNjRN5xmemDcw/WZSuZEF6K1
8zl6PJOm3Xx3CISrhLRSvlGpDYfVkbxMXfcUf9SCPGbJd1GNSOA2sQfUjm/B7c8B
uDoZxzStkNqjtjGBP2AXvK1OH2VZpxfn/wlTYchRL2bC1maRRk5zMBQbuwPTT6kw
cwgIQibW7t0YsdV2T5BT6IlY8SZS9+OZHI0iJD0sw7OaI1Uore0TFjQ25J8rTTQh
R78Sqz4KGEmNmtVVdxU7xNMJjLXzdp+g8a8MVDyKUM9KkJqaXhdrAYOgEdhVmT68
IsN10cUqkwY63lVGbff4/qVpUNUaIGPEM8ocwqq5RoGEV2YpKA6bOySP4gGre0pz
CvFZPeH3K5PmXI4ctte1IMqsrSSEYeAyGmqC8Sy6QvPuZP4nYE0v+3ZNOfaVXVtu
4k6n+x0TSLTh2ZkHY15GOiRdH9zk0JHveCNe07j/f0RcgNHnlcE3b+Qb1CPpdRoZ
RNHqhX07R7UugA0MgsBj3Bz3xcs5PkQPq1gW4wB8vxWHkqAxzJhtCDOiaPN5Gdbu
qeVmUVcxeN1d8a27w7q4C5zrVGOtJOG4CYTpyUBU5esX+7WOwXTkR5zYrDR2m5HM
fduyV70oJioF6lnYQHxiVNnEy+WOHPmFCOF3Y8ZSZTgiunxRzxfMw1EN25eKCKWL
1rvcnFSlETFvLwuuTCplceGfnfsmnZflUre0PXW889oBmuRM/Y25AX/5nqJVI8hm
GFgE+OrxCCTN0sItEHmhnlgFMwG8uDpfamaonblnkVzIBwJwXETNlQt3VPcVQOq7
MFi6WoMhrzgUvFZWn1VhziGp7/JVbZ9forhVU/Op437+W0K4eZ0UZecdKeXyt1ek
QccpvPlgzAusadi1ONvMEzqhIS8j1FX61Mo2Rphs9i3R0HceFXwEwD3l7DncBdcF
Gan36G8WzZd1C4Mz86jEhS307kMsCIhZhX+MOgfmcyl7QHhlmzpbIARNW4c/5f2D
4yDSVKmiD7LNL2f7QxIElbCOHd/uM+CGL+apaKqF+ET/9gymmZUZe9zloIDU/3M6
Mh+f/hEsgodqarm0/k+j02/dJCp/ZiKQz6/uu91vPUMD8AKwRxFZKXucS2rMQJGW
T+GNoTh4Yp45D35DqgW32YB/kAOVzC725VUCKXPXV8GY+srl/m57PMhOK+iu8jsy
RextiB+p5D1EPuUXkj+WyUMmxLNXngMER2iUM4Q/LR/EpJiZ5udhNnDvAn7882Xn
9JVixbm2ewc7DK35sPSdQhcWo4vXo8U1AKLltwLxCnxDKz9Sf2gb8RUmO0Cd8DA1
wONxgT+Nvcy+CNSi/owbOCB1CIEUEC6TW7hBZZ78LXwTEmdhKpI5VF5UmChEKoFo
ozYPM/Pc2TvFN23Vv5MO2E7V/Dk0Vps9OSdYAgHgg7q+7YbRrOcIDxF3iZluo9EI
YM7W2IsE0GPz+SuO7rJoDAsfYQ17tpVt5oDZan4Ex6S+kRur/wXGVvAGJjsfmEJ/
eZONJnnjAR2Bakkrt3vPH40ov0ZFeCDUUkAFlsp2HSnm9oZpkPRPQuQkuF1VKoz4
Tm9hmfIsSanCzMRPs0GnMVFFy6kFJ/GZsF4JNDOyRuSgFt9nddVTVQu7f2Jk+42+
Fo2u7DVY0m1NrOlaWtFVYFU4cO3a6D659hse4wKSR/sWN82cYAzvk9kWMu3W1kad
KmK126ZWcjsdY169nHj7d+gLsF29ucZVEtkzvtiovEdWmh6++HE2XVRI8tYDx3kb
2tzMOChhFRzmvMpcKhW6sp6I9xvbOzfyoPeurHnzAKKWjLRWkCaD67WT8MsZY8cV
5nx90ZBQMM0W0V4bQ291c/6N0Oj3nR0NgxXXxTm4tslpbWRfq6PwGiftgqnScrh8
pRg1cVEuuOIbvfgtBq5vHZjKdh05SqBDGL4wXF1EAeJ7iwnMcKu+EkHTIIWNmRz6
8NVW/qOx2PGK42hsJ1bb4GOvWjYlOTvQ+ZICYjuYfnT1hFCfBIQSNHU5yo4sTAVg
w4eUZ7tszcZ4cFG+iHEul6bDQBvt+lORci17TvL9mNQj9Th2AVcmStCbyG1mycXv
muRIdxWW9SKBPUS9tCk5mJ5SJUINqF/F9b7AbGUE36LGVmxYLad1yLhhsmbXgQjO
lwnVQqlf+qKfUXEH/km/SmsUnZgYgtV6CjWLfKhggUsCecpTuvEJAS5EBMEUz7Xi
BcPRDwkkqm1HklvIWMo2XUmvQoJTiQ/n6+7r97rBAFDTskZsilH4t+W5aMjl5EAJ
NZysUMfMlrEUpBoTZSvnCIG+Yo+5/WWwRCbwXhObUl8jkywtOEZZ7lrtSZK9kP2L
iAXZJxzdCTL0GcDURd/xNaOcM4FQJZU1DrerhLctNbUZXQnjKvaNlXkQpcMpvuhk
qaJ8Bg4kW/WKb4+8/wRaByQLoAccs8gZLHZhH1buHgQKv2zUASKANE4XLrcJZgGY
cyKbOY0/01DR/ZibcjpPT1wbNRKGVNfXjviFTfCrYj5WaMuasz5FD5F5fJprWZXX
DYEgadc+AAp7swquWMHdnxP/8hNBVELmuO0Kh5Xx6/uGQqaclo8xSxy0YFkUIvpd
y/I+42UBVOHk5aJR2GE/a+ASvvFJ0ZNG6wsh3hxQ+vOyaJgMkoSmoZn/KMf6tZYb
QHn8ThtC8qcs5gcAW6ea6Hy85iMrKtvXLVcr3ZVhDPpmeVC8nhj6uqRy4Q8+qXQs
+PkgHV+sSJyX6CrPvhz7qaYcAEpKkZIt6TJzU7HVAjIUA215OJ3BFmcoMvcwWuc+
Fk0blXs4gd+c4JZ+2hQtEEWUtJl+WAakfdnbjur6EFfDlUdpGTF9bcmqGiWyCL6Z
ApJpSY3nv9pjkBy5c0uiF4SPGKH2jYZLUS1CFY50BpHtQnl+LCzB3wc9NjaLfbd+
qR/3Wv2kPOE9k5uSFvIIDc16guw0Hyw5tPuA/d6tIlKI/fkOs8eAURrknMfU5AJ/
GUFWSDrxz3YeFjbQB5Oy0cgUWhtUkv6Tm26nhPUSMGTjKY5b6Rb+o0GE+Edr4+Wu
xEdf3P/J5wOM/Mi6ZcpoHnb5Jz3bRaGYQhsvVzM3UUeW3Qyf3/9aAkmqej0pzntF
pJqYtf4j0uyuq8LB9Ai5VDYKQ/aoYiLuXAY74e6y9/1bWDxSJMedah6RvoLctFva
f9hLDC9s5EbDHFxIOt1yAdH99Ug5BfOpdzbyWQGbxI/U3XBJpcrsRR5z0wqoLdK6
B31RdoawB6f8YCWnxfxYnnkafxOuaxNmpOFTzOEeCqjWUMprco6MaTSQihB3mf5A
Z57ieBvRl6+Z8824z5URt0/22+qsMKsgB6HlH13ho6urBWzY9MYzcvmnJYIBMNkb
5zvtG56vI0iQ+eEGUWhpCeL3FWThodd1X409FXlXZgOPh+G8IkRy/VfBL1Gp4HB1
rfKcKDcKtgbortCqGvUxvpFMOdKBa84QDrsX6XmG0p0yhLe3VbDuhckxQs3eOR7z
+Q7Nt3dGXJzJz51axUA/AdM4UHyZnDutD8Oo1Bm/gFuR5xYtziEfcvjPgEhagSnE
sm3JFayXo5BRzAMTod8r+/7EXnRGSt31X3E9Y5Od4IL/2OYu1iLH0msREDLTHU9k
2+BXuW15jBxgQOtkArj82aHh7aqm2v9K1BE+6Rli0RAvkgoueGD17nVcBChKW9x2
wGtRDosSs90xhmivrjYa9RxaVo9Moqf44nm7rc3El49njRzldC5mIPzDQDNL42YO
6v/L9E0dnQqF620zq0DqEIusa+v4Se+OmVODAKzgxZVriV+GWglMnlFAW8Af+7D3
14JC6guPb1/wS0qdMZUUrDMQm2atr1tLZedzXT8Wcz+jMrsCkDsbA0N5KK1Ejm6p
m79f3XWAa2KUEudMhMKX/dmaafYvYIG/h80GHv366o/KdwcJmzLMQQ6sP9JIfBNC
Y36fVKWAHQDEKLuuClQJYGqO1kUk/PDKFOQh8TaWxOOqVrLk1FmkupIFNlrLDu6v
F8AeXBIoTkmwokOdSyFWx2fQsaJSlJnKZ0une1ppdLZL5aKkUr5blZa4mTF4cDh9
e4PKFDqMPA4CuTzyw2mXBldz3nwxAx1EHYgytuzP13OY35IPpcB9kAESmJIPtEGe
iRD9/KMQ5pkpMahWJAjAkuNVO8zD49T99EOLPbcFkZlNRA1lvuJVwYDzkyjkneYp
etT5yAG05bj/j0NdMZxylCYwjr8cGOQYIpnpNMBR/uZWstEIfZjRD5zP4Oc7P/KS
h8jCx6Qn5DvwiObs5zRkRqgnPFjalcbjdPnChjUr1i/g7XGpkTW7LXoD3wdYMwhr
TAzuZvJVvh0pm9G7jrhnJoMza/rnvIWAY2iEgTyW4E/OmDJOscOaROvZ7ZreECsq
h7w1oobTa0Lb9I4ocGQWVwtrvDO97Mn8QILhUQvOm1ibGRf+fZE0n2NChTPoIHw6
XqdS76peNHGQSh3nmRaJDVoL7N6OcdiWkYCC9evMeQuE/XtfXnV8eDlW56I4Ns9D
+YRQPbypnMqVpyF2SSWYaKqc2hQnP6dr87XuI39Px1W94TWoGSGOp1IYPqGF0z5m
TrhRGSoNCh4t1YnzX6AO3uhiEydc+5USgy8MX8blAmM80lmsf28kNClGnEO4bIG/
s2p0FW3ZSnr7snIYuDrb/IJ+DIxAYSJh8ek6InsosJ29YzHbXHaPizCdC83BNcgV
i1NbQD5ljNuzpWdyvkb9ZdVkC6CJxURt1cCa7IYDMNDZ1CzPr8fuk1yw88BmtbqP
LEvafgrk2NBazY3MHroadtJWWBCpafr/IdOEyO1MrweghSoi7JG0ob99uEobbp/O
e6zer34afBQvz02z/Y8Q3jp+goK8FEf6+OSthZaZiVlZNwMRdO0b347uFg1C9IaI
CD0vmpOyfbEmNm/H6X6IA8SldalBaj3LfqU2EhM8yMFqqRaHK+ykhJS2aRrbS0vA
n+C0kjdhKSSmcpZDKNrr3zmHqYr1ov2CEmHo6ITFc9+9d1+KyNnabvxnDIkBsJek
3voY6tDbItb9ZluzImKrJszjxKBE+0HbRlVcaAiQYbkhpgu2hhEs6JUq8aP3EyKV
f5+HoubXbcsJXgw/95rig/hmmZyj8GqdNvR/T/ncLYxZD5njyHgjx5IqjageDjX9
0vbokqQ/hKOc3qZA4Cm/IWv2W+XVWVpZq8Rm54QNAi/5s/3z251MDL36nlFx/XGX
kD6mrfzq/VJ3dvUNUgce8kw7V301j36zB8ar+c7NVNCLwMqaDY8ZCNMucD3WOx7V
WAemuahJ7vcusiKuhKv8VP0MCvTA6IDKLHwBUdCbH2x4hHXMh05ZK/XTldeVf7aB
khyVvmA+haRbIc6UpyGU4ZAzv+nWDnn7Lj/4ftC/sQMJ3f06QtTplPwZQt/pXGPB
YY+QKNaNPtwhAB7aMVboRR5RPGf9Ngh8RSP8oCZ/37oi3ProFQ4MBu443T6LSfNO
eP6ah2COFAmdDMgS3YSMBerzuh0AStHTHRUFHt0ag41RNhDGWSGaNNi2mQmaN++h
R9dCjmOm6MLc7JYPVvpWm/K/VF/id2K7s58OZxgmjE3dXQLEFR2pTMaFOrrxonBU
GBNirfR3YkWG7PwfYutYilsDz3+6n/gESd+fHgFx0VnnjIE8RY0yJ62KOR9QVYUL
OB+B8zI54m4NZoVtzkKNHh5Y15/DlZWkKvNVfxig59A6kBFYEYCDNgW3Ha1IDPzn
TbUBvCmfELOdMzmd88JFTcFX0/JSn5RvyY8WfuRUifZ0YYZKxt70ee6YEi7W6K8R
YW56+gQFp/oy2WgWsm+36ymuDvbBpvSh7P/nBlN6VITyymtENmIBhs67Hth6tdUv
g0mheyb6b7cj30LaKDrQitkvVpXPX0kNPWF9EqwmPaXI0PDTxDcDYjVxkNN+lBXy
dj/zPNiy48Xb3ZTYIxY89PpFFQt369WfsJoprNTNpPR2ifmo5imyFXogm1eFRyGI
NOXLJ5YojtDG38axBA7TQNMWnxwoZZfDTEHMXMXlCa+bsQy5VC6swReRcCJ+siUB
Na1m2dA2ozq0nntw23hxPrk3bYbMHk8Hyi4BtHRhDQ98e+FuVxIHu6+IZHdXXuDm
ZG0sM6/wq1f1HsaBtrTnRG2Qw6tGdheMnlLRI5MXMTiZ4onaRymlgNhDm8HD2RXd
c3Idswd9h2D3SMjMne5DwY6KmM4qk1SPHPQ0nDmsD2x3lgIH2cMLEmBZ2IAm6oJO
0FPfkCdOcmm8fvoiAjHGvLF4w22uM1KQbJ57zO0UUTFMpzn9CTA/NXsPP/FDWQ3v
yZW/vHQHMnykLEchPc1LWvPhLoi7M+0Pg5NASeMaeqdTgs9ZFp53CDojV+jSruiV
t/quJh2eUbjUDDV43yzugkUuV+TijknxfRJi5ZP1Rydxbk3tcNswOQk/+QW+1Uaw
T7q0KdDFGXFewYHL+VLZN08wLTzM/H4Q4efTIV6DUk5fxIJ/B1nFYkwJlMvwodkM
YktjoBaic04gFhRYnTbum55Bfi+Wqg4BCgyjkwhUIVEDM/ZWMQPuKwM2OP4d0Eed
j4AA7JR3H0b7Y1cE6t/Kq4wRgZtBMWWs/HcNw9r+1BYt1nKf7u1Jp9biAS6cI9CV
mnkg0EsdDoF88Il/m3nBK0uoxTLXOTsALBw9af3a8xtsrXkrqnqZ6E1PvjpMCay/
gc36Mya1GUpl67yAztzBxtdDj/RHUYyUgnu5bDmocmMzGakBIJAfNP0pMNz5JSTj
cAwdcOHJ+Co1aPgCRlKjtO0KergyQox/xnBwd6ByEv7qso3Q31O9SjNTEMq7T5jX
xKFibjU2HeslDhX5wGKv25Slq9jiYiBIJtSe8lP3Jdvo/Jq4tfOiFjdiRKRFM0Ka
ls3FLKR8h5Vtzf065AY/beIXEzm/VeJ/CS0IaXiBGwz8vsDJSrEytnkYVJqa3+jK
z3QfAIDGUSxwT1/OOgqlsYuqup4EUW2Qc2hnyAi+saie2P++vhg+rXAFiuCoiyYE
zMA9T2h4jALOU6B5NoCbdTCFdnV+3iYIWOhDW5IRWyRGMNgvHANyYA4o6l7PCUMt
0GfeFH42D7ZYZi6NDqnAuP543lvlblYvVMLSs0Ok2x4xi8csebxqJRtq7CYypMpX
YDWtXYAbA8kIwz1tI5mm4FVek4Qjvxnz1IUEZpGdhJcW4LN7bXH7sNaXBsSGTLGu
xqwyvQaMzz3HsAgOaw5/Gf48eas37RYaBn97HIakOhoFX6gOpnoU/7JQDA3ko2YQ
c6u4bma6xnGdXbofUE8p5kihbLDdrEwYQYpu7EaZO7tKAcB4mWSdr/yTp9iXsMnw
XCoL/PciUWQv4MZgRmbaksIkZl2DSiX6qehjl5ivIKxaUwg2tB2ne8VaFAAqytqm
ZonhutQqKL/Q1YT+25HiCGdXPWvZjPL+rfwWpYmFuL3ahK/ptngf9Wp8OO1m7+jg
dLYJn2epbzvDsEJtY89UenN5Qb0itDDvt1J5wLCF59vo6rlsEU34RINUcV4CTSxc
LtJGcasZxoc+356tm1eg68DgCM6kdUpfpd3kNbBtNH21y05NZFhlyt0J1ErmIFqR
Haqiuqgn9r2AwZjaGxqy89Ixhr2S9uyGEGx57MKym82Rr+YBIezQBk0gO6Mkd3e7
CTF2oKrfBgQQgHL378WzlJ1EuLxIaEM1lQPD2EzI57a3VrAZHZ7Sh7DSewFkBYOp
+L4KdFMMMc+6TGa+cIJbHh7zq5IaWS2/v7gB2haDoHliBQUR7WQRCHY9O+MF5u8K
BjByZxgdIG3fpB/yVVxvnPDe9/31716YDrCrkX6hoIofePF+UzSh/+/9z8abF1H7
rl41miTc/O/+761Op3AEiacfeqbczOlXO2LY2CUXmJEy0c7qvwcqW7Ygt/1tmAR7
QXLxGekmcN7B1BcouXihMN9rAOMz5YbbsKQNBfNzfFraWSGHF6WAEfyGRRxldrgQ
uAJbp3BGHUXL3Ksv2tcOPDqOL7poi3GdjmZcMlhKZm4yWNJlLpQNXjLTzYxgaLwf
bbmy8bKoiwbHD3OvUN+4Nn/e8eYcjgOUwRRDPwxONgDulypJj9wSsck8x1ItZpBE
MrO09kKeTj+3v85aBp0X5jLjRYHQlJkvFHd0Au53KZqotnzbmSCbgpom5zK9uUQe
j1jIuBTd2IJcuVamTXt1yxTWNwRxz1Y8psK4u/d0nXIE0L1IHTb3b1P9gGu9KT4G
jXrOO0BmDRVHKREpcR+3K89n0K7S2i0CyMzRZ9XMIX7ABbdEZYHln+xOLTtwsjfK
fZEfSiATdaZ2hcT7dCgOdrsh35zB5qJ78grv9UV5E3qcoUvHSfPxdBSwSGvXeK2w
jllf6aW4I/2Mc5Y/xB7AFAnRLqPk6j+jKDIsyhL7OvklBvjXfk2n3dZZrXzMnbrr
kc5PtwCNH8czsuvleeQommd+OGjuA/A+Ogs/+wsAGjVrRUrnx5neHZzXqeoe89Ne
poMaTsOHnfJmRFVV7VemNVNgbmfXe8BZMezw2nETLKUKfN/Yi8VSANqNIYkxqUJF
8vQF3uF53OhVb3lc7J+VR+/HRcO3JB2DZma9U3QUjW3IcbyFyRq2xkgShUWzEYdH
1abP9acQzqzYxufi8+gtT68qke6Iza6jFNEBWd1TQSmDlREJam5j2dNJXl5DCY/n
J759omC8CSlqp7anf8hMDiMPXi8Ut+bX1LesIQnQLGuZI9F+sm+b1/ECiY4/0Ehw
xGLwjKsvMjzWgsw7T2QwP5gyG3rpysLGqLvccWzzjF9j3hxfbHKMGGh1POrvBvNe
j6plV+5gh7QMfr5RzylDIqCMLRpgY+unFu8h5oRszKr2tQ5DFuhAoOrWbFwJDHJ4
917WSqjgWnsickcbw10sl96189zwaIZyvljYwGkWmw7R3sFL3fxYH6Y0CALwlLmU
KmOh9DIV9xt42S+g56wm2nWek/5mr/eby0Mo3fQhTrx0LI6Gpu84OQ6qZK5ETK1H
nzcjatQXeRkW20wFGbWv4UNQ+WzY18zlmB2Lccp6EFgX/LMZE+7jnaDW7a1Qisbp
8ZAWcbHHm8xQ7TnXNt1dTH5zGK7qgfEXyLSzIH3uiYTQKoog/3t37+RUlDnBu7fY
y/T6H3ZJzFknXXOo8a3bBW5yI0D8rkTXDzOSx5meSnZNmH4YNiTBWsdDyOf3ztji
6oVVCtiEJpndAr93UnYEVL3XXQx0Qf7ywrOMTncVgN/9EJHmFW/dcwugvQfAEi85
22ISY9fJ8xNAALIffIKvr7e2Rm5b1G7+e6DPXigV2NuydeNxce1mYJTnQGEA1vHU
+qQpRdge6CehBZdrvxdxfGB5y6JCf7rE2wU2bqB/2snxpnZ5Vjbm4wM+ziScq15W
d8ccqpcMNi0yY/KWpBo/Tv7bQ3tnBVfFfpA+TLzC9epLnw2kqadxlluKzKubtoBG
1KYtoWVxYoQZpg39PSJ2drN2s1HkIOKPj8L75cWuz64kx30BnEMkeBtpYcBqkjhP
fGu0764lNRnDsE2tL9i1jsjVeKya3qXDZnaxy+bjpO1aXPwRahwCQSOpzkCqbl2W
XfmMbCpHGBtrhxDD/+xfGYp8fCv5nemtTEZZ7kAQw06c9nMO5lw7gKZTPXbANMVI
g8X8tE8B6GoKN5U8xZ6f5SNAuXdWlSREvFsavqkADQ55ZzrPBAqbvJol0Y1ivIed
L/T2Gnf2Wc4zWaDsktHWrinoeGhhiY/zeWB/1Xubm+HqLUFLlfR+64HDn8rvkvWi
Fgh7GH60xRinEFwIIo3XNb7kHpuisk3g9jtPC/JUKA6oyDYqlyIFuvfQoaXQDnF9
95+VWsazMFn8WzKEL4FoXgQLfNeULjd80YcBj77+EtphE+51+4yHdRWrLRHV75p2
LO+LveypECrJ7r14KmF+OYM0BSitKVPxO27WVnoVo1Chtudb75THrgof9iG5nbF+
sQ/TP8ppYNncEjPvJgXIAxbhjFpo9/yLKvsICXzNORDbMarj+Czcz5SXpB6I3yTJ
HQw+TAEtACF7z2LrlyrRUFi9/uYZIAy3YpqxwFfoADr40VhJ1Fkf1BD+lEn/7+vq
0RFPDML/xYUywplI+qrjszivFBQo3i97rnIp+PEfafWvVLp+u6EWRhjpRzXw6fdI
/ytYcAWhP+WN4XwgpPUerVV1fei33B/jhuN49GZ6moxOhm5O/Zxj+YIXZO6WSswe
Q5xbY/7Faxbgso8LPqgTi1LcL6GTc/jmdtAultmAnfzlK1zfJAunrYXPEzNaPnEH
9PVdiHiyJxN2oDXsVFnQNk3SPkfnwo4DHwdKzxkilNB7HDBpnLwiNYETaz1yBzd5
sAvAEmzSNnmlFaY2n/JvlNTtrF4eMolIZMcAKBqtArDEGHGYwvBQgDpE/Z59atCi
YlyfxA81vRVsCXGLzG20R4iujH+3zP/kTFcpwC6fltOfJ8H7jhlKlRMD2dZE7g8Z
IcbmdoC8r+0cGlcXxFdh5xAZ0VD+shaSMl8L9uoVQsogaLuQKLa1VfwcrX2hmIi4
sP/XrvdcFnm4/nUpCUfsPFXrdenHuPtiE7nxyEgE9J+ohztl8wRLKKeTUXhDZte1
IV3nRWKmNCQitFxroN6BhSMne9wIHEnrPXZXZAudzkLeBfuQYWtGbANW03ExokGK
xHZJEsPbDj3gKIe19XDwcdEmS5/xCkqAuZeZb8zU0ptO008uSNnTkdpc8pzHWTMF
QsjEHLaN8KM4aUOwmZ1aJnWxnjbqvjRqSx/eAGWG39zDJMH7uQnBSGr+S3RebcY/
CfGMPdp57XAGxww+lGDMiLT7LLjps/6yeSU0rmoLPrKWYkw6MYaLY4t1KcZ85ntF
xGvDoSaNTubeIsWgelbehRJf34ELpa1JXJASpbq+WuaHW+ITniPlDPlUxJA283FH
ziWhTPdS0ZzvGdhzaeiuW8YCVh14BaQEZTcbWv67lTsNguVlTPdJvoxx4uzi3eOa
1CrvqzeqglQhBEcSteKlkxX5uwvQkOAN/vUPcW8/CGJKvZStBo06IoFKW7SrLeYb
ZwmegNSE9o1RNH/ikl6ItRFomgoGmFjx7DELmVMwtsumIJue1R7K2NQ1G0jswDrW
gOWAuWbVeiXhNvmSytFl/LHgbwX+8tR7fqRr+ZjLZB/wf9NBAl6bBTuiHHzJAEu/
pPdNahnAB5Fsk6Q9DuYuqwm3Ixdp2q9+C1J4kVV+T8o8Z9vw3K079ln4ZJ/iXfzG
wfMyqueNyMIjvEJofxu+bHfj2ZwzZb9g1Fu2t98PlRNVq8jjiwGL6g+vFYPvyG2I
lMRsz8SZVwOZNXNeHHKjrBhOKPadi3KZZ4cVIBr9avOhZqw+gqALZMIq60DniS01
EWroZI1XpFtwmQqS63x2tgFad1DYfE8hhpytOXYp/bggPJLSBShngeN4m0eq8H5F
yiysRYrQP41iBhpwuyvfk+diIkkvGdb0yzl1nPyICCWO+w4xCoIdu9Lz0Gu5AI+2
dIIXDRzJ3ncB7AIJ8+eYrsrm5iw6Kpa52IpAKCVM6spM7ErEjk3B1fG5F+RqtnSX
p+RaJwbbFoQlhg1Q3bp3EG2VlhDKXFgJUGVAXaQCmfFfq/k+dn52bd5dUz/VylMC
3qauVdHuL0Y6fW42pzqC6//948C+nJXZtypWBI2MQjszjXiBrYWrQUKbRS2uVlIT
1x4GXO67ZepiYS3y7bHwucnyndBYR5k70VNk56bHKPdSwpMqA1ZU6Jr7GMCjnzWb
PJBvk0RRTNx/CNxd/m/2LEafzLC264eVgVgYfk9h1zaQJqOELazdctOLlGuRP0fA
PBBgsxmOJtbM3xEsIMSrvDjPlBonIo/rBFrdBVciigwNvXxNXtqHMFiePs5EQJ4a
IGOo8raR3WgnfN4loOkG9mzx6DIwzQJzXb+H2rKn7hTSoejD0dVplJpnBlD35hnd
dPUy7u7sIamNYfZP/hD+oJUfSt74dK+j+96Fk5OTLEjiow+MBwXpP2Y90R9UstjF
tRi5oLkIfEM1ofcICn0xnPKvHOjCjU2gmD4OTbZJaeT3CBFnagvKrzjOsi8CW8h6
y0kla83UTXmxzdd9WveRNylPziR/ZMeV8HrhEnJUOtZYRYRhFb8pGozY4GzlTIJa
xSe/E9bQIhH9AZyyAm3rZnv8yaofnB6m4335XbHgNrFnJr/TTtS7zTpwrc91EQ4E
3nxfKWN8QTMZE+EMCR8LmeE2SkS8CQVeiwgaSxLWhOtNfZ5+yap+MOTOcEn/vPf7
qSmFZkENHzL3Osb8h1QcY69OKo//cL1sVmKrwKIL9zA6XSEhoEnRs6eppb7GeJFy
TFuekzZ3q5d8EWh8VuynuTypBiLu/6PEYyP3gLk41NfRhC9bJTPHTR5YB07r1oYv
IaGgCuq4FW0Tjh/YnlDxpCvREiQGowHQe07MlLDgUWtPxltbXsyV51A8444KqHd9
OGSG/w5l5SB9c2Kr7nm7khy1mv8lfwNS7n/RwWdXLxdc+ZqZOQVTXeC6i5bydgHR
HaNpkcu+VmJpyc0+xjLhuBFC/eHGBxEZVlX4XidoCOwHjKtNArO0hb0YRsynzSFe
j6NXBCOnaXt2eMeEko+IVUOc4zzcEcdZJzYoWiKPljZfIyUuaVa+aIEIkw9fAu7x
v5OFDEBMBlsub76vepo3+V/0cjAHbel///oIKoj5T/H3R6XaGfa3x2l28EPKBCpV
QCTEKTzVp/l5MMuxYrhhVnTV+GSH0aBChe8AbWbsBfPsEr1LWNkVTU21a92RV3Fh
3WQJjpq/2HgWLcTnO69QH6GUz+LFhbi0eP/LOVibqiUFQaebiJ958anCZKUxYAeN
5pDAiYDEOOTw2cWH9md9tHlkkAbTyPYx6Vy55H/jHv6lfSSvHPVO8op1xc3LShNO
p6UYRW9xx8Cup9ckdwsEQX4+vPtOrP3NjtNlqv9b4DlbD9ZPS2yG16+urnGgwO55
wpYU6uF9hWniHfrptcP6zLWU/w2bZbkvPM6fYfmWBm1AWegdgKLcfgZE3CMFdRxH
CkChkaoYwf7YsDRTDWR8ZDksFqc+ahTqKeG5UpfsPDvWSnIjXWmfaEmnPl7GfQdY
qjwm0dRT49I/aSpnOEankII0q/6DYnHqdbwfuR/dBCn4qodznlLMb9nKl0XC+CjT
s4J/+/nB5SjYRQeiwpX88Qj5b/Qg1hQljB0f9AvzYtcru7YN+m42JziZ0oF6w5z8
glKzp+88FvqyZ/3M9bfde1BGH2ZzI7lveKsk0e/66qSW53zYn5tlip2QB7s/AVAx
uDgL5DgTHDsy5hgqB5E4/WYzCokNEzOC+JNqmTFbmttfYHfBGuaYmBMMMfVSFIJe
fb1Hfw4OVQvYnnOBuUCtgyM5ZV83GoEHPrx/+vxg+Mp/9UzgYq39U9aTPCgp9lFT
drx8g3SPv48oKeMcbeA9+TAG68rEmoBvVjLHvDrQOj3Cs1fLb01I+W4MVzahd8PE
e1n0pqEszj5AOFwTPG0InMMHBSsA3lst/LSMJ+h/3ZSXhZvEjPzX8jzTZbaBufPu
Lbe+ajfVCIYwL6yhtay/7V0523yB2NrRIaG9ZozrWK+ybpmuOwcM3X3VsBkMBZnz
u0cCmZVEQdM3Ldo73ntQ0Y6oFGwY+8Q2oodzwzPMTCnTA3FcMezGsN2m3ghujsNL
uisWpz+IDwOeoZjkTx8lEFfzPK0exWnAfabUZ7BY5NncIRi4uTOKnQQhGqcjFTIg
yJN6YZ/NpsDUjES3pXAa/xrqC/PHXYIgpNO2AsOl3Wo3m9W0oxzWhxkKaFqGeZmO
Rrz1ISD9RMjfvKL5pv8Yble9h53E898pq0vA55N5qch1jnhuuqkp1rgsJK3Cz9eB
UtcojjVObSSguypGwxDn05L68m1e7tGK/O11WsR2JAUKtFjhxC6RC9hSlwabiEEH
lBHkbyJTU3CcKO/GYNBlMF0k2lhKDt87B08GVnmUwhH/aU3mycZpug+rvXc9hej5
Eav9FJd0LOSiQsR7qkikRcPSw5tiSscvTOypfUAontb/uXpLCZTW1DFhJWreyWos
miCT2rJpwsUsd4mFOMnqCkgz0iKVQpW/2T3CnPW9tqPaZjytNQyJ4hJcWhzafwul
ySUvstKDzTkB8tIuncq0IyKqXeo/rdU74l75PpeFZ/wTnu/6Qg7P+fmjKd1X8cRF
n+DoxtxVIIXaJDhhR6Ad5Uey3J5FVylhBje47C4a+LVeUKSPtwdUvIKB5F1H0Qwl
8+3UqIi6/E8xLUV1iZHZbLbF+ouqC28g4jmpZe27oezh1J7QtaQW2OfKkJoGZXE1
g02YjHmi3DLOwu73a3DrwwCFmPFH5TtfrOoCGmL2HLeyU+QoT8qQzNPC5/zLR3Tb
TOt5VN4DdUT0NUx1iFXJ78FgwUn5LQoxmyNIdjZP/sFA+Mf58epV767qqfBy32Bf
tvEixy7RKOxfQbda5gPSqKsxaQD2AE4up/PpQ3yNDC2ZrB9uEwPDT9qMxmZLZz6c
Pg+pquCAXGRXgBOAZxrMtBS+e0f1SqA7RGjXnt1ZDmzT15kVSH95LJV1RFKQBkK3
qwrdeBOSSNQZbAi/0pNKAMG0WlJAXpiW4Bx4qFP84rg7DoIm/izh7TbBVrCMx32x
tF4S0j2uN++K0JLVje0nsnoBmmKWTQLiqUxEDwcUtEUQ2zs/Te5H18O9gxtLhAJi
gX8V+IOknlUUSAbbDyKcbouPqRMgyzb20GFw6ed08hM1VSOhE7PV8KvPztMAewfk
9ZnrT/k+5rjAhvv7Uoj8QJ/jWs0MI1gxy1avjPnhT0ivdBi3DaEtVIrYxOer35tH
V3eeRuF4sUrp1b5zCU25/65YX3auFTBG7rDmdtxo6AkK3MShhZwQa1YiVvSYDUY4
L4JlOaQjHE4npsUWfmlVWifRZY8sbOz1J5qSyks0dbtjSU343H1/OmWd/ITJi2qD
bf1dvomNlOKzByw3653v/lF2jNBWtq5OZUfRSSNMl8xLZA/EHznLpnEyIESjdFsH
EJILdqg76rsofoXe+PfrExY0nPANL3rI3YXDVyA9yyxyiTB7kHv93gGYZca9vxgY
HDJCoKpZW/9fZVjlN4F8FVA8+WfQecsa6AGNacbIb7KWjRtCh47z+0m10MNF0ug6
Jh55dLa5qe7mz7esPj9PYT6/k5USlT5GotHMxspW6bkXjf3Q2O83Lxr2Ewz4G8hw
Wq+sBQC62OFK63flqrhOpfqrwa8GYr+LLi4W/YglgZvTkWIGdB0uH2IIDVqBhlvL
KgdRl3gnrncj/q/ezvO3NJf2opHHbZz2kw3Sue6engapcIzD9YKeQmgNCv9NlVuN
aFnzIi0fQBelJ0MIYPvnL80E5i1UgVwVoFAWViEumJijAG7mng4kL1NQcwVXqO9A
vnzbfResBuSEjNxZQRPqN70vsOPx1DQ45mMe2p6lAKqKQN6bySQ+fWcDF5w+8d/T
AFkd3E/EZusp06GaJ3JKvsd9cBiHamobNIg3q0MCDrJNGR8tyq4DVGI44n4+3MNC
KhAxKZjpSq2jjIR/nCCEm80pVJOfvT9wXTg8hs1yyoBR6tb9GcsXWVP5Q02TP29Y
nNG5ursSSbc/kMya4MkdnZpdqe5eHUgeigBzqP/9kqFhHi0q69tI0+5zYDHljiio
t4yQmkpSsouuVQmCNfv6b7FW4KJwvLWa+0BKglF+PNKb4ow4PHyNep03RhdUaF5K
gOZfknxzVyOodJufOQmnNYvhub3hToMoIRGtRwi6l2+lTVcyF/DIQtUKD4N6VYui
zWJxd6LHIyakIe0OlngChjbg/6BZ8q+OrM/nOrF11WiOLueeJWryX1RDzpIf5qLN
dG8yUvN8WxP5ymq9Q0hA1l13GiPxdbzCQfUtTXo9qat7qd9lyIKMRLcx0tN5OmTQ
dXN1NUkbgV2nkJmMNo+M4NqYoiwm/+5XaevzrqSKiWjfegoM2/Y31dBWLhU2H1bq
luL7rlsRh+TX/b7g8kH7s93rXVs2GboTJsTOLYDWVp3s1xTL74EpElwlcnyadk8M
g32lY0F5gUsle+fXXEmZLzSQNupdoYy/WPFiWgSTKJ3kAGpCYwq0VvwNUf1Fpgua
OjBEhFRXTZJZ6R+DqD/ZL872NftkkCfhya5zCEz1fLHMfk4qioKCPDFDK978A7ac
TNP8SkyduR92X8/1Yq1YXtQdw+wfDAbqP6FNlf6uof9fCKAdyMb9uHcrfqtBvCmD
s6L7AWrGvc2vCtEcy+qdKViI27gXMjPHoTOmWmZsnxn1qXQDH4Ep3OlfAKgOvRH1
bJ16JJlARWTQSlprnGIjpNsUvLkRkG7aoBLos4yfHAVmo1bnZ00JHsL24MSFy3HX
z+8rk2Ke5QcefwgllUCvCYs98ffzsAOC0hEpQKPcBgopXwCZxbpGkjSPPCIhGQqD
eIyHueRNeRGGR9OzFjYEYSkx88lBFpHHT0Vtsur006ePai9yS1FfT4zfIW7ncRH4
4EjGxt0ojA6uSyN1+RYhKEsrQawPR7iUNxzqWsQ0zcfo3kFEkhmpbSEYGt1TO7lX
Fxt/dOWuXquoWJaveDJahJL2OWd1uTDJpOpnTPx5PT/dfWgXMl4tOF+TJDeOvtpC
931h/MNT6i7Za9RHRrRyPjUpPh0HlTvzkYfL0FSfZblCCWIL490E6nFseDasqFjZ
PaZJYDamSZYB03XhKPH24GeG4BJ/nttq06HfuF+KSwIPHw6ofLAAYsQtxi6tS6l+
06UnKdWsEZoEhVFAuyUtOVBUvzxWU0Maq/1Ut63/iL0FhxlRUl/E1eAepo2z6KAb
Pe5yPSwIuMAubLIY8McxeDoxALrsnVpcgpPPkVmtJS42pdXP9nqFKPbSlwgNSbQF
Y3KVtjffT16yrFux2mgn27ZHtFUq+b57kLxcGttm1p27XSJoM6K92p2bcbwB14JM
CsVWOQj88JQQEWkLhJznaf3KKTq+pcjT3pL2t/3ZE03vqKZFEzEtnNQxKg0RZ7cM
ZP71JZ6c6fcLqvqsrlEBQQYn/NTdCtBZLL5eQfSKh08wi0uWkIOsjtOwOvDurmvo
y1JLkpS19T3G/XS2MPgsG53Z0KLiHt1JAr5FIRz4FIsqEzZBzjkQPM2ZSyG5W1e7
IznsZj2rrjbksT9ZlRDJk9TllcKdN/4jOE2aBiz2gbr9tJy31K2H9lkuCCyzF2+T
RLu2OIRr/JncZO45HMWARb3zMz1GrgjSJwYv/oYFm9bvd8YY1thBp8JcLChGi+V1
qcSad/VlXm4chEbI0H5arr4pbnrSPvEcTP156BwyINYBuhEmALbotgc3+x7hLyco
/skZMbIyACLWZfqEDWUSs04QQ0WULCd//MW4gY0uBXAOOg73lRF0+CwcHEj4VquX
SbAjbI+Xs2FAh6Dg/wheXTd4mlCg7vOrOF0BmNtz7/DhK4azl3AVLxe17erpFd3o
CGdPzlfTJfSklfIMpB+sYn3RridJg4IA4XaVO63gO/Y2QHPYcav2tQ3E+miVC3kY
kpJOFCaEWwLowKKghcmLHdyK/lMgw3nlKS+hetve8fwiD3tmqQqOluEFfrCr7orJ
zwwjDhLJysarbfzdyHnXgSHsucZMw2NVywjRmtvm9WAeqI33ZhakUAFXa3f7aHBk
zaEsZPPI/EaPtv/yNGy9Y6yIM3Fa1SLGflJTD5FuNbnpJcI7p/kZ8a8E4Xlj/gI0
jyYZo3VIVa3jOyWOiheOTcBdXAzko5ubHAUclH11lgANiWa1R6dumgJwgrmoV6Jb
TXFsXQoa0uxNHeVP4CyVaoH2vR/Av/hDaqq3/Rjm9VRCO3RwBH9q7AT6wn8pg74A
3UqiLn79XF2ZO9lt2+5l8352HtJgSaTJEGCxon0uIUVQQfqipsG+xPsMTxLJH3cb
y/zmyw8Jy6DiiozwES3IAY4lwHai21Lx+A5tfi9pjZRDEpFP3kPnKzwpIWHWH+fd
BusgrNhbYeBnkXRKICnU5TK9fHlU7nAkfWTWcYRMdb27uTKsBhOvKxdEC5InJnz+
XBzcXWLpOKy8j0fMbwIHXmrbF0DEtuad4KS+hmIkuGwzI5MGFDhmrgLJ3BF8hVKH
M/gnZOymw9udGFsorOllEPrD+Y1X9CYc3sxLU6E6XQAXGzUFMBF2FveXOnCirz4l
4o41h0sQbPgrKx9Qfv1d3qpBprbqyH1QB0VPbbndzBbbNCkVLADw/REHzpBv6LHq
3VfR7J9m/IFsxdM7whKdjPsLhKXrU0xXdOaOx5gAb2n+36Jw6Yh8Ki58k4DlNQj4
JAU6BFght6Jl5FDaCCiGTQAzioU4kWOv+cFOJkOpYDXkS6/Xsfo4h0Z3KLjtzb4g
iOvKby9Z5ibjNBPnIDs9LTO7Y46fPiacIF80RCUIe4O5cSJ+Nb4U1ZJHZJJecMca
7WLTi08gpfsvhSZqfGEwM9E513T2OhPpYKANrWhwAkFQq8SUij2iLCCOSC8ilHzg
Jj8YANDVBNkE9shNw0qBMEBJJv/sfN9eXP/BBqIui24uG4jcopNghULaFGCLM1uh
RoRrIv644MeY2z+hoV91ET/Xk0F3F8eHgQVWuYJSxlroQSj0ipJGDAdOBnyvfkVg
VxvxoRvlTKCHC+Hrn/zQFBZeW4ROUuKiISluB13mLwkk2vb/7ZCCkBA/+cy2kQyL
ScNyIItIEOa/UODY5bdJPxLsbBN5Z+ifrsJoRVrfVDxhdy7R23+TR5KnC3Cwn9+u
pKXTthuQsQXgsGWjueiY876VviVg9wE61Wwf6bRBHVpwmpMG/+RQyOmaovETVOjP
UnNT2lFVqPQb91zOtsFhuIC9eZx6aNobQWzZG4xjZ6iqzbVqq9zLXciJzUw2xWxc
0WAknJWUA3tSZZCkM3IZxH+lS4SigaC6QDPuyJH1cyD/pCuwsX7dHWTZ2SNUpYaE
UiICzWE8v6KsCz6/5PJirwh5nBKYdzLhZaM5FHFRUew85WG0ZfIsZzxLl0+sq5gH
xrIo0165MWCfubgBLFIx9BXSNDkD2+74/VfOPs3sb8184gAHC4bKgeSF26nWXkp/
eyLArOy71BLjuhocWGXLqFx4Kmg/jHT57Mf7/GA27ziNKmV2T0U/nBdneiB9SAD0
cNonllKHFSQEBQQzqfQj57rig3Y0q26G9FahW9ncs4xwkzzi8Bqy3KCt0IhYK9Cj
w4OPbhNZOSSPMGlmCi3CxVALIPwUsE6+dE0jlB5jP084KTF+i90LLijE4obwtHos
+lkQKdurgzbfakLwbzLZn1Pp0lrIyvnMDCDuQgdnpuvzjD8vkAg73Ga3Ik9y0L1Y
BZ/wmNJTr9LreElZ6MPDVUrq7UMolwXd2kZZs/UmrOLmBAQGY6KD5q4Wxl/qSdLz
ya+SMb3Ptua9OeJq+T6eR7ZHaS/Hm8dzbKOzhHU3N2bredptyt4wtj2crTIax3JD
0vlUo1bwXRz2ShrkhX8sFZ+l5FKbZysRWgyCRVHn/TzQXwDX5r+f9rdutluEYUCk
KNowyhH/XuvAnPwspLHuQ0sSMeeOoigxC3O5UHGvBXefFMoZ0ZOZK75ad/zDmx0a
6os88bICknIcCdfr7IvvqSLOdlI846fB25XWd14ODFJj94Dx/P1T8qogaFQ3RO1W
s05MrG3gBDIUIh7KGlE6KceObt7nqUYMpUJSGelgNUQJ5uPEIffNXBOqbznAKat4
eh+vTM4HTW7VxwVj50nMNx+4eKL7lQegpNJdmtXm4Qh4bRDiECHSNWCMyX6523bJ
TfaWCE/J0dEd9pFSqJDY2YcO4oR/VLENe/VD/ZZrMMqu4ktwUgfQhwG0sMeGMT3x
vfxMVfjTvCPKOxi/L8KNeG/In6OZfrehVIxKeWUJscsmiZRXVrCRU191hseGYs+q
o3kMg/Ez47KLge6SRdszmtdevirCkJAqhNHaNusRfIDGH0Dsw5YiSw2mCMkDBu1W
HLDLxbwlBTQOTtXPLhxCvEzWdNo71Tv/5rj3u4LC55sXDb9ZFKkLv3UzKBV0uzGr
A2wUOsY+Ddajue37ZepuCfYiFZXfnnT0d0AqzxVARnz/9O5v8PvZqYOXmxbcK5F/
iNbFkn5Fdu+t6A16L/OgdGGGj3OEggABKfwRaKLKbfMZBQnyc+q9YzIfpGOi9niU
4/kauJuSW6EWZxYKPU7Pr4ShKXZCx/lXoQ9CntZYhjhziOgKAZ6vLzyaKcfu58Ef
Ovqzw/HO6vo1nyUhSQEWND+ybxYCsEkdfLpM/JYm6xdz5LL+KkKvyZ8o/bn3P8+k
sT3aJ3jUy2FxqRiXgM41erV9if1/xeq5R/nX5zzxNe7DrxRRCNoMt2mB7s7DBCmd
bAmzqAq3uWFDTFfTaHzDsqX3mHJCZEwvD65U30816O32HS7zBS1ZJhMmdcAbPPcV
tmDPs6Vd2AxM4ASFwnhHK5KDqo4xpWKOIYTjTMC+EeZL+1bG2+aFfWGrTbfKzhPz
21gHxVn6Dgorl0ExhbvLdZZ+27+e00bNvvVteOEImLfLRmT4X62wNaqwYc4rRDZQ
cwprtm1llWnp5Z6jfzrq9RMYTwSsr4g4M6aXGUd3B7hnAenKQ5SuxCLVcpJL9Pxp
Gu8hvD88p75q1uH4XRB7DdAWi5SWqwsdoUzvzE4R/it9tx8Tf8KQfi+kgKvpGQq1
dvT/xf9RMNpyxtpfaYSIjqbwJf8Ximuc12m88xz4a9yiDrqPKcYbDUXSk4jw8Hqv
kyAPuxD8J8ld4N6vfDieNImbAAY1dWj148dywWxw8xIodh4r9UVO4K8oQ2pdavQs
4iSgeVCrAfTHlG8aQoTKl3B1HCWwISnskbD5zDEKEWeWKUTyfMsHSmgtlvAl+qJo
TWMfY2EFI249z65sU7CvnFCZEVWFbAYo27dgBGKMuaa1iGFUFBPnlGnYaLrdEjjF
rEFrsU3bb9slRWrO5c4FHOR7ZCpCVxfch7QEmDVBRnjaxCNgOoMwMqMnLOnbHhwA
0sgAtHuN3jRqDcoNYtHoho65VocT+axed9G6sqbAGV8jMKRuesGXBrODS7uO9qgx
IXb9GeY/1/j8nTx+AXF1NlEgBURvI4zv8LTjdDM+VwKMBBakCpC6O9cVOg0WfPG8
a/xB7ez01tXSvbj+oCnh2iSNT619b13nJ2mvYIzfUA1O6CLHKfmsSDnD6lckt7Vz
gX3A0Q8mQPJ4+ScX3LbZTeAKrpczFWwfp3dtkxw2QX6G17wYobpuu4jScFO9t8Vw
Fc6MnP6XQjlRy8XK5m4umUFli/Nk7kV8Gkt0VR25YCgatw9NolRLaRKUJwclAAyA
mQb/WeMnXLvT5HFmYi6fQrSSt3Ed3uqktpBk3eJZfpsJYF/4101EpL4Zi/aBxdpi
CAfefCcmhpM8mTVwRbPF4E1+Mxx1mf4wuA+ns1JtBFxAkGW2NUIVepBCMRiA5qft
+REmp1pW4gvUqYvZplVO+ouV+l/4F6vpoC4AXka211kP63ZppGmfQZ4qfuOCfucX
pL8AatMG7oMAtp47Epta8A5Ol/QHtVoC90w7eRNj0Rj5EOu+q7/QagQYrU0O5Umd
pcEdMMnbU7T/J0UaBtFospbKydDnfVlEpjUVhp190DZO2kEwIYPVLRQJ0AuwEaJm
j3P5h5pILw5td0C+Tn9q0md2QgLYQ/7UPMYICmCg98VDD0Mj6zhg+AlEo9wkV1kD
UplM+gjtjM9tZpQCs6jawL58zeDA3KnTa+9JitF7R66UK9GU0PUEmCauRK0jGCi5
2o3Bbyv+8ezKqUM3B+MWsisFLMIfF/s+sy14NnZ/i13/DVenhyT/aQrPTZpDjw7b
DrRDijk4n/W17T3P8gHnr733xCmLiAeBXpzFqUEPbc3hte43nWiuzKQnBHqMJuqR
eCt0+5PqJAhRqgrSUpt/5GC8ejuuf0wgUy+LYDtv99SJ5G+irvXiAMKlW+BtT4VX
WtQfwYZkJKRiXYNfXMessY+yOdAMTiAEp0cIaGKErIz0z5sIsEbQMCkPgIYgXlIK
Zh+3fHMy407CdVmADKuLAGq7WWEcJ12nvzG11sQ6osecT6vR/Abfj/+pcY7o6edE
3Jk5rQ7pLMvvlRhzs3Pc1t3B3G+9RmFilyBJqbzhnQ3jtvi7hpoel3vYUQ6M4kiF
U+U+IHVChK/g9wGnlz/bjaeaio9I/B4Qid9ppk6bkQY6r88MPr+OXvd8BOxJzHHr
9B0WtfR8RBYFvXNsmYtqG8AA54fxIasYRc6AGNk+hRTCgS4XViKdIhH2RHsCcOkj
qUV4N3EcCBK10Q+HsJ/Q3xPOqwKlmqDiyHTRVN0gxqBQvCJFIvO5TJhOFayC+gR7
vwJ3UD+nKYTL3UMTTKiqk408lKL6eoxF7MOsc9sLJmaMMcn7YfYEcK1mS5dwWDI0
cpLtga/0K9nw5+tqplLEH6TTJVkd+RemBpsaBxi0jQGTA+ytGEUTJ9C3w232jMol
8YjWEVdTbtui5bnfVBFq9eV5qYJ+0keNicCeJj3Dz9yPf659wFeFSnzXWHU1obT7
EJYKUDNx5DrSgRiBvLfsrK/bt7pniSNqtYVKqjDMLtFcoW2yaE2QYtPXKN+hdlY+
79UycLJasrFWgbZZPRBgJ9sh6Me1mTCr3FvNGiw8L7vTxXHEPnpexSbIJc+I17co
6Ws68orMeO/nKmyE+zQwsED8pAdOSlxIho93A1N//7Ys2eNHIjXEVVK8oP5msXVU
W9behwxP/Q6tF/WSNSgIoDHYv+3YVN6tswIrao1nB1XSc45HueGN8m6wnnEaRl+g
ZF397Wz8s9bLM2SgixpvG/0K48u6NH3g0xtWxmXU6n47s19xR4ejVlZi+bFVcUkF
pBHETkubvKANGNL2he6ASteGcBPwOKPfoqYLTwfvqHQYLsP5FNst/WXDY+cbBfoW
n8PvXYDW0HlkQFu/QcLNPRowsA1uDhjMNVGGA0ApUs1APiQYw2ZeNY1EVwq7CZFQ
w6p/RsemL8fHdh5LYfcOeJZ8KEROMv/iaxZXN1hHRL/ObX2ab3WgXmr4iZ5EFVxT
JrCLrBhTfu8tcqmJ9Mdb0fYifM/q6y1zouysfzPYyeQr6mhZCwB8f7vKsuuDIQdw
ileeqSndd3fG0GsQwO1YqvnON1uMFz00+edYrnIe02K76ALnrE3o2yQlGsuf/qwt
LzYNq1JhEMB/GerK90JPK+pWEUoMkzeSh9e2Pl7BBQJp+CFyA/HqPtexFgHjIHN5
3HOqAGY5QFsKNyAIx79ni5cTdlYAXYYQSvfl/U9e65Ac6MsJXzEc2nbo/+nhQ/Zc
fFB4OTSGcHrF4tzuKGiV72KVczd0ihTtkjVBW+YNcLDuRwMM9u3wgIgkWOOEkgSS
vIzr/kRmFptYrHOhJ6RzmK5AYQH2Xw/Z7FWiNz2nX2K/QcpIrqPzv4RnZqNK4pTr
CeE7w9JyWRTYaPVefx91JQ19p+nuAWT7n5UPUk/UlCx2EaBRnV2AgJoHdGUopGIQ
2+y24vSiQpew+UTepJAhmp79g+yrbWZvNG5OLPhtJyhPY0pJl1jsheGRUfFxsqrS
yCbWOxWO6qlnyFDioGXnM8dHrnUXz17uLzwAi8zPI9MtQ6WPTj5frtTgnqOgVsoy
rYyBo0fTDE7V1GK1b1cxo0FXwcKIieEbnv7GBKHA8V+7aSle9J/ToxnVZFINvgTt
QAkFQFejbF6j1ph+KdcWRVK3pdS/8sVNwEc7TPTwK1smaBM/O5MP6humj+Dk8h9C
5QvK3j59uWTO2U1a5CHxcJn52IJLhuZ1RhwJkC8PFK00IgGsY4lEvScVOGKJOiWz
DQuUr9JA5HIbsezLhKrnFKlUmkGkgpY8mWsXNORmSVZm+S+/RWv1Ih4awFHk3h4Y
KtO/pmWzfk46/pA5cy1z/dvVHudkx07AfK+l206g4/uwC/1Sm+BOI3n6Z2x9LzxI
uk7i2pk3soOPDxMlEcZJGhmhrlu229TvMbyvhotNZ21PuBKC/x6kQaRhv4clJ04/
0fCmN9SAyVuAqrkPsJMDymLDltLeATfKNl+2WBwRNXsuDIZvOYcbAP4A3VEVvZWa
pzOdOHBAusiIv9iJzFNrE5dwRPygkskDGl0TPDH3nmlUPigl8WMCDdBI/Wfpgc0+
dAdL/8bygZWHwk5ayT6I0E32dTjR4zMDllRFvWnmRSEFWweKvObKyQEuUnFoZe1M
FKVAXIiiDiDKk8uOiL+C1nnAzJnoWtbxW10ycoVQrLyR8CxgcBgSqAWLnK657rtZ
s8ndvQ29nHCJtvP2IgUD+Yxh9LCysCf86Hr4+ZvyRxeiqHMAslPVjwo5+cBkrlOi
hHxC0lqy3RQgEZ6wW6RRoWn2LKs0SBpwl4jile09kh7L34OYbdxxQLizxawMjkuT
aE3VXWhnWb8THx52ifpVKQ/FYniN70teH86UMH9zqPo3YgcTkMuD3MvhNJ1UGIV3
3LbnGf3EIa6CUhXio0CsYWFeGgiqL2JW94jd74PnEATqKvexsSThLg0bgDMYR4SJ
jNug7IfOheJe8uIURGE1/x0B1mO9R8G3DzZQB2zcnpZyrorLwf+sP6AYoGbxRv+x
RNgm1o1Sm/BmnWyINdy9se58Hu3EKwvGd/ecmESxTyVnIaIV16m5LlyFCMjdrlSn
nDdIqofotobkwxsjReSbXp8gWl80McL+kORjvekQj/DMzCnmI7WtudPmMbJ96ly9
w4Zd64L2OB6haaqCLkISLFWWc9lHOxUNQeaEMRUt9Sy2P72zsvoU7NDY/v8t8T08
Afki6NEsU6t9TfgQwdNEwR4snC9kGemvDLNJSg7LNTQlHXKYWX50bX3lAvqgXT66
DLImTk9C1GfPO20OOs6ZNQ7045iTMeCOE3y4vgiHTitMaCyYweFiYZr7ALySTBjs
fjBcRrEmQAU6aPtPv7t8v3Gag8bjSDFf5av+CNQtga8Efk75hvaeYrcEcc8UpFM+
YrRo6dXIMgejp/kJGumNiiDauCAiOkxiTlY4xOR2rHklJCedsdn64wYjTjttrzbM
XL3X12/WQ5NiiSNNCoo5/mVwIr4cAQ8fGUjP/2y+Qydk7C17WKS0N5wxrVWON61D
yO9ZF+ge+5BrGjo81eB5soKHErjwAO2Tkjwlbc1jDG/iFx6ac+wo9cQ+DLJI1t8w
yaLUxAfkQ/+I3ZyicT0aZaWW8PSriBqFdEs5J4wYCHNZ5GGGi4cNfkMTO5YAUmib
Km/oFYR4ulMhwP3MzTQHEfq3gsQpY+U/UYkjvVa7mPWnPjlFl1ReEjyoi7VMlK79
8yaqF3tEtY3PLkMyaysZfx5FnuSoA0dAoG3FJKh4+RFVQxS8AsNxfFOiXHneJdOd
HnLdH64PKx7CBInf5Q+6Az8VlD8Z6D7JVrqxrBJCpNtJk31MV7teg6Phsy8d453B
1ThxZd0k0ls00isq69L1UQBG42H0b6N/Go17taD7jajSb1vh4T4topS/ijWOMDRq
5aArx8u5MH1FJfqQvkCbD8a0dHG8iJ7H9f9L9ftqnnwdVOMT9vKpHzzuqJTxaXPA
INTq8eaCsiHT9Ql/uDIV3MSqSTks63jva0VTnQlkt6kpOcj2kH/0qMjX1ss4jZ4b
HmXCgMuQbwaBZZlUAPwgYx1gIvy+3mEBLW+ZZKDBifRQpQ65DXpAP7yGiOQRXlIY
jOYp18thXcUgna9DHEj7DxobIZZ1wARiRsYCDEh5Fxb/xTO+JeghGXSTZMgNRSaP
jdSkRSvCKq2+4lKmLEhlCVCTORylIHDTBKwBfdZ18hq1Xg40YpFn6B4u1AWxkKCt
oW3KET4OmHk1tcgc5PatPCqHcOIUUKz/VraIQtZgKNWX7pz+DJwrUy3CeHwBpZdS
HYms5sZ0REEy7+F1vYf2KAD1zc80xHtPU4E16g0E7I7E9vKk9UdTfmtUfcRspWNa
1AFsUB4EpEor0N+mLPDbbzlyoQQBqAwAt8sK2bmfG6VyfLBA+W65zklcIQIKzytv
DcV7SFg2N6n94u1COYMEruWYW1MFc81BshQfyg7z9KQ=
`pragma protect end_protected
