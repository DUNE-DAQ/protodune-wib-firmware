// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bX8M1lcihzN4Q9yHV2kPkZqLnqSPwiA6xUsasfW0Se//ItRSbXYXmBC8Q8cQ0wyB
3GUwHStTjVYe9JTHicHJLbWkPBt1d2dwMTk0DWek7X4llM8GdrNz2IHuq2cEwyga
FutPszJJp3+WYdDtrgicAalKH6HlC6kQkTwEqoKt254=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13104)
6Sgcm+9F7lOm7jAVnpba2f16GD0CI79mYWKFW+BI7VgcNA7aJUM+9laTbQ0QH8UO
qVkIw105I8V9yQetDE75AVVLi09EULowWV0Mby43hh3LVWy8fesakDgAOMSxAkFE
ji2Uj6VbLqVg1QKbdyxehXbIZqV8wWFGNdzYGyh6wgGCqd+JhbWGb9G3sAwoMOm+
740fEc2eUGjuF7+Uu9AWkIFcJubOi57CM0ulIlwxtb6a9r5XxRXWyV6nmbqq0vAp
7s9eiQ/sbQ0VypK0r7rED14DrrsXU6//lgEhf6IArEQb5iI5ojlcY5S3QL4X2ENB
uPpqS0mpprEHYaxg+Smjcvp0z13ARcwn7ZIYOYrQCEz91c8jTVzfNfVP8MkJx7KN
AuxYwtLGXVqU51AvX0q41k6jkfyzEe6CbiklY/G04hkqsG9Spns0rsV138ui7W3u
WhUdeO97vxK3hUIHLccZLwxvZ8R3UdW+sBhqhHnVx9RF3NzCjJs7XeVJ6Ydb1pxV
bOlk3w7mYLjUAghFbRlzyWZLI0hv3ojN0fAqb/nawfzPx1WGn+c+WSKACatkS4f4
JB2fryCDyqORxHi8Du2mvRd3RFILfB4Uw0t1IWghmXFuGhTEjwQDYXacsY1y7Bq1
Ndt/Qhoi49sUP750Hy/1sYuLzvOtOCjSB3en1JyuZYYZl5ind+zKjyJ0gJ0LHiKi
jsvubZ6KUB6/SUDvx+MK0k66GqJTu+fNdhJwLP343I9C+pcD/RMpyMBmb3lc+Q6D
5f36aprFeKThCWb8LvIXhtVO8On6z2rApJuUIiCr7ZtrEU6IELo2r7Q2u13ft4N7
RaAxFTFty06WTQKhaT4MUGLmYQOX56k9+/iWmsQ4zpRJbwXHKyn+1jjfyLdTaabc
k0qEqRrZAV410ddU7AVDgiFWBDRbU7j89aYylHceQS0HHmB0ZICaDqwIq2QYgSv+
BVJCx+2ZwKiD7O1ta35FnQlWjPYZnnIwbKd+fwldWkTUllmWg8LjoiNsXk2pf8FQ
qbCQ89Pw+3+JV5XHo2gYaHUv8LsGzBfzA0vc7e8WcyEOBO6OVfKQSQ5eZGqitHBk
i8YAqz6kQWq5K6fYO5iGI85Q7MLBol3PwebKwpn9rRWpy5EQLuJOEh4FHawrIJio
GIXUT69K4dT5vKAOJq8ONbNzZRlswnkYjkiRRtrek0rDXaFM5PGm9gNXIB96Uwr7
7HI+DVyObuvjVw9t+hs5p1ZTRFyPrCZS3vaOEoguJfwDeg9N+GdnapYnsS55FId5
hVSshLwvUnapGERFpN0XaGyZ45pHbZTDYOPsJS3UQ6qGf5DL7ZwEmIdk73Myku+m
g7g2L6YlUduVTda85N82/juZHBoegngj+rOcRVj8DzXEzw6pNOcDbeZa6/hcaXGI
Cx+/4WP1SPbYfXHfn4/s2lt1yag6XE6zYvtbEkfrg7o/Oc5OJCEM5yT+OI7ZblgM
Q/rb5/KTL22Mt51cDuIPjjV+kDfNQFGqG76PqCAhBRfysa4PoRvczw1bIkL7Paq1
XfxFT93xCpTjykoJ1iNu9MWq921qRPKDnAL6IATZsdD3kwo+0u6XvLPCyrK6POcf
utFKcH43kwdTXh1veBAH/PVJ3i62TdfKkBQqSr5hivM3Cq9Mqc0w/xIkYtYIQGJO
Qoz/uFyjKvCJu7YGqL6VdqojcJkE2WA11ptFyW7OsVKbcRFM1Kd9el0M/TE8EC1A
eWBHTg4QowiVWuaGnuXUWgGuSUm4c4HpNJjmnytykHUKXyj4y8SZPHvWJFx9BJ9h
uHvc368bHo5GAKl8p1JDu1TUW2FEglTwoK2iXGVaxCFD1AMjqTxln6yzULq0+DYe
z60XZCrLgPBWhCbtC1wg5SfdTtu3QGuQ+/8jjIwfg62v2oQdHTA1qx/30azMNoZd
ABUdNo736uv0enVRsUu6GXim+QWXC+VRxH1B8c7Vl2CX9VJr4daEROiu1eBa+lQP
NE6Atvkw8umha+m/kJSsMMnaUi93//2LN0pcPVGrVCvqYHejIm4CBcGw8K+WBlbT
CkdAhZ6FOsrcYzA7Y5dlUWO24s6YCzB6kkhcIX0DPZN1QwT07Ya0BmNsLE/cwab0
NlE3rETfjHRVH3mRNtIbIR740sE9/QzfoiBpYxEb/SfeTWlYFZlIbl45ProPVlQ1
UIghQqBwn52pflIWDExDb19V7rgkHGmX1ePRj44EO7fidDS90+pMHhLvHq1Z8sJt
ihxHSxUahuw+u49ly4CiqAzBrAuakcC/AB0dDT3TvNlg+tyH5spQ6gEh+JtAiwgB
3WadPnvu/V9fdkHAEdeq7ej8BrdrsKRlPFRh73c0xYQOb2QVOPcFFphpYeUbFrzr
k7fgAOjethSKgp6lqgTMpaa9WVatYBLO5gLlkMHeKUCGyJvGE4XUUdeo+0TBacsX
L58xWpcvIjxsZ7ctp9wmkPEFSRx1HrB48jfSSdxEdO5JWE5mti69QBAISc4J8em8
mT8EMp9K9pKZ5ILNgndIak27h8knpqD/Plv/s3euuh6Z3fqlCJ1uSvlqdgsZY2SI
e/nHhh1CXfWojvZJfMK6nkCR0OamyV/ub1IuS7NeIs3cs5ASFOPK5WVwbSFOgyrY
/KytFDb+uM3vaAynlRICz20h1JRJuk9Id/jZSFRxtXdh1ibOggkLh/kaTrO2KLvF
3Ht6PMJnaiw6t4HPG577FXD7U7HEbvs7FgsjnmbAmGpymr7BufQfyW+MugMlG/qm
pHNFN+oY+nE5SnIxlLc+VNHe3Q2/7axnoDvVVUaaFjr+JhbqVhsbhUT2hssPoRmQ
iz4RFvuk8LtzSxzbJzKLMK3T9cs+s+gvknUTgYuQHcm/4J01EPMnOxinMqWBMmb0
7s78boYeUJvwao5ZBm5EKLIisKpli4Rx0PmEH8MO19EFuuSl6eHJ7TLVU+aCHDdI
sra4va2Djfw3bBVv5f2Mw65TvXwILJCVZk1WOoRlaJub/7n69ErVJiHa2ymGUFFJ
uwwFcKd8JCBPkSeisTBDTzPbkBblrzcsuhgSDJBgn8OmMPsskkp5yLTd7PMVHXjB
Gz2L6iadS5rQ6Fj3yWy3HyurgREVIZIrmOTCOX/dlhy90GXvO1CST13hcgKYBqXX
CAnZHZ1VnLx+V3ejZrFIPEDIikHX6f90m0VLCX+TvbYrxiaOf31YPr/xz7HdJM85
G6FA9tmM16b3Nx439An7PtOGtM4CuBz4k88Dq3mXS6c7PP45zn+a0LUgtUntndSu
LvlT/mPXzRNXNNrwm4b7XRqdqdgd10T9rzSpQJ63IXY1DmFPC1by1ikRlLH1pC9T
hSHyX29hsuflSTGaSAE6PsfZOjm+u38jhH5InS5SDg4yMHb/lXvfFtHCDk4vECj7
OwVsgznOuzb/IiTXLTptOUGz5fSLnbMZVPtdojXYZ2STR3SK4Wn2lssaAdWdeC1J
KeNoC+Nz3UXYOVcFOEHfg+fbrACtc8wYrNTz+MGaMM9jYV000YyAE7biy7nfIPw5
lvg/OzKINREUrPEUMzKEDQ3tbbCWLdzjHGW+dnUfaZaxwYM81gJd2S/c9+fXIPiZ
zw8j3Bj6H2mc2wa4oMN1fJfbb4J29IohBhPpD/4+z2UW1e6o8ZnWU0p6XNtUk6kF
6rAJ0KlZX4E4p9vo7V5cZ55su9O07mVKJykbN8YaiT0m31MRucCVeGDrxBDTDYkB
7AA9MZenhX9xy9hL5R5v0CCH/y5b4aSjGHcAhMtovmqrfXLB8X44naYwrUA4tt5b
L+p1f7QFMNRTXIe9OvYxZwVTIhHqemgC6MO2czqMwaq5oGkK32lNZ1bD4zqcf0yy
/vwp216PRZ4Vvhcf6dkF5N5uuBxl65hAwWtEnPe5WI874SakkXMoqOvBbXsU6rDV
gAzYE02vlR9WpoGmseT1+XI09btQD/ixTAKMlTT+4hgOf6VKZ/lChnZn++1Wkq7l
GQvrPsLWJuGiBw9KPPCDBbg8wPPY+OyHkbog57iGxuXkwG2//TOMzkBcgzXhCGCS
ZZZLwkP1nVL/oG9hhH9jH/LzV9gNBdBwdFeOGVusZ6YjZEcyBVdhVgEuX3QRr1tp
lFKlAjlnLAADrt9Sr6cyTd7k1bZVcyuc8ROe3wBcZz0vAWxgmAU++7gn4agNuyH2
can5Uw8pn8exBY4LMkmEospuewA/8EMIIZddPv5+t/0BFkpJ/X+X9MSI5rx0zWaI
bhdLO1fBVJtU+WxgAT6zG/im2FQ6u76iGmeMc1Lz9KlN+TgBmaoKY7NzzpUyjLVD
9m2Y+0KoMwHdOa9HueS80p3Okj/eg+Hsh9V/njE68aD0o+MdPRsV/zQdNqdehFLV
YjpAOd2HuCWi7v/Kixr+Q/orTCqvuxYh1ziCzt1szOj01HU5EssCSazn1ETeN080
RBLm4Vh9m6UiHM5kRRKU2L+HxOsd42Y+t/T16XqrH31v6w4NEm5YOouPLu8J5bHl
cLV6ShAQBHYDNkjtEWlnqdrsOY5E34+QAdrtwWldnlAmzT3V+AcGq2gOnB+rwAOY
vyKACgEZkk7IWPOxs83JVaT8AWo1ZULL3s0GwyLvidajiRNwbfP0xX4I2aKJooID
3wC+JVKzlwaSuyReLGO03L13IoFNLqK5h2xENZPLWG4TD3daT4CRJ4XgViXLNpjl
iLX4Hy9xmXVDd2PC357z0hFYGV3mIPnadMhazmIcPKpNbYQRGL+9iFcztVZAGWem
wZ0IkIrP//iBwQvui/Jwmcg/63Boy7cidAns1xE33vMD70FBCpFVqs0nS7Amwdny
eUJ6xUtiD5zxFmN3Yj+VSFDfJTiQqxYFWj9OZKM/7VGmX+AZXKTe5ztU2sQ09DbK
sLFV1jpgG/7hAuIq0Is9/96mRyVKXkgR4qoJJ0D0olkgfKyeZRHAA3n6tOk6rhk0
9CISwUZ2JMl9UxH4IvZy7gzIz1nuZa7uyw3XfUEJuEdZolCu9xdzSaUhfyAtaC04
qiehrYEsRiZR7aN8wZBDNEa87+ISC0s6bvvUwK68HHmAQoL1/1bRKJSQuKNT6nJE
n8uTetftggei2cUT4FTRXBAXHxC607Jve0cK8Hrb0rWBYnZAJUeL2z3I5IcqpWrZ
eOIYnAAzfG29cJ8EiA6OUEso8g3aoHXMQhnR4S4Jz06JWl7RHsJ/evDMRP0DBOL6
nmSo/a04ovS2O2kVr793p9klW8qDZRfmJ/MsOLn62dsOHEBEMuCAhH8Rd7Z5qAdu
mBgyshL5q4UOSn/F+J2bEc+Vv/wFCZxwaKpr/kO0v5vVY8lv9Ecw1R6zVuh6lAh/
3+DkMtGUhe1Knw9bjcI+Bn8zWMjVUczjrKWkICW5ZNJuefTqdK0/yhSY7mGy+a5b
DYpn392r6LgBYK7DHwg1X/t8ObLMaD0xqVTZB7iRip9WLSlitvnSTLEiq3KfsEza
QNLijC1VzzoCC6rkAJAmpyX3TyB5dTCXAQU4smSDjkI3Wsi30QKzrs9esaReNtgm
CM3wQZH7lSrVv7Zp8BilTqk3mMrB06SfIAubqHjxx0w8lhuyxUmXt0cm18Ai+BZz
2noyozUfnjYUyuF4vrXY5JCO1sQQYlZ04AClmcAoMbvGMvlCC4N1KGa+cEFQtPEF
e5NwLOMQoDFWNKyv+QBZsBow1b5kFKObAta6f8CdxWB9ZeIs3JF6Oa+eLQ3NDR8U
A7E9EaisMoqiq3Zduysy6FsSYuR0LLlLxgyMU3dCh3wdXtM8eg4gLA2BoV2eDCMx
aWcuzUqgYfHGvOphnXlTSAySa8CAIvU80SnACn33q/0scAq+zRHu4sAK33zph9p2
zu7nxWRCocIH2Dcg5DRrsK8J51gMomYpy1kDZur8tWtIiA5W2T9uwQFrraZpRyXF
zILpi+EAcVRE984R15wZ7NoKOFObH+ai6+XfEJLdCbshXmlN1xPG4FN2sndVaJGk
5hHHhyIcxRe6l0IT3iUSbE7JiIK2JsqM24+CLf3MW8Mn8MZAgLDdhGQv3Tv/38AK
LIv30olr2Tk8eh6AWmIrLWqzZF8BUDhVzJb1ISqCLuB/w6z+tJfsQrfSw0ieYiaj
166q5VRFPQ2wapPvnwsW6scr31nQOSbtj5rRiJKEIOP1OpUsIGP+eIBudnu60qz8
fWoRqdiDF+iBfJUtEVQkhwCDg8PgH8BaJKYfU/fqbHejVs5zqBydLu2BdgjyQH0J
0nABnb66dbuCUk4+vC/7IvBcw4iPAngZJiMulxL/TkDgnDZohwVu2uRY7uxkoEmj
pkIhcRYQd3+SQxaZnEX5dSqpsW31aLTka5rcgqOvPqrqBBgyslGPqFjlIUuGYLwg
rj5vO245mZODpXAs5GqtKI+ydYjeYxDFxRMaJJ0R8uWTvGMZ9L4AO3TBnlZd/MVP
BZNGQpFoDNY2v93RXJqSM5n8emh/r/5/V+G7EK/DGKdRN6fO7TDpllEjs8vhDU18
ivV/2CJCXSvjlC19MlOjV3N2G8SX87DvjnYuuPXkQL6G/5Fh0XI5n3+iY427+23+
rtiHxBVprjuDJYDxsnDBDuLWYw2XOKZgh+3vgICp2hRQxTwBJY0u3UH5nAdS8SAW
3QE1yg9H4XXsF/dt7WafI1uidp8ANaUJiCQlLpD7B2aqynNidOzl8UUt8DAxmJzH
JwzWzR72eh7AkhgCcCOyDaTPdHok2bjn4xYMSsYxReHaFJrdVeWCD1+ml+bXhIkQ
oWlqYGz1pCKNT9WsoTr/2b+tO32u9jMjwMeKwTFlZdVacBxAtqDNDzV8GqsHG1Or
+k4GHv8QLbi0Bt3Yak53sUK/XXDQmkwOziykpZd3koxzs9IXBF95lYl40sR5v1Br
w3vjYiudfe524m1wrySuIq7Be0Qz9R/2Gk7pG+ZyxFTStpBOcw/YPSuQDPzPGupt
qfZGREjbW4VJG1UFKuKEOd5ARLCXNg4SwinDj+dqr5wO+zIQ9dbo6+R9a6rUs/BH
vsrnsFu9e7lsHYTYyxQmbswfrfem1SZ9d+J3mRhHU7T6Qgqm6VN5WpySB4ntLgeI
FQ/Dsoxoek3Wi6tEzU5xRIToWi6DI1uV7wzWdN0vdKq986w4YuBsd7If8Up7hQia
+eHTdvx4Kus5VkLnohx0GOa2yTP7GxHywpq5idMFXePENqLLxffqEml56ow/bAwB
H5epATJe8PRVNItC1E0TmPbs8srBw1TRTlWPSS3pTDmeCA0CeJl8wO2IDQBRU76t
pHcd2DDSjVFX4yeoB+xQnM/dG+cc91VrBl2xs/4MYQ1Xmvyl6aAWV5qEa3HN8xcl
4MlxQE2lsfMivozo1j0wNFeIBBcuQXnOAWKW09SZN0vJvU+jdWbui5sk1NTzV3AX
z+9m1o+y3MilDnPvDhi5DKpJJWN0NvzzLP9aa+K1vhNRdgFiN2CYFn0Aev3vLYPL
UjLHGqd6kuIoJkItY0h7BsNTEwxVbfs9XDYPCrzdOBuQO7IowaBAdYT9W6u9UWn9
kI40u5WOiNQGHjuz/Mt1ZDVtJ21OGSD7V0Ejiz5WEHYh/KbDEhDIDSFswmiVFTjG
Nzt3eAGuwHEVSB+BSfbaK0HQDJFR1l3QB0AzrD8SaPQF0eKLdnqCOQWGalHW1xcD
vwFM8XXyRumgQT4necS0MlZCE4HLlNaE9YjIihOgzPUu+Ac2N+5tJog27BMRQesI
JlrlurjfSapCqjQVHhSJhoF5iXTvnJ1QzS1F8wzhdeveuKkP58+m+UqKnmr+kBBj
xavNw5l0L1Xa/KEAlJCzusDOMEPs4YNU+kxsZPr+0ixUdo5Ii0nbppW3oqH0uIX0
4N9ecIct1UxVJIhcfK51u1MaQ5UZAvke9yRYPHO1HGD6QcSGhoU+MelEc85HMTzf
8n5FkO8A2GZJky8Lty2BLdfcVKXFvlYaXTiNHsCnLVCINUmPa2JuilZURqCFBWw+
gZlBeOsHVmnApu3c+h0LTlSU1a4hgWC/F5VAwKXuV6yZUYqu6yB+9bRWBwoG2r+U
T9EL5Z/xgDKzKoi8cBb1e80hIp1qkrnIq9JzLluqaI0lobgzKRLlwtnjcg4s6stP
q+wcepr0qXn/7TAAv5tNO4kvyst6r5UVnvZQ/fs8vlMKQh06NJFwyouYXQJzKvql
YZ97ITnZGl3h3T49D8GS10JWQ9eZssmUTfuDSkyrHBajUim7daNBAeNpj4ZYiZy5
12/0cW/14ayO04T3CkUZr8yiCwK/ZyCxG3r04MvJE2p6SgAhhWoqZbaC31jy7KVe
Yp/LohOEVj5hev1p9MWCaxlhsA8HbH07cP/nCTzdiMdC22Oy41NWDmT5K+pNOGQ6
ovkGCC3sCU4v/m7RFB5OtHxFf7EPZEYNhArBc8l6Q7Ob+RD0Ay4tDf7v2E9hEqPm
FA3/qyCHQ4rDOZe31tFYquS0wGG51WpDTiJB5Lt6cAcPZW0Flagdy32kCtcYvtgt
buQcS0zjwmAj9Kg2EsJ5Tx0nD+egUJlpYRD2xJlKNw4TmDp4pBUL0w7myqheFkea
i/rctKyld2+ECU8tKCgXYZmC1Ts8XMstnKTvR0gl0eP6wW42qZg16OY9bMypTHMM
XLtcyz0Qc+XxTAUKvZQ0sDGyjuf/bV/JSB0bvfuiy8rP4ITQYaSwujeDxLXY0a0F
ENB7VWEDKchs7E4lBnMAk6UmPPUuF9grKUujDy5xrqJt4VbRl9Z3KtfCV8xpG3B/
0esGjr99o/wVJc0lKIb2bu9tZy4frN1yBkeoRtmXv6j45dGYvJY4SiiG/ze4W4vH
GxKepgyrXrkpVbzO9TPZVqw3EUqIcAnwM1tlGWzs2UsraJAKwABYsf8xEHrI6YS1
47GO0wTxgBCrYeFCNUawx/UA3jYi7vHNFZwSmTzx5Aage4Am58nGe3qwnvTYgSmz
Lj/wDrMSzbfMLny1L+vKZjczctE4L5h/xUMLQLhZUyhWk8Fr/J0jCTRmn0TTJoW6
zY3OZNIfoa6/Bf6NVF5wWdxbp1R2pnFUGdgvhLdGSMlOuvbtXOz5wcX6h4koiqDG
g8KQQk6g1ON+IoXFaXgN3y9X0upVlrnl2ousz5EW7UuqP2yqPLxCxdHGajZuS38E
TKVr/dHcEkZfCYvhmW3QU2V20vRozH2pGBk1yjphDJWXWahlmA9Ddm2xY8z/9Lfi
ri0484Wporov74olo2BmxanOVl7skrIt5gnEZPFQAKvx7Fmz2MlB3a9zsu91m0RD
A/beTC+E6gTIwz9vejAh3UG2aQWc1mGnqlhwH2HEuTFViUTnJNGY0cbDuGuxHn1R
UaPUwFzNMTJT4ChZiViYbfqH5Aldp8JAD1Ek3i4SFOuN199UXEinMldBgh1q0LTw
REqdFt77+dF6I6sEwxu49LFPnbwC6TemIBL0nOU9I+WIcA3kmuBsKte24g2Xx7+y
oGGkh8hlnDpNxJW8avWLBj8ScHgr4FM7dvX5GfNa79CXfsoRkKd9WYmo0fVksExB
YqH2wIiB9R2uXdBuPTvjFmcJmgG24HKYiG1jQlnM/HEstlb7qEWQyEx8U6nuvLMH
7atGb5/PWpkFM8k2JSkYkir/ayS58VNjoP1Z1A1RTEdajW5EBL5MAJRcfx5ecaLW
/G/XfPRD4TFEz4oOGekQqwHCPLmqIg2cYcSlgKp7iKRJs6soAayOCQwYq7Pb/w4k
JWEuX/Lp7dIvoICO1gwhHtoY+WzhnArANDyailY/KOVtqI601JmMZ2CTCx56FwN8
o/RIumDRTQ5TB0Uo4qYOdwADmx5Nf8TvedSerEk/WZYoQg70O7P5jH8t2aecNvUx
907xJGlxabFImvozKrP2VUiUJABzVrdUMwVXKhPR8CEUKHfDJguhkF2Q8RT63l6Q
zNZzLHa9UACAkiBktWdsSkWib0dS7BQBWMR/Ap4cXen741zApEavRl3EwMhsZu4w
tecojvaJfcX9RzG6OMV87m0O6AmxRiEXfdRQ40ZwmwXIagu7DRtJDwFeOFt3eWWt
q57RKnfjsDakAgtjkSz7VqwkDRZTL/dIjzOHxLlI1mj8Nc+ksE000/YIuBhp3uLe
rMCx0/w9AjLKqIreDIM5N/2ROZG5Mbx8hAxg39HVH42XJASxCF4yAPlBc18+sN0M
zx6O6QwYgDxfFEaWAnbV7EJZLcmnEwpMxirPkMYZ4qYjdXCUBw79JFWqjtrdogTv
b+AMHxSkgpjUkLCmnOWfWZyU7A+63Dj6Mgt+72US0Ky0D9UpWDzVwVrrS55CekD8
SMrhtz7sB5zeXhJmEDi8BDaY04HZdEtDMldrlz73MFEazSrcVgN3550gZOAONI+4
8qqV5RHRulD0xkCP0V450nHtboR0fBDJGVnp8+h2Xdkp1epffzcraLx6/LK0z92E
WG7JtFzSuQMMnCMi1jX3bRhj0gs7t3wS5P0e24ITaBgkGXwz6YJ2S4gFgsH4j+sQ
YG7llS0eR2I7djZSDc93zDnSjNP+buKgP7L1w0lmxxpFGFieZte9i2w/OLhm/twA
5JHXg+tyoeEdh+vgAGQY6lR8v7vc5vnXjtKjLQOdSFH8TCli+lR/CBGPxYQPn+SN
mKIVWKds7DwAZofyIieVAPF3KVye+5p5wmy8SPFTmpkqjT8xdDfHQs9kiovtO4hb
HBHSDID7GDT8MzkmPnaNo53QhNTF0AU5H5jcInJN7Qi/HZl5tZPaak7XVnLt3kD4
1M1b0tfn+tvLc9u3mIo9jj91Z5upJ4aZGZCbjr3/DReiT6MmUA83Is8TUf3YAY8o
4U/Ta9NJGVf4CE7wg51sZJpIxQRSy61jvoS022xzjFhGfIpfPU1zB8TLP+STTe8O
GuOVlSdb953xHq5wQmL2UAl2zvTvfxAt8mo/AMGxKJnMioJvXhJn9oYZ82PY6WlZ
XsWaWQOQART2+VrHDRHRFDUDvIobPRypFA2akQS44BYthNPOPnJCop6EbtUe+tbd
lft1zNfT6+JZoDQU6o6pvEImrLO1dflWP3drjgTaU1PGHzxkQg+guGeb5nP/mNqZ
S/+kKVcVFL0H5m6ZJckL2WeDei3nv/oLLdtvKPxLtkyNjMtYbCi50+gZ38dldRy7
fq2N7oeSBEV19tEtOt4PjJBUcVNutmKxgsBOFg19nUb2Rx/1X07Ie7vj7CmQfdYU
HaqmZZrrYPD2rWNjBg91kYJuSAExm50JOLcI09oZsDoHeDeEu39Nt4PMT0x26+tm
/KRESh3JAgpbQ26LHfXKLNKtQ1827z8FgHm41hHarjqQPHsuV7eEInXQwtLeP97Q
cUfjPwViKwSUBvXH3QoXgfzQCipOSQd9oWoDkq2lYj1p0d16IBqiHuq1ub1iPugf
9mVHTWIMrm5eWd4cFn99Vb0qINITbyiGt9LYuesQr5DIO9IUJ3rCBlmGRpHb7nTt
RGMJngAoTuusfB8opm5lFVH1jENO8+FLzziyleRdGRaKwcq63yrYgXrtVJU2J/zS
fP8aljhnrimkSv6lG1GJze2v5NllfsW1kupKZ/62R87GA7yoOSrPmGaEYVQeR+qd
/0xibQ/c5RouHcm3B/vPN19y0m3/UiDXhbz08cAGjHMNdI4XUTZuiAs6W+AruHAZ
0rMDfpKtpQnC4pASuJI2fL+90Nm11N9xmUhFyPUGrJBYENo+TFHLg+xxMQ88Yg5g
JMa5YGgKORJoN7D/IKIjU/lfIwBdQgvo1M7CLbfxMwJKjohhLFShaCNVPTFPoHK8
49KbCRn6nzoN+KGRpAkQXJOiHjrCUMu1EN2FvDEclKn/MWjrbKvkDvdUAS3ATYCc
faGPmnqZoauaOy4W6tbu7P5HjCGGrIKa5+SqQ9lW0R4e1auEy5VbjxFOPp8zQxKC
O+vAcRTZmmpcJm1LiNYubvRErfBrqbat9AgN0nuEpasAoVzBohFuoxQn6C8Xs4uD
zc8iYaseqUch87WzQxoU41jJn8Jnkuj342tO8l//4pj0vsocB3MHS6vxxdOY4XiP
3EST80Tu0ZYbtQshHBQsfyoRpdVS/EqdSMBOHDMpVFXdUpgn8z7TX4uXjpvOPk1b
aD07ZcacZRDdvsP9tRdEQBUgULQ+oQvjyVeWpxPmfh999TbZ4kZQ+Q2+/VAboxgk
T9FyF6yzyR7pu2doO/TPsiLJQ1QcuAc1dNF8+KCaqCx6RNQSVLrDipRGWDQt2ask
m2C4QnpakC2S8rwEqzKdwArDbaLWfozB6zqNcEW9Pj4Lsfuhd9TTtelzPr9RSq9g
RaNprYwdWwfUA/usnik1Lm3SuFnLAfKl2I6IVny+wwXVSJ5MhDWR9hRO3VT6R4Kf
lH4gQdOpB6LifcZ6wYnDmjOUO8N6QVUv6TdCmj9/O3PiCyt8vpy4PbVPzp02QRD5
70lU4L+E1rsC1+WEJIVe0s0Z5OL3DZKGA/UETB/WriJPUBY1bShSIq/dc4jflp/Q
pwCLMkaBb8x1QFv9VC3HRl/Wg/UBpRjZ9wzlNAnSZpIYjpM9csE2wpsFgzdCjh0Z
M2w+xxMeTz7ZZINPdsWrWG8ByVf8cOMK+Ien+R+KIPoNHEAuNdLMii/oLWwvemAQ
LiEKm3C2UIj37a511zmWCv9m3hi8VwnLt6VKWeq9MsuR71P5x7grPlyuKJlCEkFN
cn4fSqzyTVoIENiesf+pnBZYUUXdf8DzZhE2oqWFdty3ngchdK82DMj6a4etR7YX
hjoDdvd7zm2j8Er3U5BqagxSXD+3KFTRGTM82xZP7whKIitJiCHY2OaeX4nGhOx1
jdK12Iz7xTHvAADKJKswTnvHzZJo+UtqL+LRsS4Yfc+Ev5kHrt62WQ+wbJULHkue
pVjj3BakS5otCEtZ31twCTMfM7icz6b2Khoz4aIHM5zdqT739AjMIsHTcs5XoXkM
k1HE/pjtnjPDAD9ybDI4Ptx0Ltd3Ugstnh88LmjtdOshdI1jjwYos8a90Y3uFrI4
oTX5ERr6NDxjFvVtwSz56nlL4qWIgG37NU38FerkHDnG0i72iCi8OFAL222yq6Yk
/T8DhAU+QZsTd3BxNSfT/EYrpfBAhZ2/xSwZJHPKVi4M+eZexxzQsyeLBjrFJXRF
8OGORw67piSkNWxEPyZ+6B9crCIE0mrIlKbuzJJi4KpOJ8pgf/9ymjrjCx4/DBwk
smw4Plvq0G7b7LwIO/468rcWj3f5GnOp2N50xlJXAhG9ufNEzafJfjEEfwGmEZdH
njKDS+LCFiLE+e0kUly9tCyvPwZuNqQMsYMxFqBhdmxWHPFebdf9a8Zj/iFIKJLT
TJfMmchtgrCxlHPERgIky1pnxI/RZtyULPcpyTo0E3o7bt5up0Cr6d8OmHGdZJ3C
j1kOiSjx79y8jByAUWGxfN4h6yv4uzieucbPlW1Kc0nxXpcpvXi+XLE0XchSOitB
Kjg1Nsl1CtoUn3NO0K2ucoXvBGm1nCTuFrhidLG3KNJqy9uKq+5/wWKjx2kAHp1Z
cPp6y7tKf5ssZamE00WyMI6GaVEXi4xRo7bFL5iQsaf/xcH4vnpHG7sfgbmIWCCW
YvgTHP2jNA7m0tMyGBwGjwK78MgNgIAgInDoaAQcpeWnri1PVyNiASG2dAh0ZA8O
g0OI4OF2SLkDQ3tjsmeR4ZvLxmBuM66WOAZU64VS0gaNhffj1c7tovHMuRTXMuIZ
x3SfSSyeMytYIJZSLyg/XVwe28SFcIWSzAxNLCGgIbtFBP4f18pgVB1geE61ctfC
+CT4LDIBqZ1WHVyc0a/A9A9lm2I9fc3SrJ+BmEQ35MdPpYeuQeanAUHVxJ9rMYld
D8HFHAbzZixTIyGw01pk/bkx/Gqdj1sUna4MlWuBAvVkIPH2ZP8h/6NHQNPZGKEo
wM4UsEVYPNJqPqLZctync5DUFgQR2SnF4Vyfe5ebjhu8O7UB6CyhCeyd8dzui2Vm
ARdnTpcU4CFeL0R2kjbTi8yvnm6zCQI/fFXPNBSyqPL8PiLTSWQum35C0Uub5v0j
sQFjCK7XzVOpu9wHhFqNPeIaaonwK86pghs+gIWO0WeZlLJvSaih0YOGv1jfJpQo
n8jDRzGnBQNdY8r0uLwxtd3JOQzwqwRzDVMKP4Yk9axlkn8Upi/VGpLy+XPfWqnw
rP80i9qeDl8BZZ3bu2NOlGGIjYmHp2814ESslSZSm7Mw6t63QKN9KRv9BOcBavLs
Y+lYTFdeXBLJXWx1d5tTBBDQU3+WETHFxxcObdHOa53h681ST9M8Cbj8qm4d6kze
s0M5QiDys97C9X5LuPIBSLIG0ud+hLMD0Nv02f+JM7BZQIL0o9tEaOrNMaU2x9kB
zhSnRL4NBzC0HT7YFsLdXN++J4/l0KjtbnhDe6Ot29lIa39tKa0LgwoLvQb56AxR
U/a+qnQ4Q5OadBseHb5lTMrgxIp6211lCoe1g4LabnDScEa16K1qh9P4pCGDyBKj
DXDjaz6SIR1ar5C3ZdhGcRcVJxWbORyitpeN4+HCcEcrNaDQeu4IDfamJ5lR1E/t
vf9EFRKalAOa6pWPnuSPgNdtMPHHxrJzBWbTzoY28+ie31pIhD7QldyykHBeDSCi
7C85LK/xz27kqtLPwf8sOvKqKMcRllV0j7Hn4B8bbOs42PRJviKSHVQeMTvoGR4x
pMiQEg2rd94qkZL+d/WIfcS1qmifYlzAwMleVYUFu1tX2rWbr2Cgg6vFwpg1vdP8
5BsA6uKnqAlC53yPdidCoMgYvt7n4eFCFhQ2cz81fdrDAuF1+PWc8HEFeRgRTXbs
a29/t3Rrt1aWlvbkFYtIwkMImFe3mFm0mYuT+F+HIrm+jfR4bLuAptyCPx1VzAxt
ZZEiyHuSE3aZOsA7lolntFEvEXh2fwXytcSSHY48k5rWilO5QQ9x3dEaz6ZLXm8M
ewAZ45y23ICmiWCJp6N2Q94SVXqcIPzpHS2sIVYeRU4pmCO+9DHHB/Ys/Z8zxLui
NKRCcnEdRyw6qp8+KylhxJgOmeBsSPRyR+VJYfpd2Pw13kkCni9PBwR0BR0THcJC
HOSpO7HmzkT3m5RwNhmHUW64NCCoXnS/d+1J+U5VBQDj8X1KDaDZu+UQ2jf30gPe
KCRDLlCWN0ePfnfleaIwTviKSG0nhJwb17KpDHrUbVB+NY9k72W6CsljtFHpQl3z
7JIN9RMT0kTvQIpur4oiSFuT1gciNTqb47oomwrC2qzd3enYf73DEI+tI2/t4Vb4
OaTv750uLLXD8QfpfyxEH2JayWKmSx2cB0cCR2mtQSIO4U0oXkff9NzkhHpblVkV
c9Xd1Oj/JX/58L+uDCcw2yUTEDmlQS6VjyvqWUafIzh41tuihpAbKDYbh0q0k0yu
Xr3B4PWnheivi6z54OlEYuBB3H/V7RE9RsRqZWVnaI5i8fXPDho/g4lrZo/zmZMv
MT2xxZbh3UWL6Epjopj/sUM17semu1/wBMGvIgdA0up+z7gGIfwvrbqORd2cDjf2
FN7mc41/fcwnu2flp15a3m3u1ZlkiwcBi40jTDnkqqH+nJYFXpZg9Hn78r6N9euU
0A+6p18U/eW98i77MqAoEOcAoQ9my9D+U+gpp2u3mrHrfyeAKktVkJJk1A4tywHV
+jrlZijKIc5i5ZHx1KYgo8xcVjSPiYBrSags38NVkyEBtoXhqUx1kg7lGv6RwicS
NKTCyGzYdSdLxcjZVkA2mj3EMXWK8ffzMA3uLSF9mnAQFswAS7LP507SrpRYMYaJ
txyShiVb/VU8PjnMbvr+DTYzUA/jiZu0SakTH2m44UWmU6nzfS9CCiDWFxCXEZu/
gyxRs99Dy1JmSevfeexRVSRdpbDqkH3KV4W1miJOcct3D0z+LSapyDpkRW7xi2Ja
Q4we6322v5DzeLfDglbimmHKYq5E+RK7IKgiOThVchfZ2eA39NVMdkfiVEEYIH0E
5ysxw2cf4o75xSp0wAhvrdq9H6gJxoMkKQ3IW8r5S931YHMpOr4NvqQntRHvwS+S
AO5m6SRCDIBpEiXQeMoa1vY2M5t2b8fBggHxcome10rs10M+zU8vpBrFAngmic/g
Nu/1HV76IAt9IWqYNCfk8ADo64TTFKTmjI/5sus/tZsFmFRr5XlATAuxAC13kjm8
lW1i455ZaPF2x1LevKygnGigZ2vnH+37D6p/VVKYpb2UCJ6zzk61SHOwwPmtdySJ
iO6Xu1B2UlzVsfvs5SfZMGu1K3zjEsw31gMxj6HLhZd2O8cNRojDHOFcx2M0yd23
9nnep7+tOkWFA7Eu3HXREfEUZf/G8ZJeFcgqrMI253dmfmtjnNiN8yA0YRuMbpBD
BH38ZKczpLVOsdhgYiHQVELRmGXfiEcmg+WhRbfDAzYa7X97VURCKYMDA8rFm7Iw
uIsh02Eu0rY2x5ZPWuisyVRTmsvq6yn2Ti4zLwWIEsLVKmtqvdj2/+XJmT2rRL7J
EHOZiz7oX10PMTkHPikVeY43MIiLqv3QIgpixh2FjuGJawGXI+qw1u1SVO5+m7dx
93dDDLdms84moepoqsrjCBnDBl5OcTyJuZP84kiZUgjYDxPf99IYdZUk8ewkfbm0
PNLX32XyrKrtE4RZgaVvRVg1lEXqS5DNBZHPoNZSDGq4nYp9Xhx6AGSvuhNvWMZ9
mhH813s9T7vMSlvA6f3MF+OQ552Zqg4E9vvQ/bwwZsJeOl4yDlbFEXYDHmGhX/Vm
kkIUDMTIwbk33tD/MUc7oEZLRAIn2izXrp7aI8byh4+wQIXafNS2DBPUdzIt3Sou
i1sFvkF77cTyMJhQuFF+Da9//0RQemXr0L8MrO49SmoJcloB9iNez5ofOBEzGsVr
UEAJR+7rLu1F6mk/zPydyMrjtl1p/8N1FjVT5K+cqt9Vki27Dwc1AwCf2gGUQaKX
7Vj2dk18X7bTg1clhu1QQKQHe1ozk+KHgGn/9zoF3aPvM/IVtoMuU5JajlVBic8/
y2yiGiXRKEuZt0eZ699qGn9CYq+Fu2hY+hPpmOrap4Qyf0VYsUFVw58H8B7095pw
nBE04UXZjFAma3g/reOX68MI7Ph1Uko6nBPSMtlPWhncoUtiTCOUJAfJyqz7HhK3
yvH/7KNJ+4vO97UtXLfSjxBKfdat/AlJOLxIZzbkBe/xwbUwIqNq85V16XmpgZFK
VQRD9F0KXiKVeZnlPzCl9/9H+TL7AjB0KzAVST/u9aBN2MYSYhkecppPEbukP0Kr
D8AXDERuckFApnhleFt5LGXg6BJrcadQIJODTtOZHnFAr75ItBFqFo2raWR4eIaD
O5BAJuHi8NhyzTV5h5Vru1L0l6ZUqanL0DrH/RCRsgGydbSXXW1pFvOT9/VQQq87
V21rdyXguf22yKPgQRdhFb9M/NQRvte1ma/mFa7shCPRFeN2CDYaYl9QjS2ItdLS
ElLHf7JcxDviYd+YYeBjjGUVI2XZxtVFTYzNG19uBmXXt6D7/szO9dQc/9DvXhNa
KZ3MN8zepObWJuqittpM6CgEmIbx0O2LvftIKl0vi96xXMUFYq5wo8bZHVYRziwK
`pragma protect end_protected
