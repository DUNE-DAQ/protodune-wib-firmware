// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VRCbXnPcmnQbk4Lxv8VRaBJ2a2+WjG07BURpM4L1z60UKhODU5wThDL3QUnGo2FD
kcUPJCI0iQXW4HfvtLiaj7DHVNG3/NjoU/3L7pVvOksMH9FvcYJLZ3m0eeVD2pSk
Q73v/XmxbkTNSWAxrXlp+DwBHwb7Mtl/XpjqLE1mVGc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17984)
6V9Mpd8TNzsejuD6qRHaF63WD3gvrOZs1aWtZKL6Piafeub9gfzep4w1300ziSa+
+u8gZIQlZymHNH+pud+bvtIAJqia/A0BdPWaiXVfaM0SRFK3FihxBHBTtd3VO0Lu
ws9hnnNvbnA9zyzXmIx++L4T9xLUPpCgKKUiaATqCxH0aVbPvOtE0si49Vg3rROz
krfJV0yQ9ux4gRJbCklaGTls/8yfIimvkyE2LfdYIZ8lRrpj8jX5kA2QsuC7rX6M
IKAGwJTfQUnPE4qCt7Y01yEPGt+OJjl0OX6f/wapjXB5cmWmaP2GbXAhLwHvw9eN
bo4qkM4JR6LiSAcFaelFDOoxf6pXNH0caEZann9VH7xuCZ02cxRZ85yPKW66Ec/a
/JsuIwDMomNqW8bQnT22H/Nq7vPg57uKl4IvgB8FyXMAh/L1n9kNOcmtuGesILbS
2p15tRzdQEaSgT1dA79/K+mIgFo4eCsm9gc/EJUN/Pcmb2DhynKGBipKt6I/SGuY
Hphagst/vkPB9sHLE+NusUP1NV4L6X+bWxlF2JBPP+6Qo8vgu3Ez2Tj10WuBn7vk
Plp19d5KzhijtzGLS368pcisSMyHlWTW4lxl0VtIRoCibj4YAPUTsM/MDxQKuWKn
8eoE4TaxFGs6SF4X4st5n068yffIL9NQ11G4/g6bM17H+VALdDIHVnafSaHW2Dw4
wqUyYM5W20rPuDvxvvFR4o2FVzK8DPUxJ7z73IzGqVCBAR/gjU8/W5Xru1B18b7Q
meeat/tlCk6UVZOMbXIbBu1IzbeU4kEeipHsPWweY3xtaGuonWgiuBP92LVvdCMF
/Kb8RvbmACX/oElhY5DCQYIL//dl+EvkAhdXR8pexp+htBC+b0L+YpwiDkkqzKsg
D89SCYskePAWdeHixT93dignAJjl6Mzt7lee/6HnrlVIuxTaFsPAkSl1afl/yAeF
bTcri/qX2CGXqtxyvdauMWuoUi2LHGyBt8lLjSsorLJSAZpa+pyojmJ2ept9zv5m
94CxFqm2TOn51k0nlrWk0lbRSPPGSd28gUwsFCovHRRX86hqohU0mOkWXyHz8T69
F/b6ucETbuLKv1CfIICEHIKpOh7WFnlrAzu6oTxLYpP7/c8HkqDG7hYUAdYAg8ax
c+c4rVNJ1JvO2JiWyBONgqWBQND+sovNuHGmZNsDiRQuOyiDz2hqeGKnLL/2yvvg
Ohs5BV70cb2PP5iFLIAy46QluKn9NCAbJilTsYgovwct2OfFBIfqUUgrvpo1Uvki
1syvAEn8WJMn15bcNR0plfqbgowhZBEusiWeMRIufJ5uqEgPAGcQLVFuguZuzC6h
5cj+Gf50J/0R/hFlNVJKh9Bnc8dAWh302JoUL61QZRbFcEGp22mgznwE+VnuESz+
y7THrIpWY1cAVh5/Vjn2gd5eU/a4VzzMRHtR3ArdUWas5pdUaLIrgkIii3m1g/ir
cUoMT6ckWCFtiwNyIPIWQ6mtjXQGRkc2A+0i8vciQMGPSeT+ZgkmS/FUZXijJDdv
P5+unvt2TJzveoAxlJamf6P9TvsIESTT5zW0GBP7d+A4OEtW27yQ1UgsbUof+HKv
ypVSyqEuuwlRhLlutd/wdIyBVrh/ILKf+AHaf+6Jfe1zGecMcjkwRv0R4QVrjtLb
4qokniNWEWFUqhnIYTJLWjBpc+ja+HtjkEF4TqDb1fGVfVcvFcUNw1rlM24I5nfu
MFbFxlpA+fg+uxuypKJtPP6rrSRChiqSBluD744Yd7WGCOsyV6Rh3S8BJYN7R/Bw
S6/9OxQLzc/25NU8rT6cSpJbl/wXKHbKEFl+rmZuog8tT+PVJG6QPKEeDcni9E6B
0F/H0lRawsUKEKyndSAoaJgLc4pakqdHHfi5+2IjJ6Ug1mOYHfQsFueF4WLRUY3s
JI8DYiGxbVtpP1/FOps0fekB/NliJ3D/oVJepi0HC/vyqVC0y4paf4yPR00gtAC9
nPnzeKO/IrjDz9AonZ1lH6X+BrrzhDGWPK2/GuKB9YvLQxgqF1p+s7F+nGjkpjzQ
QsZ2+urnFVLgNPEhVC45jFumxf6ryKWcpn3vsyMI+9xEuvRQkz+QVpVtaz/EFYJS
nf59wdsXbt1QdCD/Q2KQXz56tSlkdyi0T0KWeUmtSwY2lqKLdOA1kU4ucuv1fTpS
N2kDsbRVEveNxoHu/PqFo4qG4nf8VtU1U0ugWkrYt/2iQmV7g03td5Ck3lQwRiOP
vFyhojY8T7DQpZtynotD0GorOTyQ1Ot5wCP7VyDo0CWSLnDUDzO6vALrOXKig9xa
bzYFCmvp3/aDtD4RO7mfY5KJKQZUkKY+/YyXKR2XgJNb/nsYRmhAnOEjFYJkUKd1
tnrbAJrPIr757APXppxds3QN80ZdmxQxGT0GX9qVUG2FDMhJ+o6o0eBL5IZ/SG5E
Dl459M8t6Iv6RDEHIJcN9XR/TFaFrTkOjgNu5ersK3dzdb3XrrrWtbRCs/Q5cLIy
q+Ox/sV/NLeV+SFDthBVUc1q3oKtLWTdVNhMOcwdXVed8bFshWSuTMNchhBS+mN5
edXhh+oiYLXxMv4uowqVCNThBMzC4t+541IafpDwx2IF1OpwzBez/emZT+KhuFMl
p8/34GygLMeLsU89tRYWB+UZ94WIaE3mxftO4s9sPxa3E1o++ftlHY0FQVBHHRdi
6iwRIr+vYsJ0oOYwulSA1AYOXFtESKmpjaANDBH5ASJwFfCk139UwwWJNqbUN9Of
0rSVEF9HGDi+oUwNINZYNQy1gK/qFfga5/iwGN/EWyh2dMRmV+F3jcAGiYPIv7gm
Lp/vl/QpFeoq3ads9DVAmffOIbqvPQf4rSYpsyofE1QBap4qezxAMNoweH6u/POr
+t+69LWbeZyaaX0Nu85n9FVhJs3CuaiN6IhBgLFalF9MSROjImIjRdFnxJNmP5d+
VaDMCJCcw2fLkdtyV6T2SuA3doxHKMznYf5O+cypUUKBcRD/GzHsGOuE9HIP6v3Y
kL5m8lIfQa1loI7nGFZ7/BG/u/J+oBng6okF+o33eQeS+os1X5z19BcBIdMf6Bd+
tMDm099dPT5B9/OZ58pTLtpKhnFIQnmSM8CAeh2WFRB7zlInkxAiTkGxaW0bU9CX
KUREIN/q6vJ8ctQmME18/UoI2RxuD2M0Ga+98ppgOI03RM/h0CZcHJGk4uVTKPEj
U8aefYjPKmy1z63h343k3lHwxHYhPKHCFM5wrZd2packK11VjpY6fBhgfYnI8Hvf
ThXKEhEeQYu5BVGZT/VOoGgY8l2wAU9LtQSAvy921VsXcIkguHbiBNm3ELPnzz77
AWo1C1x+pgVjmOKWRVXBEGfRSipoW5HEapxHObXip14iTeLgycj60erSsnVWoE8q
CCz8qLdOVzLvM7o2Id16zpFkfzqpQ7NyV37dmMkwPG5ulY0y5kuC4Cm+ebFmMPLa
omBx6TVXtKulYhj0Zhfa0XU17PEyN3VdPto3jup7bXPedHyfAE1cfDBSfVSDSud3
TOM8aiEX39vmkwgjk3ms/Cy1c2S1sV0V7M/+hn1FbNI1k30Fs5OSrZzuhqm+smV4
nCPRoAknQshnge0ETbOajOfweP4MvL0BNBdHmdUC+RgMSn/Yh++rbRCUk8J/wB0K
HTBPh+Wdb5+NxTIecazFaGzTyNkwbmNDqhV34WEbdYv65dxjntreO4UrTWDVZjRB
ZQBRJ7qSucv1F+o8L2COoFdWl4zoGia4YPyVQjWgrnh37Ir8Jtb/RRM0IFys01yG
Kja1rqvwYFDQuc1vY65sP92BrkBleAoI5f5dVxN3ik7Cm5lqkEjlTBa/+kY7AczZ
lKHDCHWYPhuQYbgBXPzSj4rSqWbtKZ84P3OdPrygTF0JJ6Z39tEW1Eu3DkH45YAY
yGTetmbchlta2d8v4Xg/htpEWRacla1Y6oulBxFAgSQiTQQw0WRxmovW09/20DXB
vet8rPohywxwUkpYM9OGnT6gCn5w3+7tGLZV4Nuus1ncVqdVUt4GmWp0O570hLJt
QT9v5NsMmrSBiwLsY8p87rCHtC8MrUYAAm474JkMrriJ50LXrXt/h/ppY42yF2qi
Fq1U9Hket5DLTr2FXRVP4hxNcfPsJDKYoEz76J5DfdZxfYh2kdquttAF5jUl94vK
+M6Kd/cEVYLIOhBp5zqj20gAO1KWg2fS+CLea4ya+fgnaEk4pytRmxLT4iXgdfGS
sn+M031xOLQ8QLpNIS1E7I4w1ZgW+faZKxPwxInREBOoyLOnxhOT3d9Zmd+/X2bi
7J6YkzIWHqpNV6Eloa2f/OkTAGjZLpglW91oRsorU+qWj32mAcySqiyHqmir45AS
87V8TqkKNpgTQa2VMkRANNg/uUvA8SDxW6R85FPPx7lD7/wr2XwiPz/Y7W0rvpfs
kmz/PCIWHunjJa4oUewnIm490jK8OxpnPQkZcusXdgxYUxx8h4v3EZMnUAcWFduR
xWhYfDBMNn5eicU4Zr+TL56tplnRRyNMrK6e9Oza9sKv26qQM+MUWpE/GAr/CQ6W
TraZHPYUqPSBooLhjgAFflpQmU2c18d3AxUEgQ3BNyBlKRsN7r7cCFvUnJBVtMGS
aQKUSv9f5KjPg/7a5UWQVQcbcLwBG1v/puVRZa5lrzD4AWrTyRJvobROSFlD2LU4
DBOzqqTNjoMdqj+RxpeJu04ow/ifKt/BI9TX1hAXvOxj303SeW+McUtK/rqT0+SJ
54Iu1YljmNuRn5pejxA5GKFQFaDgUSG1aFsNOstKdTquePOkKn3IbpiQLQOp/8BG
9z5AZDMOhP5PU9cSipU43dKz/cgcnKAkymxjJd6BS1GXGhMyAghwXzjjdcyUEvV+
/pgHA/W4ZQHS4oTEuOWAgEs1AKgEINKaB0lmvQvSQ7Vr4bJlhWl+Kn8CCUNXCYfB
Dpx9/oKGsQ+yw3FVKUg75TazfJFljzwjkNxT8hEyInz1Ml+aLmCd5rSRHGNOzsZn
MtHZSdWpbA3ks8qyhJ9Ti+kRn9GDPN/NecmthwqgkuQabahuM+PCZW+xQy/iVSVs
KMV0l2EPPfsXkh0IyDtGWEsg+XBFVr1U8Y4ji21JqhrliXXeIie48MjXB8M+9eEj
Cbe72nncBsBYNeK1tdB2RTekZjLNN1J25Jyvym27mQooZJ7GwXIqMCG33MLbHDsV
6IPhR6e5yIOwlSTyFkxVQBg9DyPZPRA0Sen7IVW4Zk1LuRT7O6CXzwgrUcEOEWIQ
dAOxEQKmmSTj13aApad7iZrbtnO/BEnwvUaRO4/jAeM/iacLjgqvYXSJnOcPHi3k
+Z7HL/QKYQJJHNMh+7FUWgeza4LGEPu8wMgZtLg/9/zLWSG8K2rWt2bRlCeWL6mj
AFJib4W1KKhVjDVZMDhLQ93k8nKMp11avBwyDR7M4sCxZYJG7B3TUpDs6hviT/QQ
qrCEnPgozQslkpsMI00uI4eZ3U7INMhFMRMTpidzw0y54AGsTGVSv87HWEY5N68t
0B4F7nTor5jkBFonSCU/divaABdzkEIX/UFssQwGFI8oN3yPv0iCoYSTRrK8r8Z+
EjBN4po7xsxDsll9CEFZTjEiIrPEYqYFQ8EvWlYPoH6wJ2AVwv/AWUu5DpAA2obQ
/IdMAtNnSbZlkSTGectRQpAKZVcg0dMdXNZoyPC0WipMwtPE5WOcAKIMeE8Rj28p
votnIsImW3YTExx+uXKfh/lkGndnEACr0Hh1EFmLEczhGSqPoio7F1FtOfR9kfUg
8aIJCg3oI5+Yxhkg6buLG7PJ+aC72n/j292SXf5phLxFnwTW0CHQKiohnjBwriXS
Is7qefoqGozwS9xeP2pfMIMKL1W/3TmPWmXeUMd16tjkrsApFgpkqRQOh1Y1MlbT
OzgzTCQ4iyF+6oar4owYrVNCQU/Mi+vzDRCHwbI0VUwOifpjHPAGXN4xgjNS5aA0
624/M+kUQbUuw9dUQLDocoxjFyBkHrBO5ALLXOkgQ83TBrgiixbXJm2Gs/E9YkyA
BSPquCwZW84xAntNOjh5aX0kaihegrC7eJq3qzF7fHOKyd2L7NcR1Mxyy8FX4f1f
vGJjnqpUbslpfFe4RcUEJqfX0CHvYYj7XRGMiGHihsV8p+QasmUuN5OfGrBh0m1e
E1dmwORlZElENJBX8lggOOSp/i3F8nw+x3wPcvEFKydWJ5b2+/ltf1Y296eqDRH+
OcrMkwVZssWLuXXlb/2Tr47s0Ni/qHlWGTZzE+a1MgyWBlF3TAyrVnsG1XIO9b11
PJVa+2q5fRqWZHxCN2RByY1LeGpdisf5NmLpiU3nQL/dJwxHNRgir6NoKd2cLAdI
sHNHCpq4dL+M9mk7WwEx4YlQjoV72B6O1baC8FEeQqqQQXHCg3TfIS/lUA3yuQIX
MDBn8ROuApFCuZy+8DkAPObqhzHKUn0U5qxCI9Wd4mDP6rob6RXSVTiYFp3HcGS4
xm6nOuakYwnvJh1prbFRLcwT8hcO2jZtP0MNgxZP4eYz4XIteRBe1znCDJyio7yu
i0Shf7lfuPuAYfAQq7Qy0z1GXCh2EaeL2Bgao7hWAMNB1ITWgz1NSgRQit9qjQ2Z
9598wOMHP4XKxo+SzR7lLI2eFAx0d63w5l5kt6AgX5VVTpQ1TmRRM6pLwyRgwg+U
C/RIhYhV24ZZGcYrO0ZNbfNB3FxFFvk68gG7GzI1I8BFt1v/wQbcrbnNkbKJQQNV
Pq6FlX+iV5rzPZbPYq44PVlI1o+Ld5ORVKfZeiBNoYD9KczreR/6CicESBdNa9ZO
zJMfL5VZKLshhShjtQqRG+DYQX9ankXfo79ON0AG96dT5nyhyHc4mxwZMHp/MDRg
wYIkP8T6SV5CHbOsYjYvQ38BBKJR86ug3uRy1QsWEsWnep8YmddUe09WCC8Ac8Tw
qJQq7n/taCZlQJzB9ElDSioAXsAahBwpJKHnvpT28+fv06NpZFi8mUsNzcekg6MC
WawCi/J336ABw7vlFvi88uYyE2jRL86k8T1bfdFTeDQdNokqJ11n3JqKTs7ZTzL+
P+T3qNF8WQjIl8cj2VB9YUSm8Er8ZcgHvSHHhA1ByJz8vahAJTBUHigI3twIQ1/L
VHHfGiYfvIJPz/efT24I4JlhM6zZM5BKLnpbn8qbHiTNW7j2X2t46jvvmjcLu8Pf
dxFWgT4BAvTgHx6oUWg17LLrHal5S8guhF8x6BUzqgp1IbeX78dXc28LHlhHVv0A
wq1sqoakwLkcmS8rYz7FadjO+ZZ3ZAb2HOe46LlnAFICO9Hh41G6Ntkp4UiOMWwJ
3jrAl/goWciSzYS/gVITsdZBw3/a4ZCcZG62YQw+oICZ3QOeWEW6pJDJYcB2eSIf
ZHYbLiQpeUX26F/7UvVENBZpjv2daYBD6ukqn6/zvQbJ+YpStYOIUer/3mc6qluq
ZwSMINpEXjoS/IGklKUx1wdwwl+oIzgBysrKfTku5e3qj1oq4QvIfc+bqyuXJBMw
lc8CLbbuqDzR55ibB+jY1bAvsI2JfUody1n16CtvUXsrHHDdFtIh7VANF2DBKsXx
MA/sYBB+qdpQWq+L/I4yqB+FzKeEH8zgN6BsFrmOE+vis+P6JB6zvaI47Ph/cedJ
kDraSU+MtZIYjKU7q5tMGi6RszJ/RybXaBoXTxw4vZrUHci7mVMmPC1ldxBAgbbC
VEziURz9q1l6KxWDa8d9T4J0ZF4uZ/Q0vluYU9KSdQ29Xi0MVIzx/AorY/uPuvxR
209pURuCpamZik07eccCmFFDC8VpVsElaKjOoxazNPlPkd4mayczfRTt7JXf6vuu
LUrvdj7qkv/8CqWZ0lqK2kjbBLu21yQ6/z9oEdhXDTJMDai03sIw+WkV5PCkwPhS
pMlENktErMjwllpIOWgdbef/Ffh0pgIkRqo8ze/9gvrdydGnErYTy1/Thfd/b3E0
LJqp/oE12PkDPXOCY+qMczibL4z8bXd8UiEmu8hwkNJM5S5Fwx5sc10HUCJSr3tI
34HPsDa0KLm6JiF6b+VZeGFQCK5m++uUsaTVpurj+KFgB9vDHEUveTSb5wCWfCfi
3wkAF2SOrqPMNhSzJbgYmXHC0EITcqwuyMfVCJKIBkxgG5MUp+l8zptlrI4R0i0T
6KtajcOnaf3hMT/AbyLZoMtwgvT0fDFeMJ5c7bOpv7I9Dei2mm7Jrp1OQTrIyGUr
IgJ+42yeDfsuZf1f+REt/DSixw27Y+P/DI/4fFTgh4hfA3IkU8225u8JBcncGTjW
0kwtMUT0kSkGwGmqAuhTLLHijdgjwralJZErdf83edWKcC6nS7hokCzVu7mLIfnD
3DCHBihg9lRDYLNVRNCWa2WadxCbCvCSPob11ur6f+WJe54mM3NUHhpgXizOeyeg
AK81Etg2ddChez3izAVHtWntQ6urSo9NjEjY/vA99yfbL5dg1t57XkxptB8CZuyq
S6NWB4SsOEQfrj7UOdNKpVmi0d/b3YI6C6tnU1x57FCR8b+d+pKI0vK8adYZGsrO
/i801hoNBK/PllOCr1nucy4WCJSRzfMzh77I4fZ9fJHGjGjFsx8Z+p0yibXYL8OP
u4ajd/TsX7edd2WqrIfRogkCMAQbVEx4lSUoNceUpNHm2Ozj8B6VsH9sjbIcQqo4
xCgkCTKhBhKRv0YGpPEWrK19dY0WqMQFDFadkQDzVm1/Cch0bFbSVUIyBFQdTtEh
wHcDLU9fFcjNFwbBRATXnHMCsry35B6cgo5I8TJwSE6W2/ytMu8HjVgdZRm3ENVK
GUUrEzMk/gAWSXKdt2XF4U06xBsm1j+UmgV4qXd/CQxIHdQ2/AmBNSrDyv7bPqX6
UWTLLtefy+M3WWDM0ctbadXi9s7GKj5nvYsQmd48qaQyABJPoGLChFLE1KKRjikh
fU2V32wQ26QvcZOP1ucE5Bqjck0C4LLQfNA+B8BLXdT4aXcKj5WGjh8dmuS9Y00Y
DvUEx4xaBQc3VlaH3kmCuPIuuyTZE6X3VzeXlTBCVtysgsUWaD2I1fkn14x7bVUZ
L5Yv4EAPvF5s1ZCgGuNF2GR7P2NlhXCboH/bENvn3k1DFRXaZOFflUl6iGaXe5MP
UTlvT5PkRjuLHbcn9EOLRwrHwrX4hEzTlgNjMKpFs0KZb3PSONjz8MhW3yUJ0E5e
6h3dyxTSLOv9W6Iv4MGMcEDNLjzoxgcH6yBcAY2mcRPGP4JErF22hN0aNmpfAveR
SZpnvKFpGl+elWbyl0POQcsxsVUaoI5LLcHXxv1B1hQW2APoufPtaId0+6YAPjON
GpUkgWK+R2coPiY8psCTHJsiitFIyxJUIZCVPgpnHrLE5OvawpBCKiqGjAtH9BVB
gmluRbeMAYGBsLmymCz4Yoj076aRkngP2jh6sgREnpZzoyMAbDRzLfEaRJTi3z1G
5NHGG568ecjIyuUz2JaZn1U10d1S6EFuHu1tbEeORnTXSU/vwx8WiSPSJ0vFEuD3
sykQA1GztNKDl/idi/KHjubfRyP2OxpNd1oD0czRK2gugn5f8AsrYX0o6NkHIgpX
iWLG0z7h6B50+uaJZvDXSIQ+v253Wyb6piU3Y5d3zsJzX+9acDL2U4LQcV/xlSKY
1x18nMbUFVm/QaWRirS/X/hrKLPHqvS1LpVakctbK9sagpugJUjkqBxWPuBDLHSC
E7aAsFEXwZwMnu2R4Y3hNDoiPuHsN0ljDTjOeU8BB638g0Nfj+MxF/0Ko1cgxcLY
EM5m5LvbHdz33k2SIytsKrykSZ7HtkV/gWIr0cB2VDinjwa4xNl1ouiZx96nhx30
QaDLFROCAPA5/vYX/kH/6LiU1dpxgopzZJ6HdjPC3pivuqbaF1Lkyxcvd+UOKRPL
EUJICpc+dcsUEInNewvF4+yRCh/FjQuTPBy1yLighUYXQrKjiOgCaACivxT06uVp
lPtOL+Jp0J03UyciUX67tXTHXdWnMvgciVgHL8NnjARUZs1JbN3RXJJoqLRd1CGG
EgKQ7sYQ/yNrA7kh8OO/F88TJO2ikqioArGHtLskvn292FE3qgAjpxfwXNw1Zrra
9nnSt5fVS9J2LKLmyf8umwTReZ9jKqOukLCj7ZWKSpYal1Yv4V+C6sv+fKVBjnza
rRuWZMDhXCFVDkgERcLtVpJ72gci7/hu20W9k6EyaJUCO5p6Ii6ioNkUJbbB36yY
uRTzmyqLXIL5jMoa3Szp+IdydtdQ91jGY39p16CbnMe+DdYhAgYd8r8FcpVh5fPA
WnT+r9DX3yY+q2zaLTXw0c5i/KNjoJkEGTkzgyB5GIXHw7SNTc4cdiV5iUwaRp+e
Ve5b5vjeRndfulhCyvQQ8VkmWm+XKOvWluuK1iUc9GsKa7HeZFrn1WV0BlhnpgP1
nQddAY5GLxehsHnGw9UcCpcNjQ1Tc15QL+/1n6/UzrIhIl66iy6dagBjFJFv0Mf+
9ShuHiL+X7EZo0xZhkkVnEW/6nj6KiYTz074t6zPBtPSUvNTBF9raRaADRyXuRRE
NgWsuAe9jny5fGi85L0qesRx9E19ShBQweCTGUHoTEF0cWeriwWgM1KFuPJmbaev
jV+rfBDeAFm17rrYd7UBWjrmC0YV8aUSzvjomOohz3PlMgoExA6pdiYTI3Ap/J7h
32YDjsQfWUDLuDLtCEbxGH/Tr9/vxedlermpXrp5n8jD8kPbRgpk7nuCqV3FjEqf
2uZkrJjp9H7CxBmJIbKyFazNp6NRKWyv7piNkIOy1GaWSavDcVa0JAC3GMSXtJQ1
KAIEwGFI+mq8kU9ZizaRgAyBVqfRMVLR97LLSN1p/6skiGXCU1TLsgCUSMYrrtBK
YEFpMtkKIJtmfemoQ1ouDcy5BceIk2Posyh6xNqnAjFE0sWjijpSsA3GHcOfCtHE
MxIGcn0+9+ZLklKYea92fCtfsqjb10Rpy9SB7lTpeMF8sbSHidEqOeytHX9USuKO
SHP8LILNwPvNN+MCVSceLJoeugspfGugu2yXQx3BJwZlpZyLKOsoq0at9F02/Qs1
ZNVVLfowZ3TbESkwdp1WtzyoptRTdAWvg1xheSGlFZXEcysbZkh79+YmyA2zWDP5
eQbFsoQjVJxzYvOfvze0B/OW7vYi5mfwAWI6leB8QUTIfpr5iWFvCYeBLbxGZiQN
EzhustnjwXspPeZ4FioFz/pUoaYrMLSYPFHAAO45HZP9IKVhAVSxy8H9pT7L06Vz
7i6O+alOF6T9BRrYjw21sSFnxyQBzOYpe0nIwyBBVxRIS1k+awSeAI3Hkb/rDGYk
rslTozzMUTutii+cYnD/JHaGSiPyW10sy7nUx+Khjv9CqXubHqyDm6bTtPTSCNbv
HOcw9VpiaBqqmW+ukC5/cm4m3G6btWqiC5j55lrKxuMXuewGqL0DM21VDmmZ3xQZ
/UDCcEMurwTZXE/u9JiVDb1SPG9bLSV1OSXWXSlBYyk9lK0G0fmkfkq61jk1UzSQ
zjpJA1NtyzSAUxbpcN5b+AXa1hnhxXeU/GO/QPpK+Y0pY6fnSk+9IKUSXCD3/PVG
B9c6b62phOZIE+v2km6kzJJl/jwbzjDrdFs8xOeG4k86yhIC2gQWtmkxRloDt6+e
sClZd9TYywMp7VVsMoWp88RT4PDxTmfEcKysM7S9VmkE5gPkAklp45WhTLNKdsrJ
yfcxrrnPtA1FBYbxGoV3/Zc3Wmz3fw8IqTkIMbJQOsugve9HO0aQl1yoIvxqoePC
Crnt2jAK0eMVQAE2VksZHQTPwcufbY33R+vcMdJYUKe4ma3bMvzCszoTXRREDMf/
fwtHv8QKEA9e7lQC0fq9bIozAPU45QLztAfGzW53PjItSqOGLU2y3BKJU6avQUnj
4QJHI3zhFi4nj3qF05FAq8TfVcl/ymKkpjIZ7hjg8zWY3qGU0xp2kpC0JjZjVhIE
iClYDyyyg4zB95oSGMctkk/cR/Rt3VCwp6z/PiJU/NKtSwopZMDoZOj/NJhzCd2d
QlkTKjmmLT7z5qtq2powrG8pjH/+WFD0YEK2/UPsFEN1Gs3EsZOqF1qpA0mK6+aK
Wi8k6TKibHFeDp6cX91JA51+8351o57t8JfIuQU+mupGPe15/e6OlFe9t9f74b8a
thI/F4O1fxQm6RFkXjmiYajt1l07F64unxD4Fva9QDHh1cguiYTCUsC0LQ731Wep
D4JsjsRAGnnVz/7wbwrwCWcKw4Fv8yMObSQeZoliQSUYAWkmRzU+h4kST2xJokMD
HhhM26sZZOmu8IM9UC+PyGCNxD4gEXzqLLGT95T7JO/4bQZzmLbILJimk3P/Fnc1
ZKgsAQ2MyQgFVA3z5fTeEBiRzzLQeViZWUMW0PGw/ZHtGUX3o7Nfl/hPU7xs/NE2
yxVSsYwGBKNPwUj2MCyxzPLPivj4XEKBmM8ioDUkskoz3zAvBNTAwBAwOF0T1anI
LLjMFBh/f81G4KScsUiK2ZgVGCyAnHbVTmgBIh8LnDsrieMCDnpg+fr0i2mtWLRw
1tCwB7PYhLJXhlj06gmdxnvZo+SaoktNWqY29o+NsW/SMq8aKWuMCqcyOLOthXdL
Hj15jNvUZaZ5vXLdv/cJl/8mUMApuTqpGGgLRWsUoCZImUaWJ60vYFf4lX5BqfBp
MXknTY3SltCKHK5bXHACteeJk3TTOnU9pZTGNChDKGz9a7yXfU6cL8NKvFsIHoO6
anCKlnkFYkKCII4w4FpGpHXSblzwgUBzPpl7g8mV8NGEm6JdgcPe5GEzqeRAEwg4
fI6mRdrBESZEEllTLzQjTBfxlwmrvg+vwm7u2NSU/7xyJwHnjRU1b1uEMcn56JLl
BwAJ5bgeitapB9bp7MDytbWwclcuqbT2f7X/Rci1/1QmPfaGRyl+ie/iLaCxmZrq
m6JkCFoTeT/DDBi+JcVXojl9Da9K2XLOjyjhoMEij+X46PBnDP3DX+d9a+VInaHm
oEI+iyBbqxWatp+u8g782rF2XgSFGLtVeRM5/1sYABvB06WbmFwYy+mzsVk01sFb
YXfgWB4OdCsQDxFzT7sN0pMXlVqsSiyPTpkmBETMRR6itG+PCnk2nTjEyq8t9yjU
nvI0XK+E8SwebQec95FIfpAWGI1UmM6IBwm9Q672YQDN8rQKXNk6wfqpEsXSRN3u
nkCVuE7c2kvDPJ3JAlgz06PTNgRmAExr00rr9JQT5PZzcRMWfT9aonSDA6TUcvZl
MbKOlTYlGUU6ITy0nubF+E0jIaCTBFn8xMGpli0QxIwICofgb7qncHjYxLa0HuQq
YjrJHjydaXhge2tSQBQiwX61XTvr62PMraqWrE1VO0mT8XfP6Ahdi9hw3AxrZNal
0gQoYag49hjQjWLpPX+ziei6PH1mvRHKPNxeZy7u7Il72vmRMXYtuOOPM5i4JTFT
0av+fcSG5dzU/59mG8+46EL8UriujaxTAz+wkV2GSnfPZhK2zDWr7Vqovmi7PCi3
3t2i7uEINpYKSFivTFiiNNUZrx7sZMHhkMBtl8wNHuW1xKnqznjkC+Gc8MAaRXK1
5HAn8swafo2sASoIxuHQ4FXst6DBj00lXUsCnBoUZh6WqORUCe+6a50nOkXc9Joy
4nIzuFXdvtN5rxYMpi+4VGFnEYkt3jgurKjnI+ggfsP39Hd++7Pdz3BFzx2IBxyG
n5OQQak/N7VAgDY9j5RMisQA92gBvRh5pQqwOS3PYnxlXzGyUABVFoUYMd3Ko8XJ
uuBUOtwVl28q+dve9totqYG19/gX3Mg3+V4pDVaU5kp+UAZcNWs4H7do7pIeyxaE
xIBe0fzmvvR0GT9zAocJOjBHjpwlGyv1u9HPOz1pUR9UVNfF7Jt8JvIbDn4jN5U8
uGSKhmPk7s0pbMx8P6bgp5GMgweD8iQqJTOVqGuuZmGEv2k//UjG/yhM1VpMWbQq
Lp0oQzftAvbgyFZ75D4ygupMb3dHEuKe/CaR566xfmy3hrUNH275rOHqNQOAhcGS
88a8nCuUepaqo6rBXxyLK/v75rGkMGnEdIILzjFo8QXQ6LHZoQhMJMhYqnP6P1eq
2TJ2G194819+jo0lTBI2kIWZyVYMuE0zvn/MgtQbBYbw3ri2hJ/Q65GOhPo7xI5f
DSRQwDUfd3YghRzXT3FsZQpAMVJCuPvEjdvVPxzk1Z80nu0IDRDnCm/KP4UirO1m
GFUeBfkfWvrEsfmtspYaT5ugYWA6ImUqzskRHaBM/fJ9jG6lfxTYOzwVE9m2sOZn
OU5CGJPWKwr+dwiBU7H/A6V2v9YOO+EMP5lGyzLDgaWTSi9QY3MKoC9qI/OAd8OO
8n1fHCwCnplDlcyE7HSq/x7PurlRXWIHYBlEhNClNrfJhtgCwkt/q1QOjfHoezZy
1FXrp9wV4pqMnuWu6Q+tDGDqx2WT4KwyB0GKqB5h6h+Cuqe1iRyPKyIca4vSjCu8
kVIbelLc/07jYUTxQJ6RQAP65GsNm8GUT6VoZm1zLRF3ZYT612Axq/37zuGJtzzl
y5yyJNon336FyfW8RLzQYDrT0XYS4UIgnMG9OMI57N4dqSVZM4HR3EAxYUX03saG
CkgDZifYEHKWMNc8+F8iDU4N6Tlfy92qnNElWLM0bRnehCPLgWVyLQFtSaZNUTaO
Ko7Kbw2Hs7fKLVaR+v6bgwuVEpW6BBX/9VmfUD21O0tcHfRzFpCQWNf7un+XdMPR
XdYj+ReIXy05USOyM1ejrlFX/32o5ZXd7kn5cL/d5IuUDFhAnFzdlgeBTKtQVPrN
y3JLYOwK4YnAQdrRONV2f3E8Apy6jKTGFxmpIaRlRhT5CsRUm3Q0BgIq3lnivsmY
Cz/xm3HzvVUslRUSvMv8dscJO0YLqjNwFEpuiqtSZ9dYBHAk3yVAE7iFUov5Wee0
Xj34fdav1UD+86Ye9WCpe3OR4hxDfBCXy8GmTbClVYvlMfocPfeOgpOktpcMOD6z
zFAfBXbWWFHjvo0DLAlGwPn/vAwSb3qEEoYyfHGOAIvvLU5euvRl3x5MsKnNcxur
bcTbmZhmd8alBtfFhqbu6/6U9KatdsHIFqkZRjLN5YUqzij/3NTSGAdKOY4UIHv+
nwSTVSRkuU/JOoIbSog6Lj5E22EF+sEVjWgHWSKoqmIdZpO5ooQzlfX4FaDHDC6V
d2xwd23V1Bi9X3kmoDysD7dvamVOukCVQt+/9wvOLN8phmvoE6lHz3AgfBFak+MM
JX0qfWnm6hN+R+X3Ts9zt4ywFs92bMlhXnknYD4sXd6YWVpSZkVODJ/19ZQumkHo
DxkYFZ+J9SJvd7YT/eYe8b2x2H6p/gb81WlXV53t+yrafuhieiSFqCxqCL997Ai7
V6WDcJRFNWRwVA/+5ZmtSXAlPLWQ0V9KDEtDA2JnCo6cVapC81akWYl1RAvNt8XS
Wc8NMuDR5DBAsL7DyemW6rq0QfFZWW+iTDRyj/kMMkPsFdCpc+oKqu+LmVI4aRfD
QH4oDhVHuuE1DZzHhErA7urKVJrX7H80d52bcMY7l7ny+0ed0J8jlSSLG4x9FP+n
oXwouOi/PRMzCYBOmRqy0VpEzvAsotttThz5LCZC2gUAraef9PHm/KjPDkyGjEv1
TOJKTUKHuvw4856JriUMJKO/dBVl1gIIcBCsUg39VAQqBbg/wvT+x9PmbgdHJV/8
gUVafmdYe4RHZWApDrHhrx8RzwFEZnDRzo1S+ILyUw9/ycLxWQtC+IbbZkB6amCo
PkgocJ+jI6R2qZr3VcobI1DoKQtBOc/hHPogPA1mul2GPhxVDuwoVKnmasbBoSHk
zx/qXJV+Nz22TpXtpBZZvtcFeR7cMbfy4qeVOSa0uovCX25+3AqAbJq4DuXfyJXO
Kkd2bbW+dvB5Yh8UeEAE74Wk2t5Hz3Jcz4CKVHGt/NOCFmNZ9ab4yz99WDIYLmSs
KqON2gS3w/CmKI6o9g+JZ+Uli0s6+hdixj9Y/JUfW4VC1GQh/jfBGnWv9iF1YQ+q
E02lKmt4Keu/PugnIeEF7Qhk8yKxIBYSvn2jRIVM5DRmS3BGaJtueC6yHfdlYSn8
tqqc3sto/UWoOWD5ocHCepUvu5AO3OtyVKXm6zJa6wX2yaYessdO4kXxi/Iht1+r
eCfeIk6f5X06YcLdFP6OOA/b7S44XdawlemO9dYLqiaTV2hsfjRj7JuYt0LG07aP
7HAN6IuiXJW/tJe9bmFIg1x1yt3mkGOOZ5xPkFxwU8n5OHF3tohBMY5X07H0atqN
t/sW9UojS9yg2iL0oLWkSQTAAT9rnlLnOiUWlC1g4cu/GB7+FvmqR5gkBgYkWteN
oDttCQdY+TV+03t/RSjXVNDY96Z+UA/w2bMc/Q5p5NdZb3cVrwpVaRj7cnYPcsFG
XCtnpLPv25KdooGVjhEQowgp3+K6uTLmEzEUPf8SSPXK41avtr1dWVwfa9IDfvmL
uyId7Np3bIgc9XY8SG4iUNotqXuMTT90jgf069OYcmsGi5wcrElegHr5kUlYrCTX
BoGwlaoWyrq2KwyivkB7fySY5fDU990YtUY2d5xw+txzfWGjPl0N0h8D+SCM4GbN
aWKhRslX9nMMNjWWVFrBEcCo2/+M3jSFO+gzzqJ/etd/afzbbTPDJJ3JqzIJ/412
qmgjLUJ9kywcEzE+nFN1iIL7oCrqS3FX7VJa7igcdzalGbN6q+2do++y9OqpY7tc
qCl0Wzwv/kFa5skhLNHigcapCGp9CzhWpAMsoIHLySOFIgyWedbW7yZ4K0euc9+g
f2lioZNjB3xRlrBfsSHmWnbAVsAFWkKpWAIV9pTtavKmG0vfaiRpmBTdOMQjoF2L
pNewkjz7iwu/afwG91UyrlZfVuyVzGD+yt+KIQHX5wKU5RFX2ORba5TKkhTeOCgZ
hZonJuH+1D7WoucxycJTNYH8kci5YZDIrc6pEi3ihHyDpa/P37VOhZDuGN0fhWcu
lhHWDxLWtQMJkzMsPWUrkda1kNQX3v3jFoR3LTJo1EEiyah/eyLxmbSa+y28iRDX
RG5IGAT5KWsT0/Fz1svSvM/NCMSanLjIQljMjnH5wrzWcpQvxJ6fCV9OgUr7tKWZ
euHr+5Z5C9tnF3viQN3tKMxO8IHCR4pa9GwXoCAYGNBIkkIN48qS/L2dvrVSAfW2
MHhrJwl53oreWZMUD/ZMYZGmK5Vk4ZWQ8HUt0pPAOVj7mHm/tReMcN9oebH6wCpo
YJtyyyqQXqH6cvCFLzS4WAAZOfJkuwXfr1TMLUPBFs4WX7geDuZgywzqulxo36TN
KJAJ6Cgcm8+q1SUtbIBnL/120TiGMOzfXzszZTktxAKivN+w6UesPEblfLy7eW0B
EEzOG9iab7k2ihzXQBKPkSjC+kkCE0wJZ3K8I0ynSOOtjo0lFrN3O23ukGpaTOmr
8Ug5NKmoAN/6yX9rIwl6GCfcWTkM8+/i4af+z2MaXuTYLWOFhkk0fUFS9M8V+iOm
YgMXCppnKNSgG+K1pYyn5M7V7eA+cESGsZ2Kpt7nsW0ER3nEGLNoM099D+CX6xjZ
AsqlEiQ/HrfdnrNH6NV+/oXepb2rJZjVE37l6+aQ3dpugASu+aO0jxOEeTFKM6C4
y+Uv1dZ6czxar037NTBFNCL6y7pz8fvsMH05d/6fAhp1m9uN8b6C+CXYCwWIxnKS
IHSQyWBgBtbKsR/aDhJU2p8rPSi1jFvbtKNBa0+eIX5IpYcwNuvCcyWXxUPBxbMj
+U4CMZ22/kB49oy9/Uye4W8g0w59pcrIA8bnJVEHf+7GbvHPtLndA7HZOn/FVWHR
X6bkXUSj3QF+DFSzHH3XGrvut9IjKmGvJz1cOydvAH2ADHCZe29H1QGBucc6lQ8F
uHfPrxuVjeCb9b+E6PwdimU24guRkU1cgmnuMHDhpb7YSyIJQEJh7Nl1/Cq+DgPw
HlKzhL8KHpR2RrEiZ4VICLNQVDJr1QflgEH6ae4yJf47zD0aqWe//qoN3NXHdKXK
qWIhrWV8ysc+NDpPWCCGRvx++MB/f8UAP/U1y/5ZD7r2BYJBFqvc+BXHwi4aHabw
JLPFdvCZvi++m2/dyIzEtwXryWYoAE3WgvqP6LratTmlCZOj/l3NOtPXzifPeMF5
QinpJliZGOwKhitqx9W30IiQNkPtyotgz92U5fIhKGqRN/EqKZSXtVYmzsGI1w7f
luJPyxz9wdQwPoJrvu8znc87p9uJxxrHg3/r72xYZ0TeITdNT+UZGAU98pBi2X27
rDQSsCSWBcHCd+D4JWHdkfvXWgOGqbn2wc0hcjPwkfe0tnSdCPpCuEMnxCEMwxEO
69Nugj2HbZIluNEZA2cO6QDiaat6d0pH/Eu78Oq4s/9AVJSiJhGN3loyXEj3d5Dn
+Rw0QihLWipH3N2iM2/hNYv9k1fHaYXx07CnImn41pBasgb5NGSwWqJfzB5s5VZ9
+ldMws4/VVO7DLifvwwScSL2qEg9zZx4+Hlq63iAeOrjo+vshBoONkEH4hCz/h0c
2shZdFP5SbHb+JYf/Dawv70/i+0G6BCJ7J8FNgIPONmTpmbAv8QhfJ7Auv3U2UDC
ZaU4BKixE9ifItedhITy20/AqXDEOVL9e8/YHMvgtQFzdMjVEQ2Fd2FfUGu2r17k
ymbjJ7KfQyZQhlpiuH0tNYQAjzLSYhaW5SyerWDuWfjBdCFFtWcnNMecsiH0lcuS
LbfjwlO9GR+g/WFcmTCJJIxeUsJxiq+f3MYgfNSJoLxOg5De1mEo5VA5m++OraI8
SNKlktAdRPr39dWJAvbierJ11tA5ODwHtj/l79+a7Jjd8aeFPLx6elCsrW18JHpl
gbx1pZHH0X5T6WZDaXKe8ANIl7jGae1Ckp0bOhqNk+x0SU8XvLSbfI+TnQsxvvi0
JIlhdNFk+c1HEXA4RzE+awfmay+PrUQ7tCpy/oE4B6/DA8z2TKY8n+N9AjqjBfRe
eTvUs1Ob2ntsiraM+8tpv6Z9z2H4GtfdJK1vBfjt5x6SHgoIDyJ6tY9H8C89xRb5
IQCP9rEpONYPnkoE/wdncoOI79jVNEzOxWFvRAfWnVqDT9oYKRp8qPHg6xN/kDzU
KarbF0NavPQ1rb+4jMhvO0qhlxkji83uncCNei+tUre99C7X7NLNR8X325LUcGK6
wKcQ3cw3DWsGpC5xGyWbopQlm+pCOHqSOFyVTEZ+RXI8yHqNAcZr7D0DiIAs4F5u
3f09Ff4xts8f0csDk0piDP8PI7oAxvYSZGrbWlm3jflcgreJ1+X61PdOFi1YIWqT
/zMPMUSKxI7N8WAmje/UupERNdAg8E1ZTt4TRX4fdPo0b/wnPgYKTUYur9Jzjr3U
5OhDlDPz4k1WT0U/eoP8SR7dTnhBpcoBIiqXK4uWBN+jQDIWa9y4CPYWdzoU4QTh
m/t8NScCdKPV7rkiP9YttdEhVnM6571cBt7L7Obrr/Z4Hn/jnQyzABi+3JB2dQLJ
lmfR5RQ4ozSgX+2jns6w2G/ZEpXRA/G5gTy5DkFGsmyEdqOGwAbal75mNq+qDZE5
NICUGNVC7I8KULflXCdENss+p2rKZniNWsMbvgJCVaCtvojOIRmJNI7Re1307VPA
A+Vw+6dXPR8kEcE08oLxhugiNvOzpVtrg7l+aL8v+m4XDZajbroywfzjozCsKDXl
pj/p4b33TxYmoVTGJHAeCwuDX6564+WWPa7y5GWS/CdENZ9WD9cZuipXAdrZiirD
ZHcoi5sEJjOOqhr06yDHntU64LDpzgo2Kg6c5oxAkhm6q8lNek/lIHbd2QpiVMsX
bNxP2N29mA9IHksQh8vSIpEuvah58b3MnoEiW1Ta8/91A+WSC2ozA3CShcIYR2kq
3L7Re6oO8mGhhmKC97dEyIhtwhQACjh0QI709SUlo5wVGKn+lGnhFDtGvraqPNCN
fAelWopCwz07d0Qo468NGn50tHXQ0zNwGCiOjn+T8xQN4oKZ6/lsLSzDDeL/hHhX
pyQ/WrTVlpcwPmBLSLwSLW7JQu8f9X2EHE1yu80NEjxRbe7Lmmt8qlhnCTHgasDO
f2SdtfPY49lzxJPEpxmlGRyk2+v9qDsU4kCaA6GweJP5gGerRYJnSSSypZqffCPM
mma+3OpmcSastWIaAC/r2jtmLi2uMXtBlZg0q2HpplZJZnMcFG5WdkPeK/6qRvpk
XzHRR/TOzVUZe5vyJPJyZSGIj5Iso65iJ3DL99pOU6oyY0Aq8bo1JGGDW3ARLRAI
oC4kHrclwGjmzN0P7chXnRNmZuCjjqmj5CymRawb9+GzUghwtfi69uY1BJnEvZ8U
0lpA69vBdzBHQVYO8NaDUV9vhB/8H3g4peF/d+vdOXpHvF/Sn37pEzpS+4WywQq5
ioMVi7VOvjNinDr/efHW83DRPS+k/wmMW8Bk19A2t7V20lz1nQcEbskMbf4u6z1D
FYaLuP/tKXAfavvP+o3UnY3mIKRxg2b/XlyQMR4oWqDBHAooChTAaMPbtvtyLuEw
Dl/hZLNxHumKJb4OImyzanoQUEnX7aQmav0uJxO6N7pRKhbws1DrQOSTtivPAlo+
IaBguIwzecXcupMMVcBJNeLVdtARju0lS0RISIkSru1WCkus+YTBJ3hI2LBVadZT
tFA3ZDy6FfW3q31b6oPmPO5HuUljKkiIcucDGjpExfV7EIfEZDhZrmv3Mwps6Rh3
1UrwekOkAnm0+hLmot6JQTVmVLxDdqxHJIqup3hBNQ9eSmZLFDZ7xpMWmgiVkGjj
q8kCQ57yWczs2id6SZieNqFAKYzp6OK0MOXATCIl7qWpz+CTgHwe/ghwP7f9So6b
24BSItyAhx/m0iVFAGWBXgmzVRfcTGsNqc1UfMFVKGM1nnsytxjUR8/nwMCjLvnx
glh4/02H7/6bLsgiDEFopWrwOOvKz2ueVy0EmzOsdVi2y98lxFdp5fQf5RSBe4oM
SqVeYU6vkEBh34u1DqU9K69uq0TxdBUgeoGFWeB74dE+wumpbvi98vAdCBsoT7oZ
oDa6C1nvxkfeFncAooxjRqSWm2R2S3GDQPO67jtyWpCe551Yw+HAr4iAyCVCiLc7
gX9yM2yLe+K4FB1hfMFcpmxyVfd1HEx7+/bNe5NuQnS7DiCsarHYTAmbKL47zH84
AaGPbVi2VEuLrSA2zJDaO9akiUjngbYkt/bFnkMh5scD8q07xJj4UlJ7GL9hUget
7mr7YEAvnAhUrX4PpBgzkXMg24sX70gHYJNRLlOZCJ41uvqW5iG5dpCXYjuFN7dM
cWurq+Mdc7j5DL5tOY9e5skHGwqVTYpoeL2kViHDSSvyWunowIdvnp1KvtKYVJ9+
U9702O4703tcuFVrm2R+HS0Era1IMGUDOGUgJOFm9xadYqSUh4USX3eUdtZNn2Hs
z41pRSaMz1g/cMg4+1gzMcBrAfHM6lDJE6Qi3nrC0139fiYpjLvWGwb3lbP/PXsy
Mohra2kpUHU99RjFAAi0ms83fRMt74E/n3jDMMfkfzPg6D0kiLURalE84iDGsoII
QI3duxfYpKhwmExMFUJlUvr39U6DM1MIoSuQMHM8Yc0RHSo8kTCjF6nVC7Qk76sy
3iweNgy2HhO5o5Re3nBloDrIfSCUvaUb7dba3TY3XUEPfBaJLEXCMv4Iyny4/g50
+YnT1WPKpTbNh+W5ry0+W4rs77EG84peeRKCMc1E/xUuvbgQYDjUzL0SNsiDCYD1
t2s0g+IaLuLYNVdE8gxBEPIE4umL4jC4tEFLD8AAnQRHZMmLU9lZ1cK42ANrAtvG
1BmfiF9DvzvGMIwLRZPkTVOuXhFIfSpDBTWaXE9rq2Z4V6uFWRvMYVnlcIstqNNO
1SG0Qm5PhE7UtSscYV2tn/UXOmTkYq3dA9BkeFGXE7ZSGfgnqmZwHwJ8fz2/4taq
Nc7/Bzq8DXIi6EftPIh5n/+T3jnLMlkv5FHbOFon7cwWBRkFcmCw0Qzd6+4QCYcZ
HVOdWpUjvoSJMMeZ01Zz0kVivvBI7YJuMHaIgYp4ZCfqSm51R5VaqDtF8TKcwCvz
Yti3rxz7M5idQZGCro5l2VrZdPQ3eRiDX6XcDAWCbXekmrKGCH+HjS6HYv7q1RlT
XzVpa1w3VfrfJoF3RjHd37uU4DH0pKJVylqh8SOyqPHaSudEMHqu+WUsNSveTSNf
6dp+UErb6luou1rikYb0Bk39MnXNKZVDVhFre8KIu//rdDY9dNpbKZHDAS8n6AnI
0E1jYwQhJUslJeblDQyrQ5ij71gc/lFmEzWLlCm/3J4+jUC26yxIVIxDP+84tuch
gLtozQpCOxcMHJ9xjyYKUyJmuJfuXI4nNwN/18F1MOFWlTksPJ40RcD7GeJYZU3T
cjQS7IdN8NOlyiPz+fFlm5bEwBmYR0K4rQeSQ37toXTid9azslEpIGN62zoTC5X/
jZVbVu9pTjaMZ7FAsJm8BbSr6Sy6oa9Df07iz6VzfomVUWoSTvxpdhQChBV3yaBT
NbXrbodMEVSgzvpml5HYW+CA+UVTWUbz+y3ESeQGPQist3dqgK1z21+siG/Krlo1
fKzIdqLeqiMjsfnq4sXBw4yqCTmHAg0RyhM3iBzPc3x2HYdz1UL7faZml3Ojal5I
NybuNtkGdKUwGRKU+rHsEG6Nhm2CmuQqXOAgD56b+IR4u9220Px/4o2OJ7WdNiw9
E1lKlZCxlyus+3Ui7X1XexAnwZTfPqpytPAgNVibnd8Voc2wAegf8/i0WHFdL39B
T2sBU9HweoQXhPqo3bls3kK3KWxAU9hWdZKV1hUhBuiRQECh5aScJmh2g4izaHw6
X0Yq83fzduxApE8xQTOZhR919EkkUkh+HvjNvq0nGU8jBQp3SWdG6zy42Ip6D4QV
y+MlXBASQP45YrYDbauwRBM9fjkL3NbS/ByRyMhcKaClUw5aUAXC5etH7ud5iyig
0jGqEPyoNfmhJWj1u3yhC31IE5YwS+oXLMKn6Lj7TC8CMiMT/0wrJGCON7p0YLer
pCvrPIJjKUxXhUFftXqXSCSWFix8xDwsLF4zcEQm8liS6cTjLut11izjFE1XmLZ6
e21PjGh6PFNUd0Q4Npg7ZIuj1Pzcxc8Cy/WMR8FdIiH4CGz548Pny0HVWbYtjUsT
6Zk5BNyK59JMosH+Vn+sOeRmexaf2JTtlgNVlpdHj+rZmMzGIX59ryf9vEDuQDlw
iA5i/gjlRz0aZNarP2wnYUHpBCJdIf1rvdiO1htdt9nmYVUHHNzVGESRe7hXp9cF
LRtBhAelVCzbm7r2ehy5g9MG/q/bQ8rturIRWNx7+4fRBsG5hDfQIaHMqZVaVU5g
MUMQVb3Q703r1RRYbHNb4lXc+B5zmpbTF2AhR1yTstRw6vWF9VLQDvcKlKUcaNoU
YfI+KKXEd/AbGiJpM1ugAs8VJE83KBECpp2xJoZHYAb/0astDvGPXGDIqHQ1HVYH
DY8GLoibsYjLOm0Hk66nLN4NC75s5fk0iVhXjcoC3Qbn005ld6mFUMaK3pt60oIC
wxiwQrOt/z4U84mAZIE5pGB70xkVvIJ/5jy/HxR/v5E4OXzPoMgNRUvDmZ+89+rd
viDgJ8CqsvhinAstLaseceZZuqGOTwllbzzHrXB0jyKSs9ugUc5aatQY2MCMwsc1
CAJ/UtR6cxM/IE4WSfMi9cAvD+lbyJqa/mAUQTnxoNK+VzUB4CbCSrGqXVogsxU5
i+jaT+NEhOAmX+pQIdHkLgLqKgcuyXD4sixuGigSCEwYJIPbrXNi3aiSnyBGUh9r
EVz7G173s0+SKCmEQgsN1CcWDxcwZlAVWdD1yfp2Rx54AIx2KPMQbrkQPfP+Jlr/
+HX23TCyRH9sLGddW3AO4+rsfyNnBnS553WVFd7j82tAIRW/7oJOoGL2GLG9q5IL
ZQBSzJGSdVrDPtIcF2W8i9RAmcudTP8ROChRi4w5E4uCQYJVRNMOf5mx9k9KIraI
FZL8odSCt2g8KNkC4IXtUkMXYr4wj9KUHIAYuxsjcv+lQ3BdzXg29Z/6mpaMZXzf
/weTvSm0uP537RoqvOxvA0+Dd7Y4HzmA3btlDZIaAZQ=
`pragma protect end_protected
