// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gjfuJzT7Ys/IiRXAZoB+yFmnU4y3HlJSEKzXYbgDkyXy05bz2H72w1pshCWXYvi4
qa+o/+odUENj9mOw7d6K8vyrx5z+WcCySFdiT8BZO9KBq9Gej0k21L2U9Xei6FNI
71KRu4QfZaqKN+SufGoj+fBjEUdMUkM0as8fsO3OuKY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12000)
TWYNFP9GYvuSGv4ExJZ2IOQLORlChPTEVrwZHiEaKzFriTQrI57jTYp33BYk8IRc
OjOy6+5WxPW/TyacG8XKsOJ3s4JCCNFNMzxErJWJHwD6p4VM70abSk956qDdeCNS
VKgacu3c6GafQ4E2u4f9rJVS1HJAMNFZyhd3hhgpGaZdyAQAK0Al7zyXtDo7Nnlg
sw0JQYEXCeTEXjfZMaRmuJ6Uaio0NbLCx6sI8MqHlbmvyvx+m9+1DcCgRcuH1dQp
9qtw6HzGUrSV/55ZayHiQoFwPyK2aGbO9/nkf72Eirn6nIG+DkBpQyRlHko6xhBL
iCr/7dA5dPxkfY/oT85ewY8a3g0oz3TPTBw0gIcUouS3xchuiwe70swfefhdP5rU
XOAoYtTOD2DFwD6tUPvVaY0LgZVWMcDtVvbsF4mNFObhO2Maq6M/RZX6CDuK3MYI
ItxU+Nx4mhfZScF6c6JWLy+pUdEsd3ZVodv/nvLOGEaqUj3pEAk97FH0k5Tf14cs
ZKhuSoD8GdK5SLLegoFUTPjgHw7bN3THu4fe2I7xz7loz8je1b2595m5IogRj6XJ
9Ds3xUUCpbR24wGy6t9UKe22XxY+ZHhzLGks7BioPazwy58WrGfaGZ0fHS5wtnmR
Enh1HbW0zrki4SPRKcYOxMtLDLpgdUxVWXRePD6AEpB1Jwzm3L+NknDVxq6l9zv+
+vHpZ7cRVzON8jxpw4Klcm1XsmVe0/NzIlldkX2W3Q8HjPIAKwZ9vRA1yoFAOwke
IaFgdI/uogWLZ+5RaUManrvB0a3yH9uXqJ/TBZTxe9xsQjUXeWFL+oYegOiBOb0G
K9M90bwPCb5VXSmeZQo8uZ8t62ZONp4IoDS1q4JabrNLj7gDdINCYSO4LuxnA5/T
RMR4H9qjH5kg6YBYkgzdc8X8qb5fohR9pizsxYpyIXMGWfEkRmyiXNsHdcGIfy9C
H117bQpIY6IKDWzXH9fD6QfUmJClP2vW6dJv/XRM4daA99meqhYFLopv7tRFhZyd
o0rseVIeRt+wy6/YZ0muiqP2OC1+cWI2FR/0ZBjHAHwCfiFDIGJMiHBZrY8dCWBr
575LflOe+raENWCwPKexDwdgxH/XGYlpHds323hCcoJ48TLA/of3cEeN2MWn20Pv
SwaLpYZuJbfEOlr0C8ut0Sh2A58cNiwNc7Ir02sBXtJLSrneyXx/BrA0zsqTTMbk
uS5POfi41TFzaCReri8vY7rtRAcNELORd7MJ+WOdSfhpA8DqjF/jLKngNM+vTMCn
AVletAbcD5pGno9bOHjDb3nfxjZwTeuRR/puin71hThqhp0Mtbxz4gSEIhwDXV4V
lfoty9iCjjKlDLR5PQI0uPOms+ceYL3VNZawel+73yCZ7seuAVmr/Iv4HC3SQ7zQ
RLTQS2yHHEd/cHa4hkonCG7fhOvdnh9+TI+N2JZSJeVroVqBdkTETo8NPgE97kwu
RXNBgaqLhRDYkac5BZ5mwQXgVudQAtl+yRM45KkBASeJGAgEvSPxKmjYBQS7I9OK
dlxraoT6q1L8yHBtfGMGkRP/ONBox7LBydmVNf3lG85stayoOiNqw/uazoa4fLnN
V/hJJyjjUTmaWpa9nzNgZpNGqL5BVDd1HBnyQ2NIMCfX6A7+MW+rssB+BYfhuoQJ
fdBpMTAf+o2zU99LEw1bR5kYMPnAJnfeCaey8sWKCuTl5vcYn6IgcVPfdS1J9H/V
fiWhsW+frQPNt4BKUcs9kM8dy53KD5bqEXevn7GQNQQhXrbBrbkCBJrHwIotavkm
+eQl2KZw3jpkvAl+EhqAgvyVS0NYUScQCqGyzCLBLdUu3nqciDbABI2Jve7FGkDP
9xTr4Nq2gJNKGUWw/Mnhyp5xOryHT/MR9b52sKWEgDT8DJ8oqvDfqEE0KWh4cSi9
XoclMu+BPzQBkSlpSRgKq3P8ffHKQz99CntktGzhe3aB4A20F3NC0hGxhV2ZcRm/
a9MG0RRnDePcvq/SzvY3IdpQ2XbNgk5AAXk5Cnts0EP4y0wBWArGqDjohS4lgtFo
D7eHpf6Ja9Bl3qlBJxTzZoXP1Dm5NAXxWoMcP5k1odakwCg9+yh59Ux/AVtk3Ey5
Ci22JUtceZMPePTeCxCV4CRLxI8WRnr56PnckiX4jpE6OCg+qVkibW8/ScUQKWFm
7dX3yXh6dJG12XMKeqc4UNGXzts+Ai4tZvzTMxGEFIUosHwoW/rdcrd9WPBtlgYK
qNZi8XfYg9zShScqROvZH5j0D3JEHOklgi40XPt0eyylhlS8+57YmnyuVBYBAtJH
xbiGi6Z72//Z+6ww/z3uLtYm4PrPL/6+NWUNudjcqu2R7IptKM+jpVudaMWrIbqe
n6X0jAKFbRNw9+uB16LnoEDjE26zlWLcSuevm7D6uadrqJtRxPyJ1PskN+HKenUJ
aucLGCaqfzX44CY5lpdnA0aIUsaAZHEVIt0/ssFBQI3Psi+lBVeYniNBEal00YQC
zfknfkUafsD5zF3OPVqBf9uhZ92n8VrtE95qQQipHynrgMKEwlf0fEN2V90fGATv
o8u4zubhOJfiYmkqMf1l13WgEfkgEZJPH/xek68fVBogWfiib06H9IPQIVITLsqh
Ew+UdNWpTRmI1VkjCb9HUhHGKCqBJtNml66JZEBMFIoO6dMra1FmEpmOXGKsSmGh
JtuDMZ588zTpUxk0OYWC0JbySsHWaEPEOG+I0adGENjempYiPGJFeARN9F4TlR9y
FnmNgScxRlx0j8IU8rQmJHhkKfHnN9VhmpMoodXZQ3fy0IjizTnb1EtRqPelpDNK
9vQfc1m2+0DtCnIwwS1TbBo6eTidF2TQQ7hbv+ftFxASJXexLlm/7ZmhB9qXfYOm
vzVnLgxt+D2pAsn4tF/7a2aZgEZXnoOElcPlVqMP3y+TLJcUDUJ4eHxGnHyXgnoc
OSweNIeqDvB7My71ibPATv8u+owMa/sLs1qpIiQIfR2hqXJSn3vfD0Zk2/0+yW0y
ni9Hy66miQX18sMMuTKS+1wpk+K2uo7fZ/W9QqqF4+Wz9jNZ704JrboqM/mj57uu
odLPPm8jmd5k0HDRuLUxRgzAzaD226Z+0qyrNnX1KaOqVXVmzkc4cCOLWQu4xKX3
SbCvQ+sXfZQFMBo88L5bu3SWnzR4jfrk5OYm15b938hj9mflytyJsOFWXNLf3SyU
ynvaC9YfTuk/yxBSbr2Yyv/IG7ra91/4lKA7zMgPbOpg1vYR6DEjMgfKnkdX32zZ
0l1nXf153ZHAePdl1iKwtSfvA6qnTp3uy6ERLEZdvSI/7m8vblHv14pjWREgHywT
TjxqyHM7pSMknDqBwxjE8FaniepumJrQOsNFAHC/GXFzh+g3Ny/hEXHRMe3kaH4F
yO0m7Q6Qz+mEe1cigqy0iSmVL37m8c7LmAvL6tkHbN3NHAU2FtM06jNd0NS+lPdy
Yr1IBAl+b95Mi2WY4LjffSk07DP0Y20dUz+SCaXsXBXF0iJ71nhehIwIYU490HPM
vAuAOcGYMaf6lemigknh3AdX1TvOOj0voXfWnsEE+DsLin2HAqFIFPte/04ZJJhj
zMWTWJEser887EYZ4ODBUNTv3sjroB8L+qUPYKSHRHujh2mEEY8bI11iju/6PblC
+nFUpgY4YjYF4wkJqHKwsdTfwMwAIEXzbddwAYEco+/2gVQ8JUS2TxTJ/RXXNNO+
x2BZvLWqV6NaCLYK07ebUDWfnjvRPbLSSLwo5fJW5y7bpSaripzfGzudvwWVd2H1
Arl5B5R97HA4NiR2a2Xk2ojYtebf/Ve89umxW1rZnJ2q7aUWLVX6v8RvkzSIYTJG
tXwK76TPoaxk1JuN9+3w8y9/HEnQRiaKjCRs4L53O/vsJClVEbVkt3A4wQrIas/v
/8d4VWVEcORQwxof9hA1CFgPR3FOgaZa2aAAWc7ccYiRgrzOd775lrThk2NiJVMc
B5Kn+mBdQ7I3YfPxEmS495LR7Ua+jWIYYMsejjIMiIVhpHc9uWindtdF9Ru2sQub
OF8M+SQyEJAw2AuH8uK48nlSKQGuGOFusBupiaSaXVBa3EnsaFERvTEKzJMcP+3Y
Qq/KMgmDjRg5YZTTfQYCXAlycH3K5XTmKlbjMZLjaqOJml4SsIXidN35sKF7GaQz
RSBrHPuAV5TrvO+aX5WSsXqIBlic1RmvuYZMMqz0vjRNuLJC13WNujj7R3tRN6hW
zd4VmIa352yrFtYWllvT0/Oqge306HL8QIlNMCojYdjlMv7ALfQ2aV16ztIVykWU
veVC7s09DiarX/OJ6bmpgOEalag6B3cBTVkLHtAp6+QkpoxtDbPhHanuuh2hjfTt
1sLaMxIoeQrCUBqRgxjvVxs/fEL8ZC1cqZ4HTHZIrCF0VbEs+YsmWNw1m4v69O3W
ijkLUsyUxoHIpP9+LKHtkx7ML3zwQFcE8WC7zGCWyhmY9vMyU3dxkYSqFNwxuSP/
kxOo0wC64KYDvfPYhqPl1E6+3N5DoJcfFVEZWpjY8kiVqhQkpYkHD7EokDs5ODbZ
TOYpmmtLj/PqkiE23lHKC2k+IsvZMMSmhhT2L+0f2NgcOdPMZ+vqiqIXrxXFhLQQ
xdt6i+Rxq6tCDsAyjt53N6PR5S63rQSUCImLXa0jBerx6Q2i40ehOCSutB6iN4Ay
1swIb5Tvm24PRTNEb7Nf0UmlhZlAbTWlJmQG/OBRBgZxkz5VRxya7IPEOOT1WZrF
gIPVBCw6G0VXApm7oYZXPNLVSyBpKqTUQSXVdEJQ9Y+zgHJTrDCAo05Hh5ePHxhq
K3rXz3blcDbllLbWV7JnQCuR0vFoNTGLdh9VAGro3n4BvMbORtLBlMOIN+KWGVkp
rbX7O69nf2P6q+vGr05BUKjgcebEIecUaiHLxsy2lA5KsvI9im+dGjnXPIu4k49v
YhnEHcVmnw+HUcQUlFIExQXiy9CBMCDAS8ghp6T4aKJJMiX/lMYSxCDQvu7m8In9
OaH+fsVD8CmGlGNTYQy10oKNLx0pWtar3kOomoMEi0R/SXjqqpyfRlR2+khInjbK
K+WdGUIzwCcpIvh22yUPQQrymj02jayhVoH+iXv/cWalWtllfcPb6M3BPSbeutsQ
YJw6TjD6fcPrJ4teBfuQMaPHOVc0N39nkLNsQLmawOMyFSjtx8IMFdSZ7Xm7Fcu5
GqVZoMmfVgfYC9avx+lY2IERAfGgUFW71WknWCnFWrbUukJvCh19Adg+LnRtye/m
LM0rkfblEUoJZ8/UUlWXa5z2JNXDDpWM3XFBhwXWAknszxcXptIzkZyOrZLvli+H
o4w+9gVCK5dBfsv20b5xc1ndQxqpZSohbL6QCNINiZAZ8QsqzwfcI3nmFUlSI5ye
OwFNND/+6QpT3v8K4BGkr3AyOXzJX12PdotAARsE96X9rtY+fQZpFqVE3+O7WRBH
mW67139ErruUksfjFcwXD9bOD1PUGXI6Hzxle9WdMZM0MyPEiZMCaucrDTouDmTH
NmN8St4kvuZann7KrzKwbUDc2t+4vseEvKSTNlUaWWy2PTzTVhD2IyvjJIbQl7GM
OBKoZ8QgD6W7uKmjncTQlohMbZ5iBBY6fjDg1fKtoqbyjd/tcOdbit1FelLwpc+v
IWRbYRaNKLMD95rKYQtZO0oNnDYWAvabL8hncffWHvPwGzHEF3lo36+0IJkftNup
UNJbtlnzbOsngHQXREzr+WS4sIjGjtB8yTozJ87LsDgAMQVfzRCeNWKQlGM9JBEQ
xt5oqxgQkf+H9ceDIf/lYnVqS//DqtVu9KfDUBZJoTBi8dJrSDiYqubFlhG6Rh1W
YJPxRu4372p35yKbhSY4bpKBIzS0tklD+RWo1AB5tFN5NSoyKRlWL9uwvJix0NL1
Y5zDubDZgh/tmMLq4PlnwSV6oe9wXxlnMC0b4HUH6woB7bEQm60GyKidhrjITF1O
xKJXrByEmclORC00cJxKslnwJeMr9aReES8KXgu2YzoVKpsBb1k0mDg6z+a1PJsN
MuBP2WF1uLLxkPQXYKVH1UjfZujDeMB62BK+vS0WQAei+typam0bW3qklwnsLoc4
/o3X9E1HLF8MA/GODJ+fSs+g9GgNc+ezpJK8Px9Cpdaa1lvFF3GX0uGyrs9Cp2VL
QLlWMqarM/+JwssSIEcaTdUu2XMbfoBDd4qcAu950IgMa3WjqZWNBFmqSsaLsT8t
AdCLQxKLsjgqG34fvoQY47GNvl/EQ2OhEPfdsqvK/sA8nYj3JKT6tZmkZRbMyzNs
HM3WajiG8/RNC5CdK5/ONxIYpOZaVZWvSmydtskeTR2U+PIw7Y5YlSIFs5x46iga
OOKKlCrcyMTRaHfwd6uGcbyFPbBv8gGxqKuabyy6cczP8WZIG3Zn0HEdI2YSiBe3
FJrUQ68eKMZH5FJBKvNhqlejii7tWWrUUP1m0CUZifTtxePmjZHPCX8b66lRemdx
WY6LorZiosex7dX4s58se1ihsqpbLUOWzhIWUgEKR4I5lfEJou5dJQSRX32wGjc4
LnaUlkm2iZaMXhHPG9+/CxOC4KXbVlqCQqaYlczb/lGXJSc+kS3zajNrTmnDGVUu
da48PotXfDjZvZdM8giZEzHNoQJ5BeVnQcaMJS/3X+J3Yjz5MYpp8M0tjk90HiJ7
1b1x9jKunKf+/T9zAV6rtwcanijZ4KrGKFXPEshDaa3YIidjM4UbML41XSAXymvs
LWm67nzx6VeDO0rr2aoDiYPqYA5yup801K4LnDNR8CKWB6rMlbeReEbLgJOvWnl0
xkXBZBchNS7nTeb1VnyZ4ibvrKfTAP4KsQCHnK2oHPBoBhQUcI5OpzymQ0L1zwYC
mFfMffTUSwEGRxwaPUHnICSHTNo4RJmxf+6KdRoWwuYFrMN2sN4EwlMABz8FK9eF
TDDw7KL//1j1rBia6xqq6ic4AFn1oP2Sq+AIit9CknPp0Jrex+3KtxbWQMI0FubY
fzhaAh6atFItaBycelM/pcVvLBUJCf3myp9x6l1H/Rv67LD8gLarlFtTTzP6oP8e
jS6mjRoc9VZB1afSal8P++iVBqNn9FoY1BvkqZaxOWa4meCUf90gSNKXIW59SCJ3
c0sTNWeYg85B8FODlFlUTpXYp0z4tJ2PFKJglx+OgGCOBHvTcd6GoRPt+H1pRZZi
4otA4fd1eNpO4BiXAGx1mYwLd2EaS5YXdxF+ZYh0eibRg8X8OPONDbVWjtLkc9bu
tDqZuWFOWGFEiEMp4XGGVxpkPIwjM+ztpSky43iwT2HCXlFcJrfTKRyV/Zmm4yMB
Kz4/zzvvfquwNrgn5CrRu7zJaB1INdsfYeaZ/25mAjPdFQYF2RqFJWj7IOX6BP9o
iqZ1z6+jclVn/yQqHVdkxBgIsITbmtlqYQ2uWBXhprQavIhXWrrLl3emu2xQAPas
R0z9wj4gXF7vKzqCSbJw7h4Yf8wuZ/o6Fq4YaSHmLTLjHseYezDgS9pno5pN+Htq
5NhV+FyktGkq63hwfJid4uq3lsHhhvTVcv2UVpC8hds5/3Ld3J2u2tOhJCtTvyRh
Zu6p81aclMdkxIsAtfMQbbpc80Hq74tHskC5hh3dKE0hpPbTWU9j9vYDzhg5Q3B5
ipQHNeabwp7NS1k7BpU/4qqn3WbvuqsEyTe8tL/ZvBD9KO0Gx47ZRSfEe7fPpKdc
gPnbWq+UcWJjqGG5IplAiHdXHWLffOn+3o78NXzxNpN20weJPvfL9ThV7DBQSz3J
K5BQPA3Xi4TQRaRhdujX/9xbVLnk6SKLVLALSGsVnwQPZNPmK4y1v60W+D42TmcM
F5QaKUdrBYv4eak6yqQwffRBGv1YToXBd177CWnruscWavtH2bJW7VpjQv6ZKroc
igPXc4rlEOh+Z3WBsTOBC5myGYKS7YUimNjHrl0K70Y9NDf7/rG7lf5ZbTEj48FH
p7SuBo1p/6REnr7hrC/DJT+U/4Wr4qkMuhHQeCs0/fmgtKgHdsxeCStliSbOvzvu
RSukdpZPECP5N4asLI0yA+Mp1cnMoeyf3ZH5Mn6Ri+9YtKHolbTom6/+hp2wOdy9
ffHEBU8kFnP2Gf4EFlq07EDzTte2hplTxRh5gwgt6TRNpFxHVVHHM7rFLAMbrMZZ
ivVmW7PxdSz7cMAKV4HdkXVVmTOoDt67XGjEDIceOu2gxoSoyCF/lPlTu4xKB58o
Dw/9VhuxUUE79btbdnc0Aw4LZEYnsO1XT02C9wGAscTZtOUVH2SGXbvKSzTxPDQG
/y3cz0xnp+0sI0W3dxVeG9/vfYsm+jU2kD38AvKAmeH94IEfPYWBkp1x8Ejcnpgs
bvf377MKNL44yuA/5SGbR07QVafzHwo9AnCFaCOCH1AbGMzshMfbuJFj65jjoQmv
ABnJQZWu+Q5z41Eh3ONoOl1+ZCdKbQvJN3Z30vwsl/NedJyTjLktdv7W6PC1wWl+
9OA7+QNkBOxJ/fJgpA2/4WQEFl4GQbpo3AcEdsfPjBokJ1235Hyr2jSUyj1mE9Yy
uss1H2n2waSKV83GcBxDsKPLpiHwpgf7GMwthHDGwl/uhxlcfnPTgm6/VM+Cfhsb
Eyjt9EBS39du6o5um72b861sm6AJz0qIbgQmqGFxmQVK7+sZxAcjeOWpyxySgnKr
KuxixOVxLAh76PTHKPyYGDA3NW76F4OY9bClWom/yhYXqtm1oTZ5hfO/gwkeDI7L
qRXTHOw0ue5FTDaKCBTStJCngFUwhfVyufeGTrWxbdWbdKckic/k5BfmyPuHZuBP
PCvFRui6yJxAUhpwyUl7WhjzIIDwiTjz2Hc7HgPvAu25eIrSwj7yNJtn0MWnpxry
HYJMCYKGcTm9b2i2DhFAN28o7b2qRLrFfcSEeclbSS2GsFhr9InEDgsnGTdYDrjV
bAGYomw0qF08u/iWD8KowU23re0LnEUKHziPxTlNfgJXkXIgKwO9XT0EhdGZL5Gg
XSJIxhOqJez/umqpmBMcV8txHrfESLsUBMPTz+QGpnm5nJUan2jv0ieUvPAmV3uv
2xcZpI5b2zIwFU82GJDNep6UhgOqwmzhYrewFQdbu+gMMbqe3RZGXOqw3Cp+tv3N
ILA7I+Y91olh5Y2BUOysHb11PRSXAQV+oendujZR4vIWOPSOPDPsbIc738Ck4ffq
QcsIlTsajDOUMxsGiZP6CUPtomgEAD8WxeuxMpgR6awg3d2bjqBmP0Ce6V/WKamY
dsyLmkTK2g474JscZhVvUWbcpl5kvWKSM6SujWD2gsmRTQ98eCG502sabUQ0FkxD
PTCQrJ6lLH50GyOufpjQGEfLWFySJmkvR29tPkR86B68uWvbHJNcfPCsxXJ3h3Jc
IfAzVpEaJlY+od9MS2dVxFkVyg4kjUdfMcOxFBD8uqYXdaDe59wWwWO3HnMVeKcK
OqJDOPcBNQN8XYgMMC7yIqGanUFy1uHZu/1NwQjcy2wOCD9ienYKFA9zeCKKXeWZ
zJc0zlSVAwPHP7jKnVparkgjuh2FcXO5vrXpXXmc47DxYnYq7TpU0eXel0nzpdD3
uyXr4Vdb+w/Tje8AyQs4gSZvBqB1KyF82TE/UameYUzun3uOvM3ZwQvH4IGpUHNe
yykkBawt4itq+2ZzpudEwMtUcvB6djfMFw7h/Qp8XwoAT4yb55sYcSMwLiN+k0MN
rp9jos7pjsfIuVG8ziLZyca8fZMWXOpretg2O3XAcKgBOtfKKJ01hesbe0tIucxX
ZunMVot56WmYMXTJhXN7Kz98LCDUnzMkltbNgDM6U0EaOcmmJKFOkM4HbtFa/YW/
/kApSyoFt9tnBudzxotLmp1cMU3A6UiCX7pyqXu6Izdb7hy7sDCTp4owbiRDvTL6
MqY107GG/0a8xaa+teCP+P5r2XZI33jPCt6PSYZQ5rhrvgCbQInWo3aQDHtpKUD9
7FEqTyg4ryWndvptHtwi1BstA3qpof7DrmOEKBerlRDrAniomC2g2Ashznk6mmUT
dC423FEGLl++7zAUQMmDlufdlYM/DxC8XkisavlzYrnQznFZJaK7ir0W2zucsUKn
zH0NRcJLThugPk40NBKt7LY6xhEheoZFHQoQLk4Bdj5A0JthngnHP3zpCaF+BeBC
g9j2GD4sPW1VGRZylOUKaGsn32TFTrI6Iau/VVgbnnOkrAtsx0skivEZtkn4RxWj
FHNfLMjCyptKovT1udwtlkizYTtFzOOOU8FCjLLc+R1J0f4CDYWBmRpLA8AWggs7
9GeM5MvbTwt1KWz8WQKmon3aDEAUca/28wX51y8AUSv6vgrX7XIavgnWHWXtnT2L
V7sn4h3X+pBmsaavihUjTjnRQUEv8i0zSALdBC1nWvtd5CHQOHJnKEkSUpwioqqG
+i9XcBij4UQvr1W1us+7Lfl9r8XhcPjhrU4HZaMtKy20zVKJCnGzhpu++p1nR2jE
5gwz66lDBQJKkHiYA7BJ+RpKiPB28xjATPnUVqvpe53hCxdSLHQy49yoiXpE3ABP
zEUAAVdArTrbkEpLc9we15/wkhBf3fgr5/zoBDsmR0c8xfQHaWGSxca4vR/5CCNm
nQlmoUoLyoMYwHyphVbKYzmyRulfBQ7Fzu4G+eyYpd1s1u0gOXoKF9fihYfJJO4j
M1NnZZQAkYg6oZ0csya++JWg5S8RQoJRCCUzAU6GP222KeD6+ww1/zI2pmzy6P1q
LdcsuMc0WfxegpllF0EpzlL9n+dzC4r02wZ9OAqHjVUqGLJwTCLlYIzLPmzxP7S7
s3kHTvWcJtiTMic1N5oAN0zyV+4XpviIH7JsxsE8NfGuH3J0oo95GUj/7NT/Xmyi
YvaauKrJtXHLM+EzKv5HDvQPMkPZzGTD59gyyFSJYV2BNbrKC2iYUXIv1bI9kNug
lhiEZf5UwGgCIp01tMcL/YY+9amdiveDlVW1vfGt5Kxm+jOVDElaWlsd8PeTq+V4
d1xDzmqI4QLekcygtD5sAXqajpYzHg8adJgt4vRmB5h480Bh4h45wr8sJgr5ld1k
PXK8PiJ9Man/7BYxoSaxMLxcqr5OufDgscUfSzWkx/AofthnozoX5ldo+ou0jFyL
+n/z2ClXxyZl2tnNAr961kc745sMqaqI2on/p+J6ml/Fi8J6AZw+xHwXLlE3kMx/
MTCa5PQ+JCKoN9hXOGD86cVQxUFiqmqAQypJe+BLQuol8ZP9aFyZZj3NeuniV3VA
9T1xpPcAXxBmtNbolAG98ygBy4aHhhY/1rW23kXGyIGP1Kx5LYyUGxp8XD43MnDi
jovJOAQ3Azn8j/2AgspgYfM2dAND29XA4npqfkXyqBIicSfKQdkiqSl97fzy54Pp
JwpXyEiYgu960TzkxfsvO+NhzgySLzSK16mzzYBQ7qwxCWtH3ydF+wxUsJbPtT6H
vSGTj6IAudm54QCL0p0NlhPJ50/46kWohdwnYcaAaktb/tWdYhAqhsAI1MoeaJCQ
VFakIAWNkFvVmp29a3pYR4b6qvm0R5Xzw96svKad1+jIVRt5XR71Blra7ONGpNn6
ZCOdWlHdTvAXZc6aR+x07QyWjTtuqE5TqEMlm5I9VjFW+ew4p7YMye3YSFhb9lyZ
1ZaBRTHSZc+J8twK0tH1CEdWE/6fj1N0VI6spkCXbZQiVuzdAdZPpby5hSvHrrz9
bm9/qz5pn6TtkcbsoCWGq/InvUHJP6LMAzjbZbDLvyCMaEEJjsL3FaFZWGJHj40C
y3truIoaN9U8gkhZZWN+4M9xKNpHJOMiqu/WdGITrWrUx2AaM1IRx+5ZDZEokJ0L
r/7irflurqZP5ENMAc3YSptUQvyRmBEnM5gl0osD5WCBpShIXGxaiATtGzucJh9r
sjhEb9mrvwMjh8uUcqTu0LVOEWEnTquaCo5Qtv0+UOO7HvGUGx03lgRH7tYTZqX8
ECGCceAMc41oE+vDHZ64xy7LnAFoQDEQIsnePETAHXKpbl9NTilBy2VF9u+l/5EM
ZGjhFLixFtbGz8kEWWmX81/BRJ2P+l6lHnGqQzrpHlkqdcR3KtUpOiwhBn9Wly9u
vIawXV6uSwhMQZvrz2139qeI4v58Q3nrafw3JuFaEVE2S1RjQBZosGlXBoQUcCHI
ukortqiURQILZZ0GRjSZoST8v5sIkB3GO3N7ysU6cyovGkxfeQfyFeAlZtXXRkCr
Bv019EgUC4jycmPG9RJZMnA4dEDkH2meYp8xc0zc8dX+LzoHP0QWp0+lDo5TUStW
07T9M+/ezKpsDtHTP+mlh3Df1HrGCDn2EwMGTlIb/sMcIJ3+OdnmcY9BbbkOxG0k
kdK3S5qQcKTvkMScE9OjlEJcFm+1hfEHyqM3j0+zJYLAbEIOl+O3fqDUyF5sqERR
X+9h/VCSNpgoV7y31LURmkZd8WA/H9cxvfgpYrKzt6xGjsuGgurGlxta+bmriT8m
ZZhqMH/u7QEk1m7JlWNXbolzS7yFyZATUH0Cr5vCNz5nTrleG6SjmvYhUYkTwizH
pEedtdceRoP/B1KNhmXYeaf74an/Hj8qQYwU+lVQB81Gcv9jx2Pl7t1ETpjUTkXx
WICpGM6hizankWWH4o8qDyFZev/eCGNp71+shr0WnP5eJnTt0ryir674vSAitYCf
WgsYpmsLw98dWLsxZ5aTl6K9yuH47JDhbt0CP2nDXOnJwWyUbqeiDpyOgusWvEaS
IelHtYmwK49/Y7eAngMeb54MRHMCmKme34OY207kr4RV6PmqK6mSrjIF8/cmM4Zy
ArOG0NMbN1rNAdD+5ry/py7Vkafj1Mu+pPO0fvYoxLMfx6ek4e0Pt77Ek+oEpIey
ZxSi3kituv+qwHHvWe+HC5iu9gz6yTlpl9s2FD2/NeSOXT05Xqd/qNznyZ3MEMtn
HBy9dSCHFhd6CXkjk86WCwuAluG0+OKFxA6fgeeLgmjxHNBonTrnxhLtEPHo2166
TveB3Fm6rSyRfnspBZicLJBDg4bZcNJb3SIr6HQLEFRMaj7rCEB1YH9KnnkkYXRx
eIEKaYFMkLxc9txdXlZDnbav+yk5fBxcVlOrwX4GbnoMOXpsw8uMsEqD9ll5Ccw+
jrYMPDK6V2+afFNK8/++L71kdhVttqaBO/vXdzoAOO6J9PI6X0SaUQo7QzyZcIRT
rVGfHeogl0enjLUjqVZcdrZ2HC1Ss5+Uec9H07OCHjqT6F3UmLKIsilLHQyNWJth
Q72mqjgwyRsFQ6Iz/DuZkZYZGckEDBqalLxWWqdwKV2FhoXnR7oiZfQyWCZKhofx
G1D10YWJEySOhk3faQp5AZqtu5GPl9wPkL9Llmm0aDU8sUuENBAkpEr06xqx8/WB
8wVZ6AgnmsMXPvLmmyxIOmXn1woPxdGHxPnFgfIK2NcE+qICnWfzC/SxrPHpltm+
iSxeoq5YHkN2lC0LFTONq1aefIDnfY2XFZcrZuOEhIuOiVdTSXg8HhIifA6eQAV/
Nikxjvcn94EVxj3YnKIqLmNHrl6Dc+8Kx6GUnurfwbdEVWLxGKw4wjKthGsHrx/E
xJGLhg8h2O3kpbmUjoL/r5x8mhzYJHAtMknwhtPt9uKCyrzUewB8OzHy4T1RXe+z
p9higE4RH8x7j1Ou8RVKyhyRMrTr2d4YyGCQxa7iDHBi4F309pPWMHU5vn2LJQSl
DRX5cq+wc8UvYvynfiWVuh8m63k6VXoKskcK9O0NymAch6F8REzjxJZGFA+87WSF
iBp5Njj0zIFmSgqDe/N3vsn4bVpyULNej9y43eylj7LlZhC69DILpwNI80uKc0C2
/Sa1wkSFndbPM8uXaiKsjRbFBfARTWT7zu2FbvRbmNRag6XM7K5mctUnHipeXCfN
Us2CfeMs0wPsxND/uz5J/IST93iIhbzWkp9vLd/3LLv/hCyviBukxcUuCVrQDW2l
6Ep2P31A1nZ4MJSovUZdQUn9j+P3hPOnrI9SNpHiLySSz6fWaAiwyknrPvxJ33Ar
dSPCN8m5ZcMruL/4HpwiYddF0cwrGTfIHIxF8pyDduiVdI5K5waMgWWL/Vp7kKQb
EMAvWO6ULCXxcIaqcZbcXqV3NAPeo4r2VbuLtgp13j9IvtnqL9DUo87SZZI4vW8y
+BdF4elnMefwtPGqbckCTHIWtS90BgzTTSYuhO7AfcakkqcOKhIWwh3ROzwVnmNZ
s7sLGCY05nem1LeaceyGP7ZhQEVx4mzNNY4mbNbMgUUE4N9XOFFjB8A/CwVJmAT6
FIO3q3cLN1+timQ8RBs4RNA78FU67bjVHUKAye4CKROTDKdGUzktU3RVxIPFjAWe
Zge9penlYnCQWhocHeoZmd161xh4H0Lh1nj0eSBL1mdz1PnJ5bQsSg8cOMLHwMVV
rHRpMkEUp9/36cArY7Lm8melyZpdI5aRp8IeUm+NyjSfP8sPfrzKOzvsiLyAHff6
tS2EHAYLwWQSlk9MrrSI/A0WrWQGKMmYEvHjdSeOTVngFTiq+SXtrcv9k+egzOQg
JMnd0TdwiaP/IJNwkpg98+dK9HsfUV7rs10sXo0zR7iSgBn5BMUdwR6avdbrGoNT
kyvEhikUE9mj4NfA+K+qf8ug9Dr/wvCBa+5t/fX+nEUFPVCwyyYshodWIDuSBvu1
VszLgb4jTZGrhYlz9E6FxWwQcuh8kcnfp4sQTN1u8PAXKTLxMtehMXicklVhsBqD
3ql+17EA6sDDJkC0Ll6hsJAibCn59tGNMMUVzX/Gl83PZgRJZwDP0icjXkxdIQiH
32jMOi6ObKu7QLX1S+tfG5ebcsshiBQRvagFUrSJaejhqABmGi3f2rmkexqOQl3a
WW5jBhwUtl7kWwd/LR6m4s0bugpUm7KqKWNb6MfjPu7RToRkuhf7YuND2/1ufDtP
O6lmHL0Qn1FpFPYAqIfcGB6A6E0A2Ez5nnj8tAT74rIgE0/1C9w+BeS3vx+UwONB
FtviEH7FmMriy0sfkNYI3OFPyXckLE4qv83LEKNWv8S/UITPdy7giUYEFbwY0OuC
eLZmI84zDYh+mHpxqeetOqJqSUsLAIyK7Kqoek1USN4IsFOfFd8uW1Fh6hgLoAw+
tfKwmqlE2SokhP0xh6zXA4IeI5xQlzUId3K2qZJPw2s/docAjr9J7nd3wboRbZsb
OvMI5AscKDnQVLXlTW8Eb6hqlUpE7AZJL/GZJufz6fKHHE9LRlJgyYERsUuP1MeC
lE3r9Mi9dGy5cSgPUdtm2CZUd8XLpHDdSV2vfeFbCuSe/8k6Bw3P1wF0dkef3cUD
uc8edD0p94WIm6hqtml78dg3Zv/EQPXitKfPpUvGelStFUc5/A7L08h80Cv6duDq
exwB/yOkT9YPMgHYwSNUHQ6p21FEfw1JRP+zrZYgHT2LyJhicGsBjn2i91bI+7lS
UNe4IzGOGq/S99x8bpOe4Jkw1YrvXGEUiZaW5mVmhhpIQ7CUSGH4ZZtKBjMc7H4u
V8T8OYqwWnyG51WL/vGpgVcVFtO3BKusJvPECVYZazrmtASRfERKGfL3qm2pM1PD
jsuXkTH7LF/8rrQEfDEtZIS5ZRdO7WCLbTf4qcCeqodvTkvNh89NSgy0y19/V+H0
Fw1TexJAVihz1FfYZd+vTRNB26BmDPoiz4iH0lFV3aBrMfZP/3E/LiBAynGMGvM+
3tmnI9t0TKpgpcKVjT+Qf7WGUcjmKkcEyELj7+xzpdk7nvoOBgoDv8sX72EYzZGB
ep4nLNarXvD716FFr+CP4kzAgfCpZntU3qPSTku1pHWhI85E/TTKj7u8TtJrRGGO
4/gB4ia1J8dBMGfBqEY1VroRX+PlLCj+ruc/zRE1HMIQp39dj8wo8nhj8HhirTQU
DL99P8H46FTO5Esl2X6DDY9WRTmUgpvssaRQ9E+/kiZTlQnjETWejThQQ0mHWwOj
xY7CT2YirPLeP6kzS8Ueuy3zo5hlb+80IZNoqNRnRINFnOBSK3MEZRX6LsS2AxSP
obh9gHd9cZ4gTk6fvcxmI/STOYhw8bRafdiIXPwRcAsGd31SJKXXgdQdWpdMA959
`pragma protect end_protected
