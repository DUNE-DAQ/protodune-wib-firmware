// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H^%=@R(JG72^5#OYAGY B^7?Z*94E\T6/TVN/=0WMP<PH/I,0"F4BC   
HDH4%H+KZNK/_0H>CW\^+S.%S,$NO P/$)?R5/^2JIRR\H_1 Z^#:5@  
HW[4?;/G74W6YC F%&2C91&O;@I6;*!4F*'3K0S>7J^ IUD$JT3BA"@  
H@%'Q%$B-;*=H=R_V)\L#QPY=IE%C@)"0NZ=[_C&8L'$U;-E-%N\S:   
HLM97O>Z?C*]@G<M%%=ENM?5RIGF7T+W=S&#N*P9O81JCIK(V6/G\-P  
`pragma protect encoding=(enctype="uuencode",bytes=5264        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@M.=WR6")]C7>PVHV?K.39"A6+\HV@^3F]R"L$B*==)0 
@U%PXF9T?!TZ=!JO67ZM8-A5#9=U-"1^PC]D@@Q76M;D 
@93I2X!)3'!*4UY0L[J>8:=J\Z5>L!$T"6]GY_NL__'P 
@05;IMY7'-4GAL5]E9 >@.FWYN00, !6I1?6R#<@1&;H 
@Q7UIC&8QJC[LRFL)J9#^&&8\ 9T9K&\.HK!"8O%GQ;$ 
@DZ-XCSO_J[!PL:JLG.8W5Y).%AL !^XN9$:&GMAD#F< 
@A9\))0WK,]XP$Q?RG0S]"!(PGP.PKH<0AZ0/6W[;2NX 
@@G*>R3661^DN'.D3$) _:QQG5Y5123\^7)RW>L5X>*X 
@F GB3ZVF#NE.ZU*_.2F@"U)@[D[.QQFVPLM?\?(,;^8 
@+V!8D$ JJV"&+(NI.+8ZPJ3GA-O&L7B_^Y"#3EQK8$\ 
@P\E',CC(+94>"@\.I$&7!=;&E3N0]"J\IFZG,#A0BA  
@PZ"Z;ON]"21 Q^'JPC>OX@;&I/6$K_GR]\I3'#HSKD@ 
@A29/3VM$LRNFB)N*[;B9L/X!4V<(ZK.I\AG8% =[?$L 
@7=02^-HOQ&*1$>\=T$7:.OC73A%Z"P_CZ4(\*7P=:D4 
@FSCM"C<4_*3(I"@R8TY$(Q)J&7XT09.GI(83<*&34&( 
@11/XF)1.N 63OE0FGV-O31;GRXS5!%1M.#%#8XKUU[8 
@M@@FB-D<KLWR+EBJ&:I2M0-X)JK67-9KKH72;YD1:R  
@^/0'C1R1",Y[*!8@,E@]%K_49^N_(":!//KF>+G<[/  
@*_@7U A*GSYYP\A1GV>E*;SDGD]B]P'O8KAX9>2:_*@ 
@SMKA\0 *E_%;,P:+-$O :_!7H6%)$7*!?N+J9'BAP'@ 
@#47])-O'ZY3IT![RYCHL3B7!$/:^9G1JX5A.3"H1V/< 
@X9^>S0?7(6S=A9+G;/IUI@TYA>F=![U5G,#Z"A'[$6  
@Y%TO >V36@"=[\MS=F<?<9.\A9+JI Z_[TK3LY_-"&0 
@X\'H"@"=@D^#A1];=2X0&AP.J;F66GB]:2&)?%H^4 X 
@8:J^71)42@8'EWU%^,U'8LY:05W=)\_$B*#YXG]:RH4 
@LW(<[R3V/74_LP:]ZT:YT!9<P3&C$4C/S!51W(V$<SH 
@3AI%RQS@/PAH89=H7QIQ'J,C"MC:A]ZY9=$^LH!=MO@ 
@ *Y'43#F :"2-X\2"8<](2V-SZA-<4"BX20!:/:([1, 
@:#"6PO&'D3!BK=$1)V:&36-+TL?]O_>Q@&G\1#F ^A\ 
@_-(>O7Z>D*_:J%8]6,P(X _2H%D#3UZK$EC 4[K<+EX 
@9C)(^YP>X3Q)\Q.."60Q1E3"CGO@C[2HUZ>Y[M21Y4T 
@4U$GLN<#$$77U"?=1DXBB<&9Q+U1(^$H@Q 77<_"U>8 
@XN"YZ,GE!O#/]>M+&..DCCJ,<0=]ZQ@C)T)_<Y_-[C, 
@O<*R.+R\P7!/#?PN<U>67;P4&P6JJKP#EDK$ QY3K]T 
@U!QAO"HR??X.=X='M FVVY0:Q?=K:&7)0I^PVY3(9\X 
@_LIL,+,R6_0WG'4A0C$<@W*<KB[[/BLZ$ALL%[^1P,L 
@V!JM[E$\ Y4*#]B!!H G?KU'-\XB]-+0I6/TE[&R$=4 
@NU6OGA9+3M:2A^"$@\!5ZEF;1K51+H,MK=@1Z(@&U>( 
@2W!+V:VA0QHJ/X(CD+#(=. W'&-UNV"B%XS.B",<Z.4 
@,M%N9&)H>]/[K/0D<\YF+971'9;61 85NZHQDRA:DG  
@)F9KFE?AF\ZK2CZ&V],DU+V4<8:.JR9VYV##%H]S/Q4 
@_H(D?V?Z#8RNE0^Q%(E+_##6^ZYV(,&38FD[ N_N=FP 
@P]5%'G"2<%'MZ1N?F@F7:G3M+(HM'*.7+S?Y:CF.XDH 
@Q+^7$PL;(::TK< #W6$F;I8C8 O=:"2/>*9SP37X: $ 
@^(XE&RBH"1J"O*FD1WN<!9C&EFSA[_+"H\&6L<[G !P 
@,HJ'1A5/+88>7'AU96_#S9\N3/3D'.=X>*"(U%V(-K  
@TK9IBGQSQ^5&06*:*:L$N,;6S3-AA.+<L_)OC<@]OO< 
@O%35N[VD[TB>#8FZKZV0XK5:2#_,0 Q#E!EP6.)?'B@ 
@:@)<F.J"XEI7Q-O2*= 70KO9:7?:72;PV2\;K-C/Q!8 
@E"/\H@&U5ZB^&MZZ:4\"KIV5R4EZ;_'8.<;]MY11;2@ 
@7^!YCJX'1_XB0MJ_V1'6==?]86/@RW!9HO-90>,?^_L 
@TPZWGT;W45P<Q=A9%\S3S6G*1)LM3'C9QZ\QDOF1H1\ 
@^Z,U*G:6X3%!21*!>BP/V@#4-@^9OHOY,-;9Z*/NE&T 
@-I))FQ30[O$C%K]U1I%E[D;-=(!(P[%IY;.P-9**?%\ 
@$!@&%3'=7W>4&:/X66M#%;MK'TBH=0<EXZXS#X-QC:D 
@<10&E^:I&>809]"5?=:EMM":+S6>B-L$:!$7'",4"X4 
@#FV[4-P7]-L9\=4L0;:!X.2:]B_S&1H2[]1[_??8V_D 
@-D(Y![IR.WD'EI_MOXKD>26'FQ5"V*A )\C;V4?@,]P 
@RHB^]C(<F,H;D0J9*6J0==<H-.V*'%#W0IU92P\>3'P 
@!NJ @&;FMBN)@JZ=1?D\9LTJBD"_E#PXW[8A8:BH*3, 
@^&46CBGVT\)#Y'QWB%^<H?LKN#WN<6YQUE?NZ.1NG L 
@U??VUI ,9O&O<UKYXW\[8+>LJ4(>R6,":#ME3W+]U^X 
@__/FE<R NV@/!:>\XN+-<_3X:CO0%A3VU7A*YH!(8_$ 
@H_@GU7P)]K7\"7Z=R3YP;X=CX:YGL.\B^6UQWC!EY5T 
@K1'[A]YC3YH[ZE=DSORG:;Q#0_O7XW"B5S*"XV@><MD 
@CS2%U#GL3Y\J_DCF.^4]1Y$9D_YGV!;,'4K,5^Y!H1@ 
@@6,*R)0 6W!O&T]>\VUL?Y\ P ?99]]ZP?2_EXI,850 
@Y*45S4HP:4]MM+S[A!A&M9V5!>WQ/<O[**CRW\C6FLL 
@.Z4*65$FI >%@2(,A<NVD0!G*\0V_+ D0;IB%SOKP;  
@HYIYRW7H7$P#[GKD,T0_^3P*^X6X&$ 0F/T#1AI3WM\ 
@FN_F(7BJDX<X%4NJU1=U5:C-&B)JKA.^XFL@F,*%;T\ 
@R$3-D*O$]O>*K7F*BIH:<-[RF\CDGC7F9>ZK3?Q\XF< 
@] $;@5+Z5!P_TWG,1$5 GH!&P9O*FMWH7X-Y\WPEZL0 
@@4-]JB#]]0<#41 */PPK1@/HOI1<[+IM3RA.*+I_35L 
@VK"A7L9Q<)$1+I0RYZSW#UH5X@-'FK(<!/NR819V= T 
@.ZED  ,--5NC<T\5_\I6V>B=[^$S?:?-G[+!3,OQ$D4 
@U&(<\1O@_*:^;B$]RW$H3DQC]ZJ!QH5_4Y:T#JRWO,0 
@J>;RD*==![-;7>QO%9"3!EH\?^O V7'H!0W%<]E7ELD 
@P_$B\PPBKC,_TS"P_?[5UZ8%2,*.B-V@P\V;_C<W_F\ 
@1?"84SZ&2-?5/B]),@YT6PPU/J3#M3H3*:-UWP8Q3;4 
@JMQF33/O](BN!2&_ <$FE2KW7QKCT;:C:2K15C5WL14 
@[VL(GFH@@LOE*KM57U$4Z83Z_\&1S0S.-F105X=V5!0 
@DR;E=S_DY69FTR3*((EJOR8YZ0([H2G7+(SB]KL5EN4 
@20DK[5D":RANF9PX9&!^%3U; /C=-XHN17+AP.-4Q0  
@<F!NB.TJ]Y69[Q*-"LLW:1;\H+R9(#,#:K\@I$$>=7( 
@?5(>']6W\EWF@(".T=4&3@_4;_BPG#,P";AFJIDG'/4 
@/\A)WB^%%)H04SXM35>$._@["F21_M4Q"XK?Z)="F9  
@!Q;[1SVP('2B#6L_>P!+]G#C01DI5P:Q _]GWZ&;$@  
@ETK;]L/.?*'RZ C14H "LN^/O^\0K04^;5O]3MU;IH\ 
@GT!EZ/9RK^PH@#<S&[8PQN&+F%3M&GLB2TK>0(6 VC@ 
@#A#_X(3,P[+"J,)!W(/JSSN=T;98R#+T9I^'AQ734#0 
@XQ]M_R)G[)CEGT58/!.$DMZ>%PIHR!C 3>QP0A8^E4< 
@*"=*7PO$*KP9]+R<Z>5YE7)GF@H;VS9&@6P[G68?N<H 
@Y[L8J?ME=UV00_<J?DHIX"T.Z$+J/'V2U;.VP"8!X$L 
@-4-6O\H52 _R^OE223^N"7Z0B^>M<\*P/PP97_!E)*@ 
@ZMO=$(O I-<3U'UE#6K#AEL#[=#SZ4T7L$289.*1!J@ 
@<B_101%H6L<<IY;G1IN02 H.E24"P.N<$NW-7^PG#JD 
@5M5N^^0H-T$CIF#KHKL8D0 #P.G"^L] AL'=%JWUQ+0 
@[0_GM!D6$I<\WS733MKD2TIU%6#HG(G0$G'!*2[LMJD 
@]#L3HDC5,-:BQRD94A30U& 0@_8=1;>Z#K[$O^1I":( 
@#:>Q# 7R4[W%</5$T>]^DTE]A7KE+P(+DPQG-@*;+9D 
@?T.38,?(L6+<\?.\_T9J:1B,_4>[!QJ;'D$B:&:NE-L 
@?3(#'V8_8-"$D%GZ!ZFM_:MZ7UM#-:X</DR)@C;V>6H 
@]P]0IFR;'2@GR?B[E7:\(U/W%B+[84%8)-A&EA;G U4 
@(IIR8%3 X3X*U(@?ZA!P2&B&%V1.0Z?U,.ADI//M$B$ 
@D[?0!NLDKG/(0K^.$S5QB!H>,X+Y6;WQ^%8CO1M#PVL 
@_>\!7:2>)+"H!$%EM\<Z_!2$YW]\@HD)!BYSB"XE42H 
@(>1CCKEH\%\L2):>9?9-5AH-A'<4\;"K'KR@*99F/^@ 
@WTU#N#2%R;UK[?JN<,G#T:OB?Z /]MM1O#V1)QZ!'%< 
@ .M(*^J:(:?:V$=4?/RJJ^EF8 ===.GFQQRV9 9G/4, 
@!EV^NGK7^Z)NL2+H8UQ^/45J7 NP9*RNL2K[^C*3<Z$ 
@L8@;1^3IB( X#V:2D,&8BR5K'A<GDM?\70A(\:/8Y_0 
@K%">2FY\=*OR;(XW<X/KXM<Y0FD:QA0Y/W B<LB :#< 
@WOR%;LRH+3/?9")GUSK@+4V<FMSGF['NXU!O$1'[FQ8 
@J[-@IOO&=_!OU9KB]+*!!\Z\(V_HFI-E<I8VYKVA#2, 
@.H-T/^T;,WR/5C$8S2$26I3%YOY/R='H)'.'#,&:Q2T 
@,5$WJ?GH9H1,4^+/M9D9?@J9M04\4HM[TQTZ#F_0S @ 
@6SNUL'R2F']Y3 <KYNN03_ 7";ER&\<#LG;""TA*B$\ 
@E#32'BZ!8#$3=49FP*6HY*RZDN? XNNE,ZJDIQ''@-H 
@ W!"B$2^0S8Z_\^0]2CB/JRQ5V8+M0R3<10WYD;R0=  
@9,('$0+!>IB=%NT# F050 ^]](*1$S<W6]J*B#(:MY0 
@Y)V"GXMVNGR,'M[%2UBB)X?2#&0,_@3-+8>Q4 \72"H 
@I:,$,-@41.68>AZ>G?'HLHF, Z=K2"OSFZIQLI3OF5H 
@ Y9I8HN]S0:/N3D<WKI@.NKW=.M?^=:='+8?!O/3=Q@ 
@@_/7%OQF&VK&P/;&^NHP]ZT-VT/C)&Q4-SMN#.U4S/X 
@RE&YCQ6A]LJ0JQ(M2AETI) ,0T^2^#A14FMW82IH<:, 
@29BU -#[<YC41 E=Q#T[Y217G7-'9"J 4SSG$-V]XJX 
@Z9[XT#^/[0>ZCHFA<X(VO+JXZM+!H-1J+K+#P_  MD\ 
@EB[[SF_1.<SM?$K% ;M3GV-Z7LK^>;A42SY;JK,NAE< 
@_:5J_PV5(<I0='6RN 2I9E3.09\)]7 ( #H8:U98I^$ 
@KZD]/X?Y,1*W2.SNPO>"0EMR4-]=H3XW-T+PULLBT>H 
@$WM^&4?=!1K!?<P/&(CX_GB$"RCXS+*\*ZR)W9V>[;  
@Q!'MVZ PYOJ)"^)>ZDN%(4VM06?%BS+FX^O2\9RD"KT 
@1*\P<Z^X;YC3$VL_F($&_9GJSFGRS=POH(?N7:FO6(  
@/!.:K9_0Z]@RZ]QE&#E&8#[_']3VU=$.)0T&->!*MKX 
@E!]"O^^N4DH78!W+ %2Y*TT^+;H[%RM>NL G(1%5Q!P 
@!(Q#3YX?J#R\JW=4%1ASM"NS/[ 9JW9M&V77-[^:BG0 
@&R^[@NT3L%GX5DO9YAO?^MF=303A>WWW@30[7K4:P., 
@]E(8+("["6HV[@GT%\<DBF)3@=!O%]@%:V<50",[/;( 
@IS(=<^%Z Z#![<:LX1&_"HRV*>%<!, P*U(4O2;?M/, 
@I(IAZ ILEHD$Z9;/;Y$>>W9CB? 1@E"E!]HUGB= 8K, 
@1A/?F+Y'?%=+Q \$'8_OT)AI7W  6_LFN^A-FCVAS&< 
@K[9>OEQC7(M[CUW V.T3MFO;;*1@O.M^+QBQ5/#1:=8 
@*F[7I69V$F=\S@Y+]1*%7Y(-"@+.388_V Z46="8XT\ 
@7QZGU91JLVS(^*X9<'S(L]+WV ]15O(.D7%@.L1_G$\ 
@48MG&#\KB^/D#;[@O6PY3S!/9XAFB#\CU?="+@11U&, 
@(D>:J^@9Q,6==JLZQ VXN,7FPIE->)T->GT "^X;+1@ 
@5=0UO9FK-,=-A2VV,N6/3]C/_Y33#139*?B431!C>1, 
@AR:EC44D6$47ZP9&#=,V'N(I-1%B<O079(^P 4M,B ( 
@.=LKV19 R,9L8,I>OT-\>RD*077*7B1L>I9FC!#Z+=\ 
@-.8^EK8^.@LX\'BJM&9X:&EUAQB3N$,T<?^9NKA74'$ 
@_0&HN1A+MQ-)_"9JP1F@SH#H* 7!V0S?4:_#HI-(.)@ 
@4E03[ IVOKL7-;\.A%NKRRETV<H_] 8EQ6["5HZ4SXP 
@IQ%2Q0%&7HUSYU3/+J]0B!_%,HG"\-?@\#AI^N)\)4H 
@-0OFH^C6=-[2/$36MVM-NN@;^1&.>^VNFX98Y1VI\(@ 
@0"+P%36]2O:P>??W[*K>[E5S<974\"8,WG\.M)M0%5L 
@VZ1_<?US**W#!AMI&5/;<(RCBO14)0,BO>&4=/KA<Z$ 
@WB:(Q-;&Q6+)]5=N)__W0!BV6*'RL\4*F>\)*Z3\(R0 
@]O/)9=Y<B4)T; 85X]J9UC2^<!5#4>B]XZU0I<-0E/L 
@RFN;P=+X!L"ZIC<2H[.4<'S=9?3%@/B6Q #R.G(?,24 
@L+-F._+:M\&;R_)!Y"RO(N'$#E->RBQ(OM?1^XA$?)4 
@0A4M@EQT]MRF%BIN ^W[G1/AO>*&2G"5(Q/=<'J3M.D 
@6Z8")/:;2/D_'11ET5#UUL;=S&4:EH6XGI*+,2VFHD@ 
@4W;MRS['&-A6Y-]?AJ&5_3* D')A(0=39U-XUG=@CO@ 
0"TF"7BK.8I,DE<N5=R%YP0  
`pragma protect end_protected
