-- megafunction wizard: %Arria V Transceiver Native PHY v16.0%
-- GENERATION: XML
-- COLD_DATA_RxTx.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity COLD_DATA_RxTx is
	port (
		rx_analogreset          : in  std_logic_vector(7 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(7 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(7 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_is_lockedtoref       : out std_logic_vector(7 downto 0);                      --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_is_lockedtodata      : out std_logic_vector(7 downto 0);                      --      rx_is_lockedtodata.rx_is_lockedtodata
		rx_std_coreclkin        : in  std_logic_vector(7 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		rx_std_clkout           : out std_logic_vector(7 downto 0);                      --           rx_std_clkout.rx_std_clkout
		rx_cal_busy             : out std_logic_vector(7 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(559 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(367 downto 0);                    --      reconfig_from_xcvr.reconfig_from_xcvr
		rx_parallel_data        : out std_logic_vector(63 downto 0);                     --        rx_parallel_data.rx_parallel_data
		rx_datak                : out std_logic_vector(7 downto 0);                      --                rx_datak.rx_datak
		rx_errdetect            : out std_logic_vector(7 downto 0);                      --            rx_errdetect.rx_errdetect
		rx_disperr              : out std_logic_vector(7 downto 0);                      --              rx_disperr.rx_disperr
		rx_runningdisp          : out std_logic_vector(7 downto 0);                      --          rx_runningdisp.rx_runningdisp
		rx_patterndetect        : out std_logic_vector(7 downto 0);                      --        rx_patterndetect.rx_patterndetect
		rx_syncstatus           : out std_logic_vector(7 downto 0);                      --           rx_syncstatus.rx_syncstatus
		unused_rx_parallel_data : out std_logic_vector(399 downto 0)                     -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity COLD_DATA_RxTx;

architecture rtl of COLD_DATA_RxTx is
	component altera_xcvr_native_av is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 0;
			data_path_select                : string  := "pma_direct";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 80;
			tx_pma_clk_div                  : integer := 1;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pma_bonding_mode                : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0
		);
		port (
			rx_analogreset            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_is_lockedtoref         : out std_logic_vector(7 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(7 downto 0);                      -- rx_is_lockedtodata
			rx_std_coreclkin          : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			rx_std_clkout             : out std_logic_vector(7 downto 0);                      -- rx_std_clkout
			rx_cal_busy               : out std_logic_vector(7 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(559 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(367 downto 0);                    -- reconfig_from_xcvr
			rx_parallel_data          : out std_logic_vector(511 downto 0);                    -- unused_rx_parallel_data
			pll_powerdown             : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_pma_clkout             : out std_logic_vector(7 downto 0);                      -- tx_pma_clkout
			tx_serial_data            : out std_logic_vector(7 downto 0);                      -- tx_serial_data
			tx_pma_parallel_data      : in  std_logic_vector(639 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			pll_locked                : out std_logic_vector(7 downto 0);                      -- pll_locked
			ext_pll_clk               : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_pma_clkout             : out std_logic_vector(7 downto 0);                      -- rx_pma_clkout
			rx_pma_parallel_data      : out std_logic_vector(639 downto 0);                    -- rx_pma_parallel_data
			rx_clkslip                : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_clklow                 : out std_logic_vector(7 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(7 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_seriallpbken           : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_seriallpbken
			rx_signaldetect           : out std_logic_vector(7 downto 0);                      -- rx_signaldetect
			tx_parallel_data          : in  std_logic_vector(351 downto 0) := (others => 'X'); -- tx_parallel_data
			tx_std_coreclkin          : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(7 downto 0);                      -- tx_std_clkout
			rx_std_prbs_done          : out std_logic_vector(7 downto 0);                      -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(7 downto 0);                      -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(7 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(7 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(7 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(7 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(7 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(7 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(7 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(39 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(39 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(7 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_polinv             : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_std_elecidle           : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(7 downto 0);                      -- rx_std_signaldetect
			tx_cal_busy               : out std_logic_vector(7 downto 0)                       -- tx_cal_busy
		);
	end component altera_xcvr_native_av;

	signal cold_data_rxtx_inst_rx_parallel_data : std_logic_vector(511 downto 0); -- port fragment

begin

	cold_data_rxtx_inst : component altera_xcvr_native_av
		generic map (
			tx_enable                       => 0,
			rx_enable                       => 1,
			enable_std                      => 1,
			data_path_select                => "standard",
			channels                        => 8,
			bonded_mode                     => "non_bonded",
			data_rate                       => "1280 Mbps",
			pma_width                       => 10,
			tx_pma_clk_div                  => 1,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 1,
			pll_data_rate                   => "1280 Mbps",
			pll_type                        => "CMU",
			pma_bonding_mode                => "x1",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "unused",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "128.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 0,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 10,
			std_low_latency_bypass_enable   => 0,
			std_tx_pcfifo_mode              => "register_fifo",
			std_rx_pcfifo_mode              => "register_fifo",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 9,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 0,
			std_rx_byte_deser_enable        => 0,
			std_tx_8b10b_enable             => 1,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 1,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "sync_sm",
			std_rx_word_aligner_pattern_len => 10,
			std_rx_word_aligner_pattern     => "27C",
			std_rx_word_aligner_rknumber    => 5,
			std_rx_word_aligner_renumber    => 5,
			std_rx_word_aligner_rgnumber    => 5,
			std_rx_run_length_val           => 10,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 0,
			std_rx_polinv_enable            => 0
		)
		port map (
			rx_analogreset            => rx_analogreset,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset           => rx_digitalreset,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk             => rx_cdr_refclk,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data            => rx_serial_data,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_is_lockedtoref         => rx_is_lockedtoref,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata        => rx_is_lockedtodata,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			rx_std_coreclkin          => rx_std_coreclkin,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			rx_std_clkout             => rx_std_clkout,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      --      rx_std_clkout.rx_std_clkout
			rx_cal_busy               => rx_cal_busy,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr          => reconfig_to_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr        => reconfig_from_xcvr,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			rx_parallel_data(0)       => cold_data_rxtx_inst_rx_parallel_data(0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --   rx_parallel_data.rx_parallel_data
			rx_parallel_data(1)       => cold_data_rxtx_inst_rx_parallel_data(1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .rx_parallel_data
			rx_parallel_data(2)       => cold_data_rxtx_inst_rx_parallel_data(2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .rx_parallel_data
			rx_parallel_data(3)       => cold_data_rxtx_inst_rx_parallel_data(3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .rx_parallel_data
			rx_parallel_data(4)       => cold_data_rxtx_inst_rx_parallel_data(4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .rx_parallel_data
			rx_parallel_data(5)       => cold_data_rxtx_inst_rx_parallel_data(5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .rx_parallel_data
			rx_parallel_data(6)       => cold_data_rxtx_inst_rx_parallel_data(6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .rx_parallel_data
			rx_parallel_data(7)       => cold_data_rxtx_inst_rx_parallel_data(7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .rx_parallel_data
			rx_parallel_data(8)       => cold_data_rxtx_inst_rx_parallel_data(8),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .rx_parallel_data
			rx_parallel_data(9)       => cold_data_rxtx_inst_rx_parallel_data(9),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            --                   .rx_parallel_data
			rx_parallel_data(10)      => cold_data_rxtx_inst_rx_parallel_data(10),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(11)      => cold_data_rxtx_inst_rx_parallel_data(11),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(12)      => cold_data_rxtx_inst_rx_parallel_data(12),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(13)      => cold_data_rxtx_inst_rx_parallel_data(13),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(14)      => cold_data_rxtx_inst_rx_parallel_data(14),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(15)      => cold_data_rxtx_inst_rx_parallel_data(15),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(16)      => cold_data_rxtx_inst_rx_parallel_data(16),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(17)      => cold_data_rxtx_inst_rx_parallel_data(17),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(18)      => cold_data_rxtx_inst_rx_parallel_data(18),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(19)      => cold_data_rxtx_inst_rx_parallel_data(19),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(20)      => cold_data_rxtx_inst_rx_parallel_data(20),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(21)      => cold_data_rxtx_inst_rx_parallel_data(21),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(22)      => cold_data_rxtx_inst_rx_parallel_data(22),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(23)      => cold_data_rxtx_inst_rx_parallel_data(23),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(24)      => cold_data_rxtx_inst_rx_parallel_data(24),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(25)      => cold_data_rxtx_inst_rx_parallel_data(25),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(26)      => cold_data_rxtx_inst_rx_parallel_data(26),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(27)      => cold_data_rxtx_inst_rx_parallel_data(27),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(28)      => cold_data_rxtx_inst_rx_parallel_data(28),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(29)      => cold_data_rxtx_inst_rx_parallel_data(29),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(30)      => cold_data_rxtx_inst_rx_parallel_data(30),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(31)      => cold_data_rxtx_inst_rx_parallel_data(31),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(32)      => cold_data_rxtx_inst_rx_parallel_data(32),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(33)      => cold_data_rxtx_inst_rx_parallel_data(33),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(34)      => cold_data_rxtx_inst_rx_parallel_data(34),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(35)      => cold_data_rxtx_inst_rx_parallel_data(35),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(36)      => cold_data_rxtx_inst_rx_parallel_data(36),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(37)      => cold_data_rxtx_inst_rx_parallel_data(37),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(38)      => cold_data_rxtx_inst_rx_parallel_data(38),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(39)      => cold_data_rxtx_inst_rx_parallel_data(39),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(40)      => cold_data_rxtx_inst_rx_parallel_data(40),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(41)      => cold_data_rxtx_inst_rx_parallel_data(41),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(42)      => cold_data_rxtx_inst_rx_parallel_data(42),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(43)      => cold_data_rxtx_inst_rx_parallel_data(43),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(44)      => cold_data_rxtx_inst_rx_parallel_data(44),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(45)      => cold_data_rxtx_inst_rx_parallel_data(45),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(46)      => cold_data_rxtx_inst_rx_parallel_data(46),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(47)      => cold_data_rxtx_inst_rx_parallel_data(47),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(48)      => cold_data_rxtx_inst_rx_parallel_data(48),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(49)      => cold_data_rxtx_inst_rx_parallel_data(49),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(50)      => cold_data_rxtx_inst_rx_parallel_data(50),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(51)      => cold_data_rxtx_inst_rx_parallel_data(51),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(52)      => cold_data_rxtx_inst_rx_parallel_data(52),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(53)      => cold_data_rxtx_inst_rx_parallel_data(53),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(54)      => cold_data_rxtx_inst_rx_parallel_data(54),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(55)      => cold_data_rxtx_inst_rx_parallel_data(55),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(56)      => cold_data_rxtx_inst_rx_parallel_data(56),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(57)      => cold_data_rxtx_inst_rx_parallel_data(57),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(58)      => cold_data_rxtx_inst_rx_parallel_data(58),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(59)      => cold_data_rxtx_inst_rx_parallel_data(59),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(60)      => cold_data_rxtx_inst_rx_parallel_data(60),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(61)      => cold_data_rxtx_inst_rx_parallel_data(61),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(62)      => cold_data_rxtx_inst_rx_parallel_data(62),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(63)      => cold_data_rxtx_inst_rx_parallel_data(63),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(64)      => cold_data_rxtx_inst_rx_parallel_data(64),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(65)      => cold_data_rxtx_inst_rx_parallel_data(65),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(66)      => cold_data_rxtx_inst_rx_parallel_data(66),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(67)      => cold_data_rxtx_inst_rx_parallel_data(67),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(68)      => cold_data_rxtx_inst_rx_parallel_data(68),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(69)      => cold_data_rxtx_inst_rx_parallel_data(69),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(70)      => cold_data_rxtx_inst_rx_parallel_data(70),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(71)      => cold_data_rxtx_inst_rx_parallel_data(71),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(72)      => cold_data_rxtx_inst_rx_parallel_data(72),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(73)      => cold_data_rxtx_inst_rx_parallel_data(73),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(74)      => cold_data_rxtx_inst_rx_parallel_data(74),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(75)      => cold_data_rxtx_inst_rx_parallel_data(75),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(76)      => cold_data_rxtx_inst_rx_parallel_data(76),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(77)      => cold_data_rxtx_inst_rx_parallel_data(77),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(78)      => cold_data_rxtx_inst_rx_parallel_data(78),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(79)      => cold_data_rxtx_inst_rx_parallel_data(79),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(80)      => cold_data_rxtx_inst_rx_parallel_data(80),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(81)      => cold_data_rxtx_inst_rx_parallel_data(81),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(82)      => cold_data_rxtx_inst_rx_parallel_data(82),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(83)      => cold_data_rxtx_inst_rx_parallel_data(83),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(84)      => cold_data_rxtx_inst_rx_parallel_data(84),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(85)      => cold_data_rxtx_inst_rx_parallel_data(85),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(86)      => cold_data_rxtx_inst_rx_parallel_data(86),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(87)      => cold_data_rxtx_inst_rx_parallel_data(87),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(88)      => cold_data_rxtx_inst_rx_parallel_data(88),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(89)      => cold_data_rxtx_inst_rx_parallel_data(89),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(90)      => cold_data_rxtx_inst_rx_parallel_data(90),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(91)      => cold_data_rxtx_inst_rx_parallel_data(91),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(92)      => cold_data_rxtx_inst_rx_parallel_data(92),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(93)      => cold_data_rxtx_inst_rx_parallel_data(93),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(94)      => cold_data_rxtx_inst_rx_parallel_data(94),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(95)      => cold_data_rxtx_inst_rx_parallel_data(95),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(96)      => cold_data_rxtx_inst_rx_parallel_data(96),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(97)      => cold_data_rxtx_inst_rx_parallel_data(97),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(98)      => cold_data_rxtx_inst_rx_parallel_data(98),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(99)      => cold_data_rxtx_inst_rx_parallel_data(99),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           --                   .rx_parallel_data
			rx_parallel_data(100)     => cold_data_rxtx_inst_rx_parallel_data(100),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(101)     => cold_data_rxtx_inst_rx_parallel_data(101),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(102)     => cold_data_rxtx_inst_rx_parallel_data(102),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(103)     => cold_data_rxtx_inst_rx_parallel_data(103),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(104)     => cold_data_rxtx_inst_rx_parallel_data(104),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(105)     => cold_data_rxtx_inst_rx_parallel_data(105),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(106)     => cold_data_rxtx_inst_rx_parallel_data(106),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(107)     => cold_data_rxtx_inst_rx_parallel_data(107),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(108)     => cold_data_rxtx_inst_rx_parallel_data(108),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(109)     => cold_data_rxtx_inst_rx_parallel_data(109),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(110)     => cold_data_rxtx_inst_rx_parallel_data(110),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(111)     => cold_data_rxtx_inst_rx_parallel_data(111),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(112)     => cold_data_rxtx_inst_rx_parallel_data(112),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(113)     => cold_data_rxtx_inst_rx_parallel_data(113),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(114)     => cold_data_rxtx_inst_rx_parallel_data(114),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(115)     => cold_data_rxtx_inst_rx_parallel_data(115),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(116)     => cold_data_rxtx_inst_rx_parallel_data(116),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(117)     => cold_data_rxtx_inst_rx_parallel_data(117),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(118)     => cold_data_rxtx_inst_rx_parallel_data(118),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(119)     => cold_data_rxtx_inst_rx_parallel_data(119),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(120)     => cold_data_rxtx_inst_rx_parallel_data(120),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(121)     => cold_data_rxtx_inst_rx_parallel_data(121),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(122)     => cold_data_rxtx_inst_rx_parallel_data(122),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(123)     => cold_data_rxtx_inst_rx_parallel_data(123),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(124)     => cold_data_rxtx_inst_rx_parallel_data(124),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(125)     => cold_data_rxtx_inst_rx_parallel_data(125),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(126)     => cold_data_rxtx_inst_rx_parallel_data(126),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(127)     => cold_data_rxtx_inst_rx_parallel_data(127),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(128)     => cold_data_rxtx_inst_rx_parallel_data(128),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(129)     => cold_data_rxtx_inst_rx_parallel_data(129),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(130)     => cold_data_rxtx_inst_rx_parallel_data(130),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(131)     => cold_data_rxtx_inst_rx_parallel_data(131),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(132)     => cold_data_rxtx_inst_rx_parallel_data(132),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(133)     => cold_data_rxtx_inst_rx_parallel_data(133),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(134)     => cold_data_rxtx_inst_rx_parallel_data(134),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(135)     => cold_data_rxtx_inst_rx_parallel_data(135),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(136)     => cold_data_rxtx_inst_rx_parallel_data(136),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(137)     => cold_data_rxtx_inst_rx_parallel_data(137),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(138)     => cold_data_rxtx_inst_rx_parallel_data(138),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(139)     => cold_data_rxtx_inst_rx_parallel_data(139),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(140)     => cold_data_rxtx_inst_rx_parallel_data(140),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(141)     => cold_data_rxtx_inst_rx_parallel_data(141),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(142)     => cold_data_rxtx_inst_rx_parallel_data(142),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(143)     => cold_data_rxtx_inst_rx_parallel_data(143),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(144)     => cold_data_rxtx_inst_rx_parallel_data(144),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(145)     => cold_data_rxtx_inst_rx_parallel_data(145),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(146)     => cold_data_rxtx_inst_rx_parallel_data(146),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(147)     => cold_data_rxtx_inst_rx_parallel_data(147),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(148)     => cold_data_rxtx_inst_rx_parallel_data(148),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(149)     => cold_data_rxtx_inst_rx_parallel_data(149),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(150)     => cold_data_rxtx_inst_rx_parallel_data(150),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(151)     => cold_data_rxtx_inst_rx_parallel_data(151),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(152)     => cold_data_rxtx_inst_rx_parallel_data(152),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(153)     => cold_data_rxtx_inst_rx_parallel_data(153),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(154)     => cold_data_rxtx_inst_rx_parallel_data(154),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(155)     => cold_data_rxtx_inst_rx_parallel_data(155),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(156)     => cold_data_rxtx_inst_rx_parallel_data(156),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(157)     => cold_data_rxtx_inst_rx_parallel_data(157),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(158)     => cold_data_rxtx_inst_rx_parallel_data(158),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(159)     => cold_data_rxtx_inst_rx_parallel_data(159),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(160)     => cold_data_rxtx_inst_rx_parallel_data(160),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(161)     => cold_data_rxtx_inst_rx_parallel_data(161),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(162)     => cold_data_rxtx_inst_rx_parallel_data(162),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(163)     => cold_data_rxtx_inst_rx_parallel_data(163),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(164)     => cold_data_rxtx_inst_rx_parallel_data(164),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(165)     => cold_data_rxtx_inst_rx_parallel_data(165),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(166)     => cold_data_rxtx_inst_rx_parallel_data(166),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(167)     => cold_data_rxtx_inst_rx_parallel_data(167),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(168)     => cold_data_rxtx_inst_rx_parallel_data(168),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(169)     => cold_data_rxtx_inst_rx_parallel_data(169),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(170)     => cold_data_rxtx_inst_rx_parallel_data(170),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(171)     => cold_data_rxtx_inst_rx_parallel_data(171),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(172)     => cold_data_rxtx_inst_rx_parallel_data(172),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(173)     => cold_data_rxtx_inst_rx_parallel_data(173),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(174)     => cold_data_rxtx_inst_rx_parallel_data(174),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(175)     => cold_data_rxtx_inst_rx_parallel_data(175),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(176)     => cold_data_rxtx_inst_rx_parallel_data(176),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(177)     => cold_data_rxtx_inst_rx_parallel_data(177),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(178)     => cold_data_rxtx_inst_rx_parallel_data(178),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(179)     => cold_data_rxtx_inst_rx_parallel_data(179),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(180)     => cold_data_rxtx_inst_rx_parallel_data(180),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(181)     => cold_data_rxtx_inst_rx_parallel_data(181),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(182)     => cold_data_rxtx_inst_rx_parallel_data(182),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(183)     => cold_data_rxtx_inst_rx_parallel_data(183),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(184)     => cold_data_rxtx_inst_rx_parallel_data(184),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(185)     => cold_data_rxtx_inst_rx_parallel_data(185),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(186)     => cold_data_rxtx_inst_rx_parallel_data(186),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(187)     => cold_data_rxtx_inst_rx_parallel_data(187),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(188)     => cold_data_rxtx_inst_rx_parallel_data(188),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(189)     => cold_data_rxtx_inst_rx_parallel_data(189),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(190)     => cold_data_rxtx_inst_rx_parallel_data(190),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(191)     => cold_data_rxtx_inst_rx_parallel_data(191),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(192)     => cold_data_rxtx_inst_rx_parallel_data(192),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(193)     => cold_data_rxtx_inst_rx_parallel_data(193),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(194)     => cold_data_rxtx_inst_rx_parallel_data(194),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(195)     => cold_data_rxtx_inst_rx_parallel_data(195),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(196)     => cold_data_rxtx_inst_rx_parallel_data(196),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(197)     => cold_data_rxtx_inst_rx_parallel_data(197),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(198)     => cold_data_rxtx_inst_rx_parallel_data(198),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(199)     => cold_data_rxtx_inst_rx_parallel_data(199),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(200)     => cold_data_rxtx_inst_rx_parallel_data(200),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(201)     => cold_data_rxtx_inst_rx_parallel_data(201),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(202)     => cold_data_rxtx_inst_rx_parallel_data(202),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(203)     => cold_data_rxtx_inst_rx_parallel_data(203),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(204)     => cold_data_rxtx_inst_rx_parallel_data(204),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(205)     => cold_data_rxtx_inst_rx_parallel_data(205),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(206)     => cold_data_rxtx_inst_rx_parallel_data(206),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(207)     => cold_data_rxtx_inst_rx_parallel_data(207),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(208)     => cold_data_rxtx_inst_rx_parallel_data(208),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(209)     => cold_data_rxtx_inst_rx_parallel_data(209),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(210)     => cold_data_rxtx_inst_rx_parallel_data(210),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(211)     => cold_data_rxtx_inst_rx_parallel_data(211),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(212)     => cold_data_rxtx_inst_rx_parallel_data(212),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(213)     => cold_data_rxtx_inst_rx_parallel_data(213),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(214)     => cold_data_rxtx_inst_rx_parallel_data(214),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(215)     => cold_data_rxtx_inst_rx_parallel_data(215),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(216)     => cold_data_rxtx_inst_rx_parallel_data(216),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(217)     => cold_data_rxtx_inst_rx_parallel_data(217),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(218)     => cold_data_rxtx_inst_rx_parallel_data(218),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(219)     => cold_data_rxtx_inst_rx_parallel_data(219),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(220)     => cold_data_rxtx_inst_rx_parallel_data(220),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(221)     => cold_data_rxtx_inst_rx_parallel_data(221),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(222)     => cold_data_rxtx_inst_rx_parallel_data(222),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(223)     => cold_data_rxtx_inst_rx_parallel_data(223),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(224)     => cold_data_rxtx_inst_rx_parallel_data(224),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(225)     => cold_data_rxtx_inst_rx_parallel_data(225),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(226)     => cold_data_rxtx_inst_rx_parallel_data(226),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(227)     => cold_data_rxtx_inst_rx_parallel_data(227),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(228)     => cold_data_rxtx_inst_rx_parallel_data(228),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(229)     => cold_data_rxtx_inst_rx_parallel_data(229),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(230)     => cold_data_rxtx_inst_rx_parallel_data(230),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(231)     => cold_data_rxtx_inst_rx_parallel_data(231),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(232)     => cold_data_rxtx_inst_rx_parallel_data(232),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(233)     => cold_data_rxtx_inst_rx_parallel_data(233),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(234)     => cold_data_rxtx_inst_rx_parallel_data(234),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(235)     => cold_data_rxtx_inst_rx_parallel_data(235),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(236)     => cold_data_rxtx_inst_rx_parallel_data(236),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(237)     => cold_data_rxtx_inst_rx_parallel_data(237),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(238)     => cold_data_rxtx_inst_rx_parallel_data(238),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(239)     => cold_data_rxtx_inst_rx_parallel_data(239),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(240)     => cold_data_rxtx_inst_rx_parallel_data(240),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(241)     => cold_data_rxtx_inst_rx_parallel_data(241),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(242)     => cold_data_rxtx_inst_rx_parallel_data(242),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(243)     => cold_data_rxtx_inst_rx_parallel_data(243),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(244)     => cold_data_rxtx_inst_rx_parallel_data(244),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(245)     => cold_data_rxtx_inst_rx_parallel_data(245),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(246)     => cold_data_rxtx_inst_rx_parallel_data(246),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(247)     => cold_data_rxtx_inst_rx_parallel_data(247),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(248)     => cold_data_rxtx_inst_rx_parallel_data(248),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(249)     => cold_data_rxtx_inst_rx_parallel_data(249),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(250)     => cold_data_rxtx_inst_rx_parallel_data(250),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(251)     => cold_data_rxtx_inst_rx_parallel_data(251),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(252)     => cold_data_rxtx_inst_rx_parallel_data(252),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(253)     => cold_data_rxtx_inst_rx_parallel_data(253),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(254)     => cold_data_rxtx_inst_rx_parallel_data(254),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(255)     => cold_data_rxtx_inst_rx_parallel_data(255),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(256)     => cold_data_rxtx_inst_rx_parallel_data(256),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(257)     => cold_data_rxtx_inst_rx_parallel_data(257),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(258)     => cold_data_rxtx_inst_rx_parallel_data(258),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(259)     => cold_data_rxtx_inst_rx_parallel_data(259),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(260)     => cold_data_rxtx_inst_rx_parallel_data(260),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(261)     => cold_data_rxtx_inst_rx_parallel_data(261),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(262)     => cold_data_rxtx_inst_rx_parallel_data(262),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(263)     => cold_data_rxtx_inst_rx_parallel_data(263),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(264)     => cold_data_rxtx_inst_rx_parallel_data(264),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(265)     => cold_data_rxtx_inst_rx_parallel_data(265),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(266)     => cold_data_rxtx_inst_rx_parallel_data(266),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(267)     => cold_data_rxtx_inst_rx_parallel_data(267),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(268)     => cold_data_rxtx_inst_rx_parallel_data(268),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(269)     => cold_data_rxtx_inst_rx_parallel_data(269),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(270)     => cold_data_rxtx_inst_rx_parallel_data(270),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(271)     => cold_data_rxtx_inst_rx_parallel_data(271),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(272)     => cold_data_rxtx_inst_rx_parallel_data(272),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(273)     => cold_data_rxtx_inst_rx_parallel_data(273),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(274)     => cold_data_rxtx_inst_rx_parallel_data(274),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(275)     => cold_data_rxtx_inst_rx_parallel_data(275),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(276)     => cold_data_rxtx_inst_rx_parallel_data(276),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(277)     => cold_data_rxtx_inst_rx_parallel_data(277),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(278)     => cold_data_rxtx_inst_rx_parallel_data(278),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(279)     => cold_data_rxtx_inst_rx_parallel_data(279),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(280)     => cold_data_rxtx_inst_rx_parallel_data(280),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(281)     => cold_data_rxtx_inst_rx_parallel_data(281),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(282)     => cold_data_rxtx_inst_rx_parallel_data(282),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(283)     => cold_data_rxtx_inst_rx_parallel_data(283),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(284)     => cold_data_rxtx_inst_rx_parallel_data(284),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(285)     => cold_data_rxtx_inst_rx_parallel_data(285),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(286)     => cold_data_rxtx_inst_rx_parallel_data(286),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(287)     => cold_data_rxtx_inst_rx_parallel_data(287),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(288)     => cold_data_rxtx_inst_rx_parallel_data(288),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(289)     => cold_data_rxtx_inst_rx_parallel_data(289),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(290)     => cold_data_rxtx_inst_rx_parallel_data(290),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(291)     => cold_data_rxtx_inst_rx_parallel_data(291),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(292)     => cold_data_rxtx_inst_rx_parallel_data(292),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(293)     => cold_data_rxtx_inst_rx_parallel_data(293),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(294)     => cold_data_rxtx_inst_rx_parallel_data(294),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(295)     => cold_data_rxtx_inst_rx_parallel_data(295),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(296)     => cold_data_rxtx_inst_rx_parallel_data(296),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(297)     => cold_data_rxtx_inst_rx_parallel_data(297),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(298)     => cold_data_rxtx_inst_rx_parallel_data(298),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(299)     => cold_data_rxtx_inst_rx_parallel_data(299),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(300)     => cold_data_rxtx_inst_rx_parallel_data(300),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(301)     => cold_data_rxtx_inst_rx_parallel_data(301),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(302)     => cold_data_rxtx_inst_rx_parallel_data(302),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(303)     => cold_data_rxtx_inst_rx_parallel_data(303),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(304)     => cold_data_rxtx_inst_rx_parallel_data(304),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(305)     => cold_data_rxtx_inst_rx_parallel_data(305),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(306)     => cold_data_rxtx_inst_rx_parallel_data(306),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(307)     => cold_data_rxtx_inst_rx_parallel_data(307),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(308)     => cold_data_rxtx_inst_rx_parallel_data(308),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(309)     => cold_data_rxtx_inst_rx_parallel_data(309),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(310)     => cold_data_rxtx_inst_rx_parallel_data(310),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(311)     => cold_data_rxtx_inst_rx_parallel_data(311),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(312)     => cold_data_rxtx_inst_rx_parallel_data(312),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(313)     => cold_data_rxtx_inst_rx_parallel_data(313),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(314)     => cold_data_rxtx_inst_rx_parallel_data(314),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(315)     => cold_data_rxtx_inst_rx_parallel_data(315),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(316)     => cold_data_rxtx_inst_rx_parallel_data(316),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(317)     => cold_data_rxtx_inst_rx_parallel_data(317),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(318)     => cold_data_rxtx_inst_rx_parallel_data(318),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(319)     => cold_data_rxtx_inst_rx_parallel_data(319),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(320)     => cold_data_rxtx_inst_rx_parallel_data(320),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(321)     => cold_data_rxtx_inst_rx_parallel_data(321),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(322)     => cold_data_rxtx_inst_rx_parallel_data(322),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(323)     => cold_data_rxtx_inst_rx_parallel_data(323),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(324)     => cold_data_rxtx_inst_rx_parallel_data(324),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(325)     => cold_data_rxtx_inst_rx_parallel_data(325),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(326)     => cold_data_rxtx_inst_rx_parallel_data(326),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(327)     => cold_data_rxtx_inst_rx_parallel_data(327),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(328)     => cold_data_rxtx_inst_rx_parallel_data(328),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(329)     => cold_data_rxtx_inst_rx_parallel_data(329),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(330)     => cold_data_rxtx_inst_rx_parallel_data(330),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(331)     => cold_data_rxtx_inst_rx_parallel_data(331),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(332)     => cold_data_rxtx_inst_rx_parallel_data(332),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(333)     => cold_data_rxtx_inst_rx_parallel_data(333),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(334)     => cold_data_rxtx_inst_rx_parallel_data(334),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(335)     => cold_data_rxtx_inst_rx_parallel_data(335),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(336)     => cold_data_rxtx_inst_rx_parallel_data(336),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(337)     => cold_data_rxtx_inst_rx_parallel_data(337),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(338)     => cold_data_rxtx_inst_rx_parallel_data(338),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(339)     => cold_data_rxtx_inst_rx_parallel_data(339),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(340)     => cold_data_rxtx_inst_rx_parallel_data(340),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(341)     => cold_data_rxtx_inst_rx_parallel_data(341),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(342)     => cold_data_rxtx_inst_rx_parallel_data(342),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(343)     => cold_data_rxtx_inst_rx_parallel_data(343),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(344)     => cold_data_rxtx_inst_rx_parallel_data(344),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(345)     => cold_data_rxtx_inst_rx_parallel_data(345),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(346)     => cold_data_rxtx_inst_rx_parallel_data(346),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(347)     => cold_data_rxtx_inst_rx_parallel_data(347),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(348)     => cold_data_rxtx_inst_rx_parallel_data(348),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(349)     => cold_data_rxtx_inst_rx_parallel_data(349),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(350)     => cold_data_rxtx_inst_rx_parallel_data(350),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(351)     => cold_data_rxtx_inst_rx_parallel_data(351),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(352)     => cold_data_rxtx_inst_rx_parallel_data(352),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(353)     => cold_data_rxtx_inst_rx_parallel_data(353),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(354)     => cold_data_rxtx_inst_rx_parallel_data(354),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(355)     => cold_data_rxtx_inst_rx_parallel_data(355),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(356)     => cold_data_rxtx_inst_rx_parallel_data(356),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(357)     => cold_data_rxtx_inst_rx_parallel_data(357),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(358)     => cold_data_rxtx_inst_rx_parallel_data(358),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(359)     => cold_data_rxtx_inst_rx_parallel_data(359),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(360)     => cold_data_rxtx_inst_rx_parallel_data(360),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(361)     => cold_data_rxtx_inst_rx_parallel_data(361),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(362)     => cold_data_rxtx_inst_rx_parallel_data(362),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(363)     => cold_data_rxtx_inst_rx_parallel_data(363),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(364)     => cold_data_rxtx_inst_rx_parallel_data(364),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(365)     => cold_data_rxtx_inst_rx_parallel_data(365),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(366)     => cold_data_rxtx_inst_rx_parallel_data(366),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(367)     => cold_data_rxtx_inst_rx_parallel_data(367),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(368)     => cold_data_rxtx_inst_rx_parallel_data(368),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(369)     => cold_data_rxtx_inst_rx_parallel_data(369),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(370)     => cold_data_rxtx_inst_rx_parallel_data(370),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(371)     => cold_data_rxtx_inst_rx_parallel_data(371),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(372)     => cold_data_rxtx_inst_rx_parallel_data(372),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(373)     => cold_data_rxtx_inst_rx_parallel_data(373),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(374)     => cold_data_rxtx_inst_rx_parallel_data(374),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(375)     => cold_data_rxtx_inst_rx_parallel_data(375),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(376)     => cold_data_rxtx_inst_rx_parallel_data(376),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(377)     => cold_data_rxtx_inst_rx_parallel_data(377),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(378)     => cold_data_rxtx_inst_rx_parallel_data(378),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(379)     => cold_data_rxtx_inst_rx_parallel_data(379),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(380)     => cold_data_rxtx_inst_rx_parallel_data(380),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(381)     => cold_data_rxtx_inst_rx_parallel_data(381),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(382)     => cold_data_rxtx_inst_rx_parallel_data(382),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(383)     => cold_data_rxtx_inst_rx_parallel_data(383),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(384)     => cold_data_rxtx_inst_rx_parallel_data(384),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(385)     => cold_data_rxtx_inst_rx_parallel_data(385),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(386)     => cold_data_rxtx_inst_rx_parallel_data(386),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(387)     => cold_data_rxtx_inst_rx_parallel_data(387),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(388)     => cold_data_rxtx_inst_rx_parallel_data(388),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(389)     => cold_data_rxtx_inst_rx_parallel_data(389),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(390)     => cold_data_rxtx_inst_rx_parallel_data(390),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(391)     => cold_data_rxtx_inst_rx_parallel_data(391),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(392)     => cold_data_rxtx_inst_rx_parallel_data(392),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(393)     => cold_data_rxtx_inst_rx_parallel_data(393),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(394)     => cold_data_rxtx_inst_rx_parallel_data(394),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(395)     => cold_data_rxtx_inst_rx_parallel_data(395),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(396)     => cold_data_rxtx_inst_rx_parallel_data(396),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(397)     => cold_data_rxtx_inst_rx_parallel_data(397),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(398)     => cold_data_rxtx_inst_rx_parallel_data(398),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(399)     => cold_data_rxtx_inst_rx_parallel_data(399),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(400)     => cold_data_rxtx_inst_rx_parallel_data(400),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(401)     => cold_data_rxtx_inst_rx_parallel_data(401),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(402)     => cold_data_rxtx_inst_rx_parallel_data(402),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(403)     => cold_data_rxtx_inst_rx_parallel_data(403),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(404)     => cold_data_rxtx_inst_rx_parallel_data(404),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(405)     => cold_data_rxtx_inst_rx_parallel_data(405),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(406)     => cold_data_rxtx_inst_rx_parallel_data(406),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(407)     => cold_data_rxtx_inst_rx_parallel_data(407),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(408)     => cold_data_rxtx_inst_rx_parallel_data(408),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(409)     => cold_data_rxtx_inst_rx_parallel_data(409),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(410)     => cold_data_rxtx_inst_rx_parallel_data(410),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(411)     => cold_data_rxtx_inst_rx_parallel_data(411),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(412)     => cold_data_rxtx_inst_rx_parallel_data(412),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(413)     => cold_data_rxtx_inst_rx_parallel_data(413),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(414)     => cold_data_rxtx_inst_rx_parallel_data(414),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(415)     => cold_data_rxtx_inst_rx_parallel_data(415),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(416)     => cold_data_rxtx_inst_rx_parallel_data(416),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(417)     => cold_data_rxtx_inst_rx_parallel_data(417),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(418)     => cold_data_rxtx_inst_rx_parallel_data(418),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(419)     => cold_data_rxtx_inst_rx_parallel_data(419),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(420)     => cold_data_rxtx_inst_rx_parallel_data(420),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(421)     => cold_data_rxtx_inst_rx_parallel_data(421),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(422)     => cold_data_rxtx_inst_rx_parallel_data(422),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(423)     => cold_data_rxtx_inst_rx_parallel_data(423),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(424)     => cold_data_rxtx_inst_rx_parallel_data(424),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(425)     => cold_data_rxtx_inst_rx_parallel_data(425),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(426)     => cold_data_rxtx_inst_rx_parallel_data(426),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(427)     => cold_data_rxtx_inst_rx_parallel_data(427),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(428)     => cold_data_rxtx_inst_rx_parallel_data(428),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(429)     => cold_data_rxtx_inst_rx_parallel_data(429),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(430)     => cold_data_rxtx_inst_rx_parallel_data(430),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(431)     => cold_data_rxtx_inst_rx_parallel_data(431),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(432)     => cold_data_rxtx_inst_rx_parallel_data(432),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(433)     => cold_data_rxtx_inst_rx_parallel_data(433),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(434)     => cold_data_rxtx_inst_rx_parallel_data(434),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(435)     => cold_data_rxtx_inst_rx_parallel_data(435),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(436)     => cold_data_rxtx_inst_rx_parallel_data(436),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(437)     => cold_data_rxtx_inst_rx_parallel_data(437),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(438)     => cold_data_rxtx_inst_rx_parallel_data(438),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(439)     => cold_data_rxtx_inst_rx_parallel_data(439),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(440)     => cold_data_rxtx_inst_rx_parallel_data(440),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(441)     => cold_data_rxtx_inst_rx_parallel_data(441),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(442)     => cold_data_rxtx_inst_rx_parallel_data(442),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(443)     => cold_data_rxtx_inst_rx_parallel_data(443),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(444)     => cold_data_rxtx_inst_rx_parallel_data(444),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(445)     => cold_data_rxtx_inst_rx_parallel_data(445),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(446)     => cold_data_rxtx_inst_rx_parallel_data(446),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(447)     => cold_data_rxtx_inst_rx_parallel_data(447),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(448)     => cold_data_rxtx_inst_rx_parallel_data(448),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(449)     => cold_data_rxtx_inst_rx_parallel_data(449),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(450)     => cold_data_rxtx_inst_rx_parallel_data(450),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(451)     => cold_data_rxtx_inst_rx_parallel_data(451),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(452)     => cold_data_rxtx_inst_rx_parallel_data(452),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(453)     => cold_data_rxtx_inst_rx_parallel_data(453),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(454)     => cold_data_rxtx_inst_rx_parallel_data(454),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(455)     => cold_data_rxtx_inst_rx_parallel_data(455),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(456)     => cold_data_rxtx_inst_rx_parallel_data(456),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(457)     => cold_data_rxtx_inst_rx_parallel_data(457),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(458)     => cold_data_rxtx_inst_rx_parallel_data(458),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(459)     => cold_data_rxtx_inst_rx_parallel_data(459),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(460)     => cold_data_rxtx_inst_rx_parallel_data(460),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(461)     => cold_data_rxtx_inst_rx_parallel_data(461),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(462)     => cold_data_rxtx_inst_rx_parallel_data(462),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(463)     => cold_data_rxtx_inst_rx_parallel_data(463),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(464)     => cold_data_rxtx_inst_rx_parallel_data(464),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(465)     => cold_data_rxtx_inst_rx_parallel_data(465),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(466)     => cold_data_rxtx_inst_rx_parallel_data(466),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(467)     => cold_data_rxtx_inst_rx_parallel_data(467),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(468)     => cold_data_rxtx_inst_rx_parallel_data(468),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(469)     => cold_data_rxtx_inst_rx_parallel_data(469),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(470)     => cold_data_rxtx_inst_rx_parallel_data(470),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(471)     => cold_data_rxtx_inst_rx_parallel_data(471),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(472)     => cold_data_rxtx_inst_rx_parallel_data(472),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(473)     => cold_data_rxtx_inst_rx_parallel_data(473),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(474)     => cold_data_rxtx_inst_rx_parallel_data(474),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(475)     => cold_data_rxtx_inst_rx_parallel_data(475),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(476)     => cold_data_rxtx_inst_rx_parallel_data(476),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(477)     => cold_data_rxtx_inst_rx_parallel_data(477),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(478)     => cold_data_rxtx_inst_rx_parallel_data(478),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(479)     => cold_data_rxtx_inst_rx_parallel_data(479),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(480)     => cold_data_rxtx_inst_rx_parallel_data(480),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(481)     => cold_data_rxtx_inst_rx_parallel_data(481),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(482)     => cold_data_rxtx_inst_rx_parallel_data(482),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(483)     => cold_data_rxtx_inst_rx_parallel_data(483),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(484)     => cold_data_rxtx_inst_rx_parallel_data(484),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(485)     => cold_data_rxtx_inst_rx_parallel_data(485),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(486)     => cold_data_rxtx_inst_rx_parallel_data(486),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(487)     => cold_data_rxtx_inst_rx_parallel_data(487),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(488)     => cold_data_rxtx_inst_rx_parallel_data(488),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(489)     => cold_data_rxtx_inst_rx_parallel_data(489),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(490)     => cold_data_rxtx_inst_rx_parallel_data(490),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(491)     => cold_data_rxtx_inst_rx_parallel_data(491),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(492)     => cold_data_rxtx_inst_rx_parallel_data(492),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(493)     => cold_data_rxtx_inst_rx_parallel_data(493),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(494)     => cold_data_rxtx_inst_rx_parallel_data(494),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(495)     => cold_data_rxtx_inst_rx_parallel_data(495),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(496)     => cold_data_rxtx_inst_rx_parallel_data(496),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(497)     => cold_data_rxtx_inst_rx_parallel_data(497),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(498)     => cold_data_rxtx_inst_rx_parallel_data(498),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(499)     => cold_data_rxtx_inst_rx_parallel_data(499),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(500)     => cold_data_rxtx_inst_rx_parallel_data(500),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(501)     => cold_data_rxtx_inst_rx_parallel_data(501),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(502)     => cold_data_rxtx_inst_rx_parallel_data(502),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(503)     => cold_data_rxtx_inst_rx_parallel_data(503),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(504)     => cold_data_rxtx_inst_rx_parallel_data(504),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(505)     => cold_data_rxtx_inst_rx_parallel_data(505),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(506)     => cold_data_rxtx_inst_rx_parallel_data(506),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(507)     => cold_data_rxtx_inst_rx_parallel_data(507),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(508)     => cold_data_rxtx_inst_rx_parallel_data(508),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(509)     => cold_data_rxtx_inst_rx_parallel_data(509),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(510)     => cold_data_rxtx_inst_rx_parallel_data(510),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			rx_parallel_data(511)     => cold_data_rxtx_inst_rx_parallel_data(511),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          --                   .rx_parallel_data
			pll_powerdown             => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			tx_analogreset            => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			tx_digitalreset           => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			tx_pll_refclk             => "0",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
			tx_pma_clkout             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_serial_data            => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_parallel_data      => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			pll_locked                => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			ext_pll_clk               => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_pma_clkout             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_parallel_data      => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_clkslip                => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_clklow                 => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_fref                   => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_set_locktodata         => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_set_locktoref          => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_seriallpbken           => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_signaldetect           => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_parallel_data          => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                 --        (terminated)
			tx_std_coreclkin          => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			tx_std_clkout             => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_done          => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_err           => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_byteorder_ena      => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_std_byteorder_flag     => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_full        => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign    => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_std_wa_a1a2size        => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			tx_std_bitslipboundarysel => "0000000000000000000000000000000000000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_std_bitslipboundarysel => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitslip            => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_std_runlength_err      => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena         => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_std_byterev_ena        => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			tx_std_polinv             => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_std_polinv             => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			tx_std_elecidle           => "00000000",                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         --        (terminated)
			rx_std_signaldetect       => open,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_cal_busy               => open                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --        (terminated)
		);

	rx_errdetect <= COLD_DATA_RxTx_inst_rx_parallel_data(457) & COLD_DATA_RxTx_inst_rx_parallel_data(393) & COLD_DATA_RxTx_inst_rx_parallel_data(329) & COLD_DATA_RxTx_inst_rx_parallel_data(265) & COLD_DATA_RxTx_inst_rx_parallel_data(201) & COLD_DATA_RxTx_inst_rx_parallel_data(137) & COLD_DATA_RxTx_inst_rx_parallel_data(73) & COLD_DATA_RxTx_inst_rx_parallel_data(9);

	rx_parallel_data <= COLD_DATA_RxTx_inst_rx_parallel_data(455) & COLD_DATA_RxTx_inst_rx_parallel_data(454) & COLD_DATA_RxTx_inst_rx_parallel_data(453) & COLD_DATA_RxTx_inst_rx_parallel_data(452) & COLD_DATA_RxTx_inst_rx_parallel_data(451) & COLD_DATA_RxTx_inst_rx_parallel_data(450) & COLD_DATA_RxTx_inst_rx_parallel_data(449) & COLD_DATA_RxTx_inst_rx_parallel_data(448) & COLD_DATA_RxTx_inst_rx_parallel_data(391) & COLD_DATA_RxTx_inst_rx_parallel_data(390) & COLD_DATA_RxTx_inst_rx_parallel_data(389) & COLD_DATA_RxTx_inst_rx_parallel_data(388) & COLD_DATA_RxTx_inst_rx_parallel_data(387) & COLD_DATA_RxTx_inst_rx_parallel_data(386) & COLD_DATA_RxTx_inst_rx_parallel_data(385) & COLD_DATA_RxTx_inst_rx_parallel_data(384) & COLD_DATA_RxTx_inst_rx_parallel_data(327) & COLD_DATA_RxTx_inst_rx_parallel_data(326) & COLD_DATA_RxTx_inst_rx_parallel_data(325) & COLD_DATA_RxTx_inst_rx_parallel_data(324) & COLD_DATA_RxTx_inst_rx_parallel_data(323) & COLD_DATA_RxTx_inst_rx_parallel_data(322) & COLD_DATA_RxTx_inst_rx_parallel_data(321) & COLD_DATA_RxTx_inst_rx_parallel_data(320) & COLD_DATA_RxTx_inst_rx_parallel_data(263) & COLD_DATA_RxTx_inst_rx_parallel_data(262) & COLD_DATA_RxTx_inst_rx_parallel_data(261) & COLD_DATA_RxTx_inst_rx_parallel_data(260) & COLD_DATA_RxTx_inst_rx_parallel_data(259) & COLD_DATA_RxTx_inst_rx_parallel_data(258) & COLD_DATA_RxTx_inst_rx_parallel_data(257) & COLD_DATA_RxTx_inst_rx_parallel_data(256) & COLD_DATA_RxTx_inst_rx_parallel_data(199) & COLD_DATA_RxTx_inst_rx_parallel_data(198) & COLD_DATA_RxTx_inst_rx_parallel_data(197) & COLD_DATA_RxTx_inst_rx_parallel_data(196) & COLD_DATA_RxTx_inst_rx_parallel_data(195) & COLD_DATA_RxTx_inst_rx_parallel_data(194) & COLD_DATA_RxTx_inst_rx_parallel_data(193) & COLD_DATA_RxTx_inst_rx_parallel_data(192) & COLD_DATA_RxTx_inst_rx_parallel_data(135) & COLD_DATA_RxTx_inst_rx_parallel_data(134) & COLD_DATA_RxTx_inst_rx_parallel_data(133) & COLD_DATA_RxTx_inst_rx_parallel_data(132) & COLD_DATA_RxTx_inst_rx_parallel_data(131) & COLD_DATA_RxTx_inst_rx_parallel_data(130) & COLD_DATA_RxTx_inst_rx_parallel_data(129) & COLD_DATA_RxTx_inst_rx_parallel_data(128) & COLD_DATA_RxTx_inst_rx_parallel_data(71) & COLD_DATA_RxTx_inst_rx_parallel_data(70) & COLD_DATA_RxTx_inst_rx_parallel_data(69) & COLD_DATA_RxTx_inst_rx_parallel_data(68) & COLD_DATA_RxTx_inst_rx_parallel_data(67) & COLD_DATA_RxTx_inst_rx_parallel_data(66) & COLD_DATA_RxTx_inst_rx_parallel_data(65) & COLD_DATA_RxTx_inst_rx_parallel_data(64) & COLD_DATA_RxTx_inst_rx_parallel_data(7) & COLD_DATA_RxTx_inst_rx_parallel_data(6) & COLD_DATA_RxTx_inst_rx_parallel_data(5) & COLD_DATA_RxTx_inst_rx_parallel_data(4) & COLD_DATA_RxTx_inst_rx_parallel_data(3) & COLD_DATA_RxTx_inst_rx_parallel_data(2) & COLD_DATA_RxTx_inst_rx_parallel_data(1) & COLD_DATA_RxTx_inst_rx_parallel_data(0);

	rx_datak <= COLD_DATA_RxTx_inst_rx_parallel_data(456) & COLD_DATA_RxTx_inst_rx_parallel_data(392) & COLD_DATA_RxTx_inst_rx_parallel_data(328) & COLD_DATA_RxTx_inst_rx_parallel_data(264) & COLD_DATA_RxTx_inst_rx_parallel_data(200) & COLD_DATA_RxTx_inst_rx_parallel_data(136) & COLD_DATA_RxTx_inst_rx_parallel_data(72) & COLD_DATA_RxTx_inst_rx_parallel_data(8);

	rx_disperr <= COLD_DATA_RxTx_inst_rx_parallel_data(459) & COLD_DATA_RxTx_inst_rx_parallel_data(395) & COLD_DATA_RxTx_inst_rx_parallel_data(331) & COLD_DATA_RxTx_inst_rx_parallel_data(267) & COLD_DATA_RxTx_inst_rx_parallel_data(203) & COLD_DATA_RxTx_inst_rx_parallel_data(139) & COLD_DATA_RxTx_inst_rx_parallel_data(75) & COLD_DATA_RxTx_inst_rx_parallel_data(11);

	unused_rx_parallel_data <= COLD_DATA_RxTx_inst_rx_parallel_data(511) & COLD_DATA_RxTx_inst_rx_parallel_data(510) & COLD_DATA_RxTx_inst_rx_parallel_data(509) & COLD_DATA_RxTx_inst_rx_parallel_data(508) & COLD_DATA_RxTx_inst_rx_parallel_data(507) & COLD_DATA_RxTx_inst_rx_parallel_data(506) & COLD_DATA_RxTx_inst_rx_parallel_data(505) & COLD_DATA_RxTx_inst_rx_parallel_data(504) & COLD_DATA_RxTx_inst_rx_parallel_data(503) & COLD_DATA_RxTx_inst_rx_parallel_data(502) & COLD_DATA_RxTx_inst_rx_parallel_data(501) & COLD_DATA_RxTx_inst_rx_parallel_data(500) & COLD_DATA_RxTx_inst_rx_parallel_data(499) & COLD_DATA_RxTx_inst_rx_parallel_data(498) & COLD_DATA_RxTx_inst_rx_parallel_data(497) & COLD_DATA_RxTx_inst_rx_parallel_data(496) & COLD_DATA_RxTx_inst_rx_parallel_data(495) & COLD_DATA_RxTx_inst_rx_parallel_data(494) & COLD_DATA_RxTx_inst_rx_parallel_data(493) & COLD_DATA_RxTx_inst_rx_parallel_data(492) & COLD_DATA_RxTx_inst_rx_parallel_data(491) & COLD_DATA_RxTx_inst_rx_parallel_data(490) & COLD_DATA_RxTx_inst_rx_parallel_data(489) & COLD_DATA_RxTx_inst_rx_parallel_data(488) & COLD_DATA_RxTx_inst_rx_parallel_data(487) & COLD_DATA_RxTx_inst_rx_parallel_data(486) & COLD_DATA_RxTx_inst_rx_parallel_data(485) & COLD_DATA_RxTx_inst_rx_parallel_data(484) & COLD_DATA_RxTx_inst_rx_parallel_data(483) & COLD_DATA_RxTx_inst_rx_parallel_data(482) & COLD_DATA_RxTx_inst_rx_parallel_data(481) & COLD_DATA_RxTx_inst_rx_parallel_data(480) & COLD_DATA_RxTx_inst_rx_parallel_data(479) & COLD_DATA_RxTx_inst_rx_parallel_data(478) & COLD_DATA_RxTx_inst_rx_parallel_data(477) & COLD_DATA_RxTx_inst_rx_parallel_data(476) & COLD_DATA_RxTx_inst_rx_parallel_data(475) & COLD_DATA_RxTx_inst_rx_parallel_data(474) & COLD_DATA_RxTx_inst_rx_parallel_data(473) & COLD_DATA_RxTx_inst_rx_parallel_data(472) & COLD_DATA_RxTx_inst_rx_parallel_data(471) & COLD_DATA_RxTx_inst_rx_parallel_data(470) & COLD_DATA_RxTx_inst_rx_parallel_data(469) & COLD_DATA_RxTx_inst_rx_parallel_data(468) & COLD_DATA_RxTx_inst_rx_parallel_data(467) & COLD_DATA_RxTx_inst_rx_parallel_data(466) & COLD_DATA_RxTx_inst_rx_parallel_data(465) & COLD_DATA_RxTx_inst_rx_parallel_data(464) & COLD_DATA_RxTx_inst_rx_parallel_data(462) & COLD_DATA_RxTx_inst_rx_parallel_data(461) & COLD_DATA_RxTx_inst_rx_parallel_data(447) & COLD_DATA_RxTx_inst_rx_parallel_data(446) & COLD_DATA_RxTx_inst_rx_parallel_data(445) & COLD_DATA_RxTx_inst_rx_parallel_data(444) & COLD_DATA_RxTx_inst_rx_parallel_data(443) & COLD_DATA_RxTx_inst_rx_parallel_data(442) & COLD_DATA_RxTx_inst_rx_parallel_data(441) & COLD_DATA_RxTx_inst_rx_parallel_data(440) & COLD_DATA_RxTx_inst_rx_parallel_data(439) & COLD_DATA_RxTx_inst_rx_parallel_data(438) & COLD_DATA_RxTx_inst_rx_parallel_data(437) & COLD_DATA_RxTx_inst_rx_parallel_data(436) & COLD_DATA_RxTx_inst_rx_parallel_data(435) & COLD_DATA_RxTx_inst_rx_parallel_data(434) & COLD_DATA_RxTx_inst_rx_parallel_data(433) & COLD_DATA_RxTx_inst_rx_parallel_data(432) & COLD_DATA_RxTx_inst_rx_parallel_data(431) & COLD_DATA_RxTx_inst_rx_parallel_data(430) & COLD_DATA_RxTx_inst_rx_parallel_data(429) & COLD_DATA_RxTx_inst_rx_parallel_data(428) & COLD_DATA_RxTx_inst_rx_parallel_data(427) & COLD_DATA_RxTx_inst_rx_parallel_data(426) & COLD_DATA_RxTx_inst_rx_parallel_data(425) & COLD_DATA_RxTx_inst_rx_parallel_data(424) & COLD_DATA_RxTx_inst_rx_parallel_data(423) & COLD_DATA_RxTx_inst_rx_parallel_data(422) & COLD_DATA_RxTx_inst_rx_parallel_data(421) & COLD_DATA_RxTx_inst_rx_parallel_data(420) & COLD_DATA_RxTx_inst_rx_parallel_data(419) & COLD_DATA_RxTx_inst_rx_parallel_data(418) & COLD_DATA_RxTx_inst_rx_parallel_data(417) & COLD_DATA_RxTx_inst_rx_parallel_data(416) & COLD_DATA_RxTx_inst_rx_parallel_data(415) & COLD_DATA_RxTx_inst_rx_parallel_data(414) & COLD_DATA_RxTx_inst_rx_parallel_data(413) & COLD_DATA_RxTx_inst_rx_parallel_data(412) & COLD_DATA_RxTx_inst_rx_parallel_data(411) & COLD_DATA_RxTx_inst_rx_parallel_data(410) & COLD_DATA_RxTx_inst_rx_parallel_data(409) & COLD_DATA_RxTx_inst_rx_parallel_data(408) & COLD_DATA_RxTx_inst_rx_parallel_data(407) & COLD_DATA_RxTx_inst_rx_parallel_data(406) & COLD_DATA_RxTx_inst_rx_parallel_data(405) & COLD_DATA_RxTx_inst_rx_parallel_data(404) & COLD_DATA_RxTx_inst_rx_parallel_data(403) & COLD_DATA_RxTx_inst_rx_parallel_data(402) & COLD_DATA_RxTx_inst_rx_parallel_data(401) & COLD_DATA_RxTx_inst_rx_parallel_data(400) & COLD_DATA_RxTx_inst_rx_parallel_data(398) & COLD_DATA_RxTx_inst_rx_parallel_data(397) & COLD_DATA_RxTx_inst_rx_parallel_data(383) & COLD_DATA_RxTx_inst_rx_parallel_data(382) & COLD_DATA_RxTx_inst_rx_parallel_data(381) & COLD_DATA_RxTx_inst_rx_parallel_data(380) & COLD_DATA_RxTx_inst_rx_parallel_data(379) & COLD_DATA_RxTx_inst_rx_parallel_data(378) & COLD_DATA_RxTx_inst_rx_parallel_data(377) & COLD_DATA_RxTx_inst_rx_parallel_data(376) & COLD_DATA_RxTx_inst_rx_parallel_data(375) & COLD_DATA_RxTx_inst_rx_parallel_data(374) & COLD_DATA_RxTx_inst_rx_parallel_data(373) & COLD_DATA_RxTx_inst_rx_parallel_data(372) & COLD_DATA_RxTx_inst_rx_parallel_data(371) & COLD_DATA_RxTx_inst_rx_parallel_data(370) & COLD_DATA_RxTx_inst_rx_parallel_data(369) & COLD_DATA_RxTx_inst_rx_parallel_data(368) & COLD_DATA_RxTx_inst_rx_parallel_data(367) & COLD_DATA_RxTx_inst_rx_parallel_data(366) & COLD_DATA_RxTx_inst_rx_parallel_data(365) & COLD_DATA_RxTx_inst_rx_parallel_data(364) & COLD_DATA_RxTx_inst_rx_parallel_data(363) & COLD_DATA_RxTx_inst_rx_parallel_data(362) & COLD_DATA_RxTx_inst_rx_parallel_data(361) & COLD_DATA_RxTx_inst_rx_parallel_data(360) & COLD_DATA_RxTx_inst_rx_parallel_data(359) & COLD_DATA_RxTx_inst_rx_parallel_data(358) & COLD_DATA_RxTx_inst_rx_parallel_data(357) & COLD_DATA_RxTx_inst_rx_parallel_data(356) & COLD_DATA_RxTx_inst_rx_parallel_data(355) & COLD_DATA_RxTx_inst_rx_parallel_data(354) & COLD_DATA_RxTx_inst_rx_parallel_data(353) & COLD_DATA_RxTx_inst_rx_parallel_data(352) & COLD_DATA_RxTx_inst_rx_parallel_data(351) & COLD_DATA_RxTx_inst_rx_parallel_data(350) & COLD_DATA_RxTx_inst_rx_parallel_data(349) & COLD_DATA_RxTx_inst_rx_parallel_data(348) & COLD_DATA_RxTx_inst_rx_parallel_data(347) & COLD_DATA_RxTx_inst_rx_parallel_data(346) & COLD_DATA_RxTx_inst_rx_parallel_data(345) & COLD_DATA_RxTx_inst_rx_parallel_data(344) & COLD_DATA_RxTx_inst_rx_parallel_data(343) & COLD_DATA_RxTx_inst_rx_parallel_data(342) & COLD_DATA_RxTx_inst_rx_parallel_data(341) & COLD_DATA_RxTx_inst_rx_parallel_data(340) & COLD_DATA_RxTx_inst_rx_parallel_data(339) & COLD_DATA_RxTx_inst_rx_parallel_data(338) & COLD_DATA_RxTx_inst_rx_parallel_data(337) & COLD_DATA_RxTx_inst_rx_parallel_data(336) & COLD_DATA_RxTx_inst_rx_parallel_data(334) & COLD_DATA_RxTx_inst_rx_parallel_data(333) & COLD_DATA_RxTx_inst_rx_parallel_data(319) & COLD_DATA_RxTx_inst_rx_parallel_data(318) & COLD_DATA_RxTx_inst_rx_parallel_data(317) & COLD_DATA_RxTx_inst_rx_parallel_data(316) & COLD_DATA_RxTx_inst_rx_parallel_data(315) & COLD_DATA_RxTx_inst_rx_parallel_data(314) & COLD_DATA_RxTx_inst_rx_parallel_data(313) & COLD_DATA_RxTx_inst_rx_parallel_data(312) & COLD_DATA_RxTx_inst_rx_parallel_data(311) & COLD_DATA_RxTx_inst_rx_parallel_data(310) & COLD_DATA_RxTx_inst_rx_parallel_data(309) & COLD_DATA_RxTx_inst_rx_parallel_data(308) & COLD_DATA_RxTx_inst_rx_parallel_data(307) & COLD_DATA_RxTx_inst_rx_parallel_data(306) & COLD_DATA_RxTx_inst_rx_parallel_data(305) & COLD_DATA_RxTx_inst_rx_parallel_data(304) & COLD_DATA_RxTx_inst_rx_parallel_data(303) & COLD_DATA_RxTx_inst_rx_parallel_data(302) & COLD_DATA_RxTx_inst_rx_parallel_data(301) & COLD_DATA_RxTx_inst_rx_parallel_data(300) & COLD_DATA_RxTx_inst_rx_parallel_data(299) & COLD_DATA_RxTx_inst_rx_parallel_data(298) & COLD_DATA_RxTx_inst_rx_parallel_data(297) & COLD_DATA_RxTx_inst_rx_parallel_data(296) & COLD_DATA_RxTx_inst_rx_parallel_data(295) & COLD_DATA_RxTx_inst_rx_parallel_data(294) & COLD_DATA_RxTx_inst_rx_parallel_data(293) & COLD_DATA_RxTx_inst_rx_parallel_data(292) & COLD_DATA_RxTx_inst_rx_parallel_data(291) & COLD_DATA_RxTx_inst_rx_parallel_data(290) & COLD_DATA_RxTx_inst_rx_parallel_data(289) & COLD_DATA_RxTx_inst_rx_parallel_data(288) & COLD_DATA_RxTx_inst_rx_parallel_data(287) & COLD_DATA_RxTx_inst_rx_parallel_data(286) & COLD_DATA_RxTx_inst_rx_parallel_data(285) & COLD_DATA_RxTx_inst_rx_parallel_data(284) & COLD_DATA_RxTx_inst_rx_parallel_data(283) & COLD_DATA_RxTx_inst_rx_parallel_data(282) & COLD_DATA_RxTx_inst_rx_parallel_data(281) & COLD_DATA_RxTx_inst_rx_parallel_data(280) & COLD_DATA_RxTx_inst_rx_parallel_data(279) & COLD_DATA_RxTx_inst_rx_parallel_data(278) & COLD_DATA_RxTx_inst_rx_parallel_data(277) & COLD_DATA_RxTx_inst_rx_parallel_data(276) & COLD_DATA_RxTx_inst_rx_parallel_data(275) & COLD_DATA_RxTx_inst_rx_parallel_data(274) & COLD_DATA_RxTx_inst_rx_parallel_data(273) & COLD_DATA_RxTx_inst_rx_parallel_data(272) & COLD_DATA_RxTx_inst_rx_parallel_data(270) & COLD_DATA_RxTx_inst_rx_parallel_data(269) & COLD_DATA_RxTx_inst_rx_parallel_data(255) & COLD_DATA_RxTx_inst_rx_parallel_data(254) & COLD_DATA_RxTx_inst_rx_parallel_data(253) & COLD_DATA_RxTx_inst_rx_parallel_data(252) & COLD_DATA_RxTx_inst_rx_parallel_data(251) & COLD_DATA_RxTx_inst_rx_parallel_data(250) & COLD_DATA_RxTx_inst_rx_parallel_data(249) & COLD_DATA_RxTx_inst_rx_parallel_data(248) & COLD_DATA_RxTx_inst_rx_parallel_data(247) & COLD_DATA_RxTx_inst_rx_parallel_data(246) & COLD_DATA_RxTx_inst_rx_parallel_data(245) & COLD_DATA_RxTx_inst_rx_parallel_data(244) & COLD_DATA_RxTx_inst_rx_parallel_data(243) & COLD_DATA_RxTx_inst_rx_parallel_data(242) & COLD_DATA_RxTx_inst_rx_parallel_data(241) & COLD_DATA_RxTx_inst_rx_parallel_data(240) & COLD_DATA_RxTx_inst_rx_parallel_data(239) & COLD_DATA_RxTx_inst_rx_parallel_data(238) & COLD_DATA_RxTx_inst_rx_parallel_data(237) & COLD_DATA_RxTx_inst_rx_parallel_data(236) & COLD_DATA_RxTx_inst_rx_parallel_data(235) & COLD_DATA_RxTx_inst_rx_parallel_data(234) & COLD_DATA_RxTx_inst_rx_parallel_data(233) & COLD_DATA_RxTx_inst_rx_parallel_data(232) & COLD_DATA_RxTx_inst_rx_parallel_data(231) & COLD_DATA_RxTx_inst_rx_parallel_data(230) & COLD_DATA_RxTx_inst_rx_parallel_data(229) & COLD_DATA_RxTx_inst_rx_parallel_data(228) & COLD_DATA_RxTx_inst_rx_parallel_data(227) & COLD_DATA_RxTx_inst_rx_parallel_data(226) & COLD_DATA_RxTx_inst_rx_parallel_data(225) & COLD_DATA_RxTx_inst_rx_parallel_data(224) & COLD_DATA_RxTx_inst_rx_parallel_data(223) & COLD_DATA_RxTx_inst_rx_parallel_data(222) & COLD_DATA_RxTx_inst_rx_parallel_data(221) & COLD_DATA_RxTx_inst_rx_parallel_data(220) & COLD_DATA_RxTx_inst_rx_parallel_data(219) & COLD_DATA_RxTx_inst_rx_parallel_data(218) & COLD_DATA_RxTx_inst_rx_parallel_data(217) & COLD_DATA_RxTx_inst_rx_parallel_data(216) & COLD_DATA_RxTx_inst_rx_parallel_data(215) & COLD_DATA_RxTx_inst_rx_parallel_data(214) & COLD_DATA_RxTx_inst_rx_parallel_data(213) & COLD_DATA_RxTx_inst_rx_parallel_data(212) & COLD_DATA_RxTx_inst_rx_parallel_data(211) & COLD_DATA_RxTx_inst_rx_parallel_data(210) & COLD_DATA_RxTx_inst_rx_parallel_data(209) & COLD_DATA_RxTx_inst_rx_parallel_data(208) & COLD_DATA_RxTx_inst_rx_parallel_data(206) & COLD_DATA_RxTx_inst_rx_parallel_data(205) & COLD_DATA_RxTx_inst_rx_parallel_data(191) & COLD_DATA_RxTx_inst_rx_parallel_data(190) & COLD_DATA_RxTx_inst_rx_parallel_data(189) & COLD_DATA_RxTx_inst_rx_parallel_data(188) & COLD_DATA_RxTx_inst_rx_parallel_data(187) & COLD_DATA_RxTx_inst_rx_parallel_data(186) & COLD_DATA_RxTx_inst_rx_parallel_data(185) & COLD_DATA_RxTx_inst_rx_parallel_data(184) & COLD_DATA_RxTx_inst_rx_parallel_data(183) & COLD_DATA_RxTx_inst_rx_parallel_data(182) & COLD_DATA_RxTx_inst_rx_parallel_data(181) & COLD_DATA_RxTx_inst_rx_parallel_data(180) & COLD_DATA_RxTx_inst_rx_parallel_data(179) & COLD_DATA_RxTx_inst_rx_parallel_data(178) & COLD_DATA_RxTx_inst_rx_parallel_data(177) & COLD_DATA_RxTx_inst_rx_parallel_data(176) & COLD_DATA_RxTx_inst_rx_parallel_data(175) & COLD_DATA_RxTx_inst_rx_parallel_data(174) & COLD_DATA_RxTx_inst_rx_parallel_data(173) & COLD_DATA_RxTx_inst_rx_parallel_data(172) & COLD_DATA_RxTx_inst_rx_parallel_data(171) & COLD_DATA_RxTx_inst_rx_parallel_data(170) & COLD_DATA_RxTx_inst_rx_parallel_data(169) & COLD_DATA_RxTx_inst_rx_parallel_data(168) & COLD_DATA_RxTx_inst_rx_parallel_data(167) & COLD_DATA_RxTx_inst_rx_parallel_data(166) & COLD_DATA_RxTx_inst_rx_parallel_data(165) & COLD_DATA_RxTx_inst_rx_parallel_data(164) & COLD_DATA_RxTx_inst_rx_parallel_data(163) & COLD_DATA_RxTx_inst_rx_parallel_data(162) & COLD_DATA_RxTx_inst_rx_parallel_data(161) & COLD_DATA_RxTx_inst_rx_parallel_data(160) & COLD_DATA_RxTx_inst_rx_parallel_data(159) & COLD_DATA_RxTx_inst_rx_parallel_data(158) & COLD_DATA_RxTx_inst_rx_parallel_data(157) & COLD_DATA_RxTx_inst_rx_parallel_data(156) & COLD_DATA_RxTx_inst_rx_parallel_data(155) & COLD_DATA_RxTx_inst_rx_parallel_data(154) & COLD_DATA_RxTx_inst_rx_parallel_data(153) & COLD_DATA_RxTx_inst_rx_parallel_data(152) & COLD_DATA_RxTx_inst_rx_parallel_data(151) & COLD_DATA_RxTx_inst_rx_parallel_data(150) & COLD_DATA_RxTx_inst_rx_parallel_data(149) & COLD_DATA_RxTx_inst_rx_parallel_data(148) & COLD_DATA_RxTx_inst_rx_parallel_data(147) & COLD_DATA_RxTx_inst_rx_parallel_data(146) & COLD_DATA_RxTx_inst_rx_parallel_data(145) & COLD_DATA_RxTx_inst_rx_parallel_data(144) & COLD_DATA_RxTx_inst_rx_parallel_data(142) & COLD_DATA_RxTx_inst_rx_parallel_data(141) & COLD_DATA_RxTx_inst_rx_parallel_data(127) & COLD_DATA_RxTx_inst_rx_parallel_data(126) & COLD_DATA_RxTx_inst_rx_parallel_data(125) & COLD_DATA_RxTx_inst_rx_parallel_data(124) & COLD_DATA_RxTx_inst_rx_parallel_data(123) & COLD_DATA_RxTx_inst_rx_parallel_data(122) & COLD_DATA_RxTx_inst_rx_parallel_data(121) & COLD_DATA_RxTx_inst_rx_parallel_data(120) & COLD_DATA_RxTx_inst_rx_parallel_data(119) & COLD_DATA_RxTx_inst_rx_parallel_data(118) & COLD_DATA_RxTx_inst_rx_parallel_data(117) & COLD_DATA_RxTx_inst_rx_parallel_data(116) & COLD_DATA_RxTx_inst_rx_parallel_data(115) & COLD_DATA_RxTx_inst_rx_parallel_data(114) & COLD_DATA_RxTx_inst_rx_parallel_data(113) & COLD_DATA_RxTx_inst_rx_parallel_data(112) & COLD_DATA_RxTx_inst_rx_parallel_data(111) & COLD_DATA_RxTx_inst_rx_parallel_data(110) & COLD_DATA_RxTx_inst_rx_parallel_data(109) & COLD_DATA_RxTx_inst_rx_parallel_data(108) & COLD_DATA_RxTx_inst_rx_parallel_data(107) & COLD_DATA_RxTx_inst_rx_parallel_data(106) & COLD_DATA_RxTx_inst_rx_parallel_data(105) & COLD_DATA_RxTx_inst_rx_parallel_data(104) & COLD_DATA_RxTx_inst_rx_parallel_data(103) & COLD_DATA_RxTx_inst_rx_parallel_data(102) & COLD_DATA_RxTx_inst_rx_parallel_data(101) & COLD_DATA_RxTx_inst_rx_parallel_data(100) & COLD_DATA_RxTx_inst_rx_parallel_data(99) & COLD_DATA_RxTx_inst_rx_parallel_data(98) & COLD_DATA_RxTx_inst_rx_parallel_data(97) & COLD_DATA_RxTx_inst_rx_parallel_data(96) & COLD_DATA_RxTx_inst_rx_parallel_data(95) & COLD_DATA_RxTx_inst_rx_parallel_data(94) & COLD_DATA_RxTx_inst_rx_parallel_data(93) & COLD_DATA_RxTx_inst_rx_parallel_data(92) & COLD_DATA_RxTx_inst_rx_parallel_data(91) & COLD_DATA_RxTx_inst_rx_parallel_data(90) & COLD_DATA_RxTx_inst_rx_parallel_data(89) & COLD_DATA_RxTx_inst_rx_parallel_data(88) & COLD_DATA_RxTx_inst_rx_parallel_data(87) & COLD_DATA_RxTx_inst_rx_parallel_data(86) & COLD_DATA_RxTx_inst_rx_parallel_data(85) & COLD_DATA_RxTx_inst_rx_parallel_data(84) & COLD_DATA_RxTx_inst_rx_parallel_data(83) & COLD_DATA_RxTx_inst_rx_parallel_data(82) & COLD_DATA_RxTx_inst_rx_parallel_data(81) & COLD_DATA_RxTx_inst_rx_parallel_data(80) & COLD_DATA_RxTx_inst_rx_parallel_data(78) & COLD_DATA_RxTx_inst_rx_parallel_data(77) & COLD_DATA_RxTx_inst_rx_parallel_data(63) & COLD_DATA_RxTx_inst_rx_parallel_data(62) & COLD_DATA_RxTx_inst_rx_parallel_data(61) & COLD_DATA_RxTx_inst_rx_parallel_data(60) & COLD_DATA_RxTx_inst_rx_parallel_data(59) & COLD_DATA_RxTx_inst_rx_parallel_data(58) & COLD_DATA_RxTx_inst_rx_parallel_data(57) & COLD_DATA_RxTx_inst_rx_parallel_data(56) & COLD_DATA_RxTx_inst_rx_parallel_data(55) & COLD_DATA_RxTx_inst_rx_parallel_data(54) & COLD_DATA_RxTx_inst_rx_parallel_data(53) & COLD_DATA_RxTx_inst_rx_parallel_data(52) & COLD_DATA_RxTx_inst_rx_parallel_data(51) & COLD_DATA_RxTx_inst_rx_parallel_data(50) & COLD_DATA_RxTx_inst_rx_parallel_data(49) & COLD_DATA_RxTx_inst_rx_parallel_data(48) & COLD_DATA_RxTx_inst_rx_parallel_data(47) & COLD_DATA_RxTx_inst_rx_parallel_data(46) & COLD_DATA_RxTx_inst_rx_parallel_data(45) & COLD_DATA_RxTx_inst_rx_parallel_data(44) & COLD_DATA_RxTx_inst_rx_parallel_data(43) & COLD_DATA_RxTx_inst_rx_parallel_data(42) & COLD_DATA_RxTx_inst_rx_parallel_data(41) & COLD_DATA_RxTx_inst_rx_parallel_data(40) & COLD_DATA_RxTx_inst_rx_parallel_data(39) & COLD_DATA_RxTx_inst_rx_parallel_data(38) & COLD_DATA_RxTx_inst_rx_parallel_data(37) & COLD_DATA_RxTx_inst_rx_parallel_data(36) & COLD_DATA_RxTx_inst_rx_parallel_data(35) & COLD_DATA_RxTx_inst_rx_parallel_data(34) & COLD_DATA_RxTx_inst_rx_parallel_data(33) & COLD_DATA_RxTx_inst_rx_parallel_data(32) & COLD_DATA_RxTx_inst_rx_parallel_data(31) & COLD_DATA_RxTx_inst_rx_parallel_data(30) & COLD_DATA_RxTx_inst_rx_parallel_data(29) & COLD_DATA_RxTx_inst_rx_parallel_data(28) & COLD_DATA_RxTx_inst_rx_parallel_data(27) & COLD_DATA_RxTx_inst_rx_parallel_data(26) & COLD_DATA_RxTx_inst_rx_parallel_data(25) & COLD_DATA_RxTx_inst_rx_parallel_data(24) & COLD_DATA_RxTx_inst_rx_parallel_data(23) & COLD_DATA_RxTx_inst_rx_parallel_data(22) & COLD_DATA_RxTx_inst_rx_parallel_data(21) & COLD_DATA_RxTx_inst_rx_parallel_data(20) & COLD_DATA_RxTx_inst_rx_parallel_data(19) & COLD_DATA_RxTx_inst_rx_parallel_data(18) & COLD_DATA_RxTx_inst_rx_parallel_data(17) & COLD_DATA_RxTx_inst_rx_parallel_data(16) & COLD_DATA_RxTx_inst_rx_parallel_data(14) & COLD_DATA_RxTx_inst_rx_parallel_data(13);

	rx_runningdisp <= COLD_DATA_RxTx_inst_rx_parallel_data(463) & COLD_DATA_RxTx_inst_rx_parallel_data(399) & COLD_DATA_RxTx_inst_rx_parallel_data(335) & COLD_DATA_RxTx_inst_rx_parallel_data(271) & COLD_DATA_RxTx_inst_rx_parallel_data(207) & COLD_DATA_RxTx_inst_rx_parallel_data(143) & COLD_DATA_RxTx_inst_rx_parallel_data(79) & COLD_DATA_RxTx_inst_rx_parallel_data(15);

	rx_patterndetect <= COLD_DATA_RxTx_inst_rx_parallel_data(460) & COLD_DATA_RxTx_inst_rx_parallel_data(396) & COLD_DATA_RxTx_inst_rx_parallel_data(332) & COLD_DATA_RxTx_inst_rx_parallel_data(268) & COLD_DATA_RxTx_inst_rx_parallel_data(204) & COLD_DATA_RxTx_inst_rx_parallel_data(140) & COLD_DATA_RxTx_inst_rx_parallel_data(76) & COLD_DATA_RxTx_inst_rx_parallel_data(12);

	rx_syncstatus <= COLD_DATA_RxTx_inst_rx_parallel_data(458) & COLD_DATA_RxTx_inst_rx_parallel_data(394) & COLD_DATA_RxTx_inst_rx_parallel_data(330) & COLD_DATA_RxTx_inst_rx_parallel_data(266) & COLD_DATA_RxTx_inst_rx_parallel_data(202) & COLD_DATA_RxTx_inst_rx_parallel_data(138) & COLD_DATA_RxTx_inst_rx_parallel_data(74) & COLD_DATA_RxTx_inst_rx_parallel_data(10);

end architecture rtl; -- of COLD_DATA_RxTx
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_xcvr_native_av" version="16.0" >
-- Retrieval info: 	<generic name="device_family" value="Arria V" />
-- Retrieval info: 	<generic name="show_advanced_features" value="0" />
-- Retrieval info: 	<generic name="device_speedgrade" value="fastest" />
-- Retrieval info: 	<generic name="message_level" value="error" />
-- Retrieval info: 	<generic name="tx_enable" value="0" />
-- Retrieval info: 	<generic name="rx_enable" value="1" />
-- Retrieval info: 	<generic name="enable_std" value="1" />
-- Retrieval info: 	<generic name="set_data_path_select" value="standard" />
-- Retrieval info: 	<generic name="channels" value="8" />
-- Retrieval info: 	<generic name="bonded_mode" value="non_bonded" />
-- Retrieval info: 	<generic name="enable_simple_interface" value="1" />
-- Retrieval info: 	<generic name="set_data_rate" value="1280" />
-- Retrieval info: 	<generic name="pma_direct_width" value="80" />
-- Retrieval info: 	<generic name="tx_pma_clk_div" value="1" />
-- Retrieval info: 	<generic name="pll_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="pll_external_enable" value="1" />
-- Retrieval info: 	<generic name="plls" value="1" />
-- Retrieval info: 	<generic name="pll_select" value="0" />
-- Retrieval info: 	<generic name="pll_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="cdr_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_refclk_select" value="0" />
-- Retrieval info: 	<generic name="set_cdr_refclk_freq" value="128.0 MHz" />
-- Retrieval info: 	<generic name="rx_ppm_detect_threshold" value="1000" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_clkout" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtodata" value="1" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtoref" value="1" />
-- Retrieval info: 	<generic name="enable_ports_rx_manual_cdr_mode" value="0" />
-- Retrieval info: 	<generic name="rx_clkslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_seriallpbken" value="0" />
-- Retrieval info: 	<generic name="std_protocol_hint" value="basic" />
-- Retrieval info: 	<generic name="std_pcs_pma_width" value="10" />
-- Retrieval info: 	<generic name="std_low_latency_bypass_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_pcfifo_mode" value="register_fifo" />
-- Retrieval info: 	<generic name="std_rx_pcfifo_mode" value="register_fifo" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_mode" value="manual" />
-- Retrieval info: 	<generic name="std_rx_byte_order_symbol_count" value="1" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pattern" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pad" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_flag" value="0" />
-- Retrieval info: 	<generic name="std_tx_byte_ser_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_deser_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_8b10b_enable" value="1" />
-- Retrieval info: 	<generic name="std_tx_8b10b_disp_ctrl_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_8b10b_enable" value="1" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_p" value="00000" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_n" value="00000" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_mode" value="sync_sm" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern_len" value="10" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern" value="27C" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rknumber" value="5" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_renumber" value="5" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rgnumber" value="5" />
-- Retrieval info: 	<generic name="std_rx_run_length_val" value="10" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_patternalign" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_a1a2size" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_runlength_err" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitrev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byterev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_polinv" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_polinv" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_elecidle" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_prbs_status" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="125 Mhz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_clk_network" value="xN" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_clk_network" value="xN" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_clk_network" value="xN" />
-- Retrieval info: </instance>
-- IPFS_FILES : COLD_DATA_RxTx.vho
-- RELATED_FILES: COLD_DATA_RxTx.vhd, altera_xcvr_functions.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_native_av_functions_h.sv, altera_xcvr_native_av.sv, altera_xcvr_data_adapter_av.sv
