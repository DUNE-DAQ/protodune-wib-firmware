// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:51 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZIPLgkArVotGSohqEkUR+64TVQFde4jSlsBay/qMP6KT7OHoB7HyDxtY2i2j/BsD
T825dwKB2jpTOwk0HjlG8W8X+W/3MQFbxvti3wf3zTomA4wM2TSTThyXkmdqKIfx
3bLf/yfHZFlY9q9Xbu/YU1YrBFEiyGBfsXB60ZBw9PI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21968)
A7HiJzHwdRgXZz+71kV7lfHyWY7lWyGicAUfFmA388kNwUEmzTU6QL/6mTtJUPFD
ygKNVU8SA4CrbCauyGfQUo2YpAooOON2vN1b51eMzLfhK4zBHFCxIxr0D8rNF4Me
cr8C+H5RZVynvajIiJA+bt8pVPb5pHHduIx8DhDaDKPmH+DoF+twSe3KipWYM/vF
aFgaweVkrVC8qf7ypcmimMxRjvkTSz9Ut1ngtUxcyEFN6jEngqTAjmRHFd9P8Ov1
88ug4+bAldXzggoh21Satyg/9PJ/V5C5w8CEUbZVVn61XfqYR+xBuoIupQI8/gsY
WMl5Z35w8IcCLJwwp4ZUZD3NC5Nt3MRUJo9lX8z74VGAQ0oqobWVeqHYNMFPAmLZ
Pa/SJbRLN8yqY7eLlO5K6wru0K2vkpj6G1W+dZBr323S4M5U1Ia3oKrzMW+HeQj2
TvaPn1aRZCTVtBIU8f6tFk96TlOSgnlATQe0YMltC9i4NMAYhdEYc4fakCV+V8Sb
u5TjGc1nJbRZdUO4uNJNsj+ivCHAUVLRpliK9RW1NiTuRQkcrYUdJVgaMipSVj/q
WQzP4P9mMGrE5SgpEOo0gKGoXO2o5paO146Ktwd1aBCAaPHUloorMygV9kCOPG5x
tinMiQ7f488FLtVY9vhVI9s+02G7kyRA5NmRJJC1t/y0TFLv/KlCcJWzCdR9xLMu
974v7OX1Y2ebXMu0vP2rvrxyPMSC/7eSzFf7GAjjwaDUQGIwMSzLBanik1gVfucH
DC74W8JS1u1II4GGGMHLAMU8Qhs02OEFFMsaqgk935mACWhdZsbSV9cVGWfX2/K9
lPwKxRYXGNGFsFZbNZdvuctxk3jGgPX91WJ1atlJt+0YAvn7Xd6sz+SnJn+khzNo
l+4767GBKT69x5Lv15mWuYLAfD+87GzxELHGkJrikR5UAFyFwsIK2tO8VON2Atzg
NtizN9VkiIohER7Msb/zOhQ5hEDEFhGhDxpw/n7WWleDWYmDnEUZiDLfI7cLuGiJ
xqSgjZJWDSwH211ZHy29eQNafEwWhZKfWOE72u7VSojQHc62wo4Er1ZxBubsQSPX
bA62LrksbiLnMof91L294zmvxaWpiWDH4m6tPaniG50ugYrWIM/SktdCEYG3u3Qj
FHBEtnZWODik3BOLEmtEL1S//9nlqusGRmjv2EtrXBJpkroWqoMubCRer9Hjmzl0
CBKz2GrEC1JOxV9NcfBnvOXdbsq6rW8d+IlAe7/zR/XqauIpaOnwhWZW4jG7Z9+4
SIvpajRjNGhmBpP3d/D+/oEfKqT9yvLVV+KEZar/MI8QWnSwFCyahIy2k5FU4thr
NGWemvx2U5dQ4RC9HTItZT6KhitRtllApWIxwPRBAc+R9ZT5tO/OBy7PHqsi1XFJ
m/6F4yskkvYhp2C9gC1ys4cjxVCgHwRjUMccQ01ppgAbu3BCM0N6rf53GnRhJmI6
us354PEKpI48NwWZv2MhRvFdKLtELXsf3jls/w9M8zVSTOZMg0X4zRqXQBe5dbYo
Y/ks4w+nGauo3aCcZizu3BaxwcUhgOfVM+dkN2S3l64YYWTW9avNF0Uo4GW0WvR5
1nJZSuMAvJEvuHuHngFPq7y2L5zM32lduCH7X+7OKk/9AtGBYuM/Q8NbFgpfgxEU
TMlVQt/2SxEnp2mwbalnommwtsjVeeTU41KB3iwOY7RxmTck8937atBZj60evit7
twFRNjCFQ/C1pwOia+l+GmFBZNTwcZkcnjn8A1NjeqsjngFozNgiaogmNy0d16lK
mqeS5ztjp8XqQVfrnvskMw3GhEkZX1M8oVWfWZ3QZtHZPDumJvfHK47XBUY5fxqk
W76FA2/ZtgeL+RI3s7TBO25G6B1FrBHIOodmI9aJfgQ7ZzzjBpVIoYgl4LsI2U1l
XiApfCbJSasadndAaxa/OmR8FHpmivxP0MAimAYA5EFpOywpblqDVRqCSgif4XdD
xy1UzEFo3UcFOuKo8uie6EOpBVxTBRKKIOtYS0zLW/pwZMXyjo81vri/BYE2utS6
8DHdZkL6k0eQ2AWYbvGALZTjlbNrVIuRygiowX29cM6kLgFuX6LeTp3XpQNI32u0
gIa/JTYB53YPW1rVP1+WaQjthk4cX8qCxqUod6wS5g+puLOjRrsH1fgG92Gmhui9
9YBJDPyiHfMzsBvIlrSoDcS0b9JfhKC5jXaV+WyGa7vF69A4EHW0jDt+yxWMAEan
hwF+VJsYluyg/9zY2mDm/yKlZyncPe3WwEmmlmcrRLPWEtU29AK/mVeiCQL9ylqv
YmYTA36DWwUCdjwtOGOeKBJ/QquGeC/A7tMm3BzzTzM/+G+xKhm5i5iv/UcQO2KP
A0bZmO1HaAhiJxZqI2lsxqHLAIZ4ZAj5gn+JAnGtxgb+aQifetD1o30Zxc542+WV
ncwF/9VNyWifYbsmb6S1I2H2oYLXVvFle9D6goGkkCHT6qhTJRbnqFsfYmRz90t2
fryPZPKngDsSCT7fKZyLEjEazpNLCL0WTbH5p/68oPYP1z8LCzHvBA68vzlMionf
Qu9A0pbIXHDA1wYg9QQOznREQxWAKYd8qM+pK6lmrQtsYbsikvvCHvFJeeum7fmv
rU2sJppRb8biykaVUDPh/3Hy/fHXMnb+kwmquoxb5YJ2gIk68iKm4ic95Lh/vTBw
GtJ9JLOF7tXGI7V8/aREFgBiVJHXo3HbteDvLjXDmivYLaeyV0Cm6htYyhrLsm/6
Cva+w9gdjEfNX44WM9//YHPw374yGjEeMwyYoPISNUfBkwync7aPmxnyKKrZuhvP
NLzj5Ph2ezkOzEUSRSLdmIvXOeyub7+xxrNxQ8D9Ae6SeIPzWRKzZeR5wmEo3me/
IQvqcpJgyAlnr2a1fF5sFP5VkDw3UXEDZKBLy+xwnIba9R5cil2Kl83tWbbArPKh
3YJPxRhqHI88/aNiz+aOrhuck9l+8t3ev+xAmmuWUxlywp0UsvYsHxBTLC4VVtsU
18/bSq7Yg5nhigAs8vvOp7vvMuNWqx2t/16X8Jv0iS+9ye8pYsYWwlYCWKWeIZVg
Tx2lkoqcwA5l/SQFnB+hTOdEKMm0lnLKfIOeGRIlT45eTtoCeCOMr6Z09PnItjgA
tSH3UUQQlIuER2I/yLy0cjOUuoMWMUYHWel31k0ZIcYqGo5eWKAniDWIdVk3cEJT
baXETeKD/qml6pShuBiBHtdOf5XT5TQYHhs2Q6L66V4VqH5fccriQz+cIqhzjVGL
nfPMfcZf/zrijP9tCJ3zbA94GJufG+okVgENQAH0ivezhS3NkbH7A9jcnVvlhvnH
hdJtSKipJWD9k/GfLHNAA9/zNleqNwxsH+plhY4U8mnv0ohSMd2R5sFDKLtCiiDc
p/am0TOROrjJm5ZgkYssynKMrz8zV17AuHqPrrlay6g5NjrvmBaBrCwGf+ur5KKU
llwNkdaMPOl3eab9mTiEd9p641KPISvKoa4Sq+paqm3T6jcsfIIUEVRlVHClkPYw
MxKmu02CCUSKLV+2eERVdthgZ2blGTHzFlH9g81KGqubrE/6GktBLWX2DAWKLdJT
AW2UYsVDM7zScr/rZSFuPAMf6/EBScgCDm/GK63B1aNDV/EH3F0F6tinszllRZ80
wn27m2OnTKG5houMkeqvx7btsR4CE9T29Po+yeJNEQuJ7uGvaz3h63vCJao9sCGB
yYN/0k1oOl6c5BpHVKkx7mi8cNPveH2vr4li13FLSL+me/clDJqSg5o0Le3iqZ+U
MB9/vnjA2gMxBkm/6b3C5vjZOVWlWbdwjHR2rNBI3LkQDpFsAuyJSa0nT8UePW5q
OHr/BnIFT8+ShY04xFYFqDN6B8MfVl0l1qhFrvnjBU49iCgMeTZYH/1guD6Jzv97
GEDPiY1gw2XtsMg1CLIAedpOPNfISlqxXJUKx8rNlxxv3QLg/tvXhISwYv9pQugM
FXx0+IVOBBBc1f/MnsXtkGIKsrYyjUzJQggKD0XmsdjOi/4ytuGuVVHeO8jYK2Sd
qxLXtSlNjmHPgC+J85b+EZ9yyxbOIw9f2N5rf0It/74xhaQuhUG5m147p+o+uXcQ
VKs+mTRoMRSRJUTfD2d+R/ONdQ9E/6qIHJx7+XxLqiczcSFISeVILL7YD4ntuLwD
tH3rtE/l49pN8rr6hwLFFsf7IRMBGIejYaUmogSWqzRbUE/xHesGy96Xj7q2RN29
0rhlPBDOvR1DuaJjd3glywPVonNQCQHhwxZt6sKjof18S2es6sM6G2v4Ntoc1Sh4
/gIOjLXVs1bdjzc6Q4PVMlSZgXB3tQ0RwSJGVS/HLyK1Pt7bkx3NyV2M4bPwS3Jj
ea7QH0nAoUEV5H7bORMZFwqarAGy10bYymJQkLSRwGBQfh7SqdSziYBsLq/IMcqD
bwIU/Bk4yFpykOac0yjV1uymmsH1JcYz5mPbd2i3AyK2P7R76XRcpKlgP6wCCz3E
sDzdzeRSPLLkwcj+I+b+xxkk7/J/JF54gbK9xqYj1MYq5U4WtGRe6TeYlJyWyJ7U
KMLkFT1YYCwWLzoD9iolThvBh14xIkYjJRTNWUfptfvG0fz/GLSAzO8oHpFdZB43
Ay+U9PBkvSDDkeizABac8rW6jyQ74uaaelgmoLxpowtwqXE6IsCKtM5L225+D07s
8vUew6qo+CbR0Jh6aa1sDHxfWn9E0ZDKg2XDlCJpiCmpBiU0A/vz3FgAIp1RdoGZ
QmvqlXNSuYepD2aSDY0F1guXE8kJ0COOd8wVc+lRNM0YdIAJ2QAELPYmRmKp8PN2
eXRfy7I80ZMZCxXaPNEdH/RzJD4NfsMiirCUEeOO5Mjz+Rabp8Cjcr7Yq11j9aox
IC+v29VLUlyQMg3dZXBU2R7auVQLaiKnO7NM3zJRPYURfR5k6IvOyF/5g6uR2Kg/
y+RCNCZNAIbidkaCdgCdb2WxUZBp3RVhIskxyQ9UsQYYDse/jN2FgNKObZfC6+jM
GzLgMvHT1dahuWa7jrMzdtgdyjeNmBXAsJDMPSouSfMWWxYWlqZFERjqnHRPVk7O
kBueZGVSF9EjaLMlqGRsmBzUwvskCw2hfTwH4uuipTtwKfohen2ctUG3I8FUPmjh
dhcb3z68/r50noVH9Rtr27LRAwwN4ZYdFoIeyfJ9d+Nj9LpEaZxI3k9OwWADRiu/
+eg9TIr2QV9Jk2/S/G9Fgl9yB3XzCq9vTzq/ou7nJByXtt7mzUdoKLebbRaczUWq
xQv3ccfoasH7FOALJhJ0KZouGOAkjkpboO8fqzCyNp7HpW7vSzH4p9eDY/DcVHdh
R/YjR6HRavT0iDWy3rMO0+Vc1Of4qGyIBFoPNRh+XL4k+e9MuEX3ekWeknY8Ask1
FGFvulTIacvkwmAhYXr/FKagZ3jHycRN4M35MPgePr1sWN4rCEW+ayp/FQ+RlW0V
QV3DoRHXw48bhjtj3vjJEmt0hGxaEHPLX8XxL0D8Bzu6hf1drSWWtZtSS/apTm68
MUVk7ak19pqFTcri1sNWqVuRdp5aBYZVE58VBKqOmM0xLPJpbh9DeL4qnXe5Y+mv
Tfna7fCalZy+753ATgEvcC/q4RCd4RApM8yu37R1WfaOY5N0srdFGrvwRmNwngA4
Vn34OIDotQ4qgoq1xKGXhGpSVcZbcKnFzwbu4nVTyGK5le+/OiwkkJ5z0UmlDNgn
kqD/FFmsLB+oX66AlrqUy/FccoGu4v22CYezXrWAnYDxTQOWOFGg0hAx1pdEolyt
FRQt/LXyQUyvCRNfsMQ02vf6EWIcND0ry7MkNBwZjL2rZudvLCgyJRECL+uH+v3+
wvcVW0pvskouXaKk3o1C6cQOEPxwnkmA+T/WOqJseVzb3f8/mCTgAKgAfCmlTmje
aIR0BdzcYgMaGCLD6uX+cMC/iGj7Z9Iq99iTOrQFBxbSeUDgTHGN+89jPUPbW1Hj
y18rPfu2sP6LbtP0mguyiZsNBoXGf8OIovwWUP9Yt0POn1cZYeZxX5rwSWtsBS9O
7LcaUdDWkH0s9Y2H9ArrfcBYYZcdpspNFKFrRx2PCVQEdQOqorl36J5PSoyDCS3r
mcuSCiauxp/NUlqbUIQ/cnnQaZolRZ0gLUpk8HUOAaw92yHwG+FGYTs5EmzQctnD
5PC5nV9tJJVivhXLzxnLhAh1LHVOfSZf3DMFvlLu2L11pWxWBU9icSvI/edATjHc
MVDL8l0ubKDXmtgu8GYhNfWtXjI7uhn6RMrJJluV1knQvAYcOyFekoETUiJip23J
88BMxDUWn+42HeEk31/a4/0CMmzGG3CLNd0/tBqkwsKk+BvG01b/vNzHMQtAuxks
+XCuzu8RI4Rxv9b7kDzpKqyu1PnRvKGFdN5dVk3XL/zz3ft2lp+K113sOD4oP9ak
t6KKKq8QEBwaoluazjNxO6sC9yhwf/u28U89W78Mv2XlB6CWAI2VeaQhjWiZZxYx
soMVBrFbFhceuQ618DHHVVVd6Z07NeAy70myqGIceBUSMMwaesm7T4S4FgKDMole
bNNfeiPD9C31GgDh60BRLMVWvd/HMhtZeXAqxGJuz10DFk6UfMUwdTbdmOWdYZms
UugKup6T6iq3AiCay73Wk8mAt2Cto+Y3YFL18xQVAU51hUIsbKv11UDAuAmawfHt
y47MXbonyyMacU1A4591Hj5AMdSB4XGOrhe3eIK1CG+ZXtX+doTOCRZEq6PqluxR
HN3gEIg34Imriu2c454tWkQh30uyJodtLyHEkrrpfEh/CTTIJ+7tP5uMtWCyc6lD
eD8BcDU6Eg2JBK51d8waa9x1M4mKplvLSThzN0DahhmQc4tonccG0JHkEVN/pL2P
VKyXqYP7tB8aZGdVLQclfhRSKyGWVSg1JKHCXfyiYUWSs0ntFn1i3lIJ4w8Hvk6n
KJSgCGT3DQUb4OJomHf/h6B0J/RjymdRHZ/ckT8GIPLLFwx3UUhMvzRZJmZXtgBK
2f9PihWcVgxS2AO4xw05fmkielCNTrRMhXAxtFJmGejhq/Lnuz8ENccsfpjnI+G8
XunNi2KMX70ADhDYyAOXC2aGRbZkyC6J1W6r5QDfi8UhJ4xW49n5VOOUar4WGAAS
BZrIxM/KhKogI/4T9QY8OMsrkvZQj3qU50cw/+F2iF95ZJk93W8xslHSfdQZkPN3
/qat4qzyZCtp3QYEDrBMrXbUXpJLA+e8XZMq8mviqsHWAgg4zlS27L8avo4p1Eeg
pD84qsvrqj3Blh8VepvGQt8k10NG04RNNj9e1YOUXLEg0g8EUnKC3Mh7giJZT/dh
O8Rx5t4s8dc8vKzu+qwRJ2GixDowqEHszQX2lLFOPOdoujt/ryfQhK3w2wKLo3iu
xiD+UW8nOiwYF3ucjLZR2jwTFc6yiIKlQm65ILlhiQQj2Wqs/hMWd5E1Pu0+mQZF
tiKl/2E+b+ebnwPrx6FlU/QpiXozmRKeT2gx7AReGRbIdQ8x6PnLd5w4PjD1ZXZt
zb6P6jex/dAx5PeYP2wSkI4IokzBbFMS1rKJqY7d7D51b5B+yy8VlQLKFHJb+93W
jPcgb5wSUMAVM8ihOBHWrT3Pmgzf/GiGkZ5BZWeVBiBMNE48Tk3ypGG6iXzq/1ty
XtzPAkg6TF/LHqIj8cF14mBvPjacnwdVpSoV+abzDvG8b/fpdiPcm2dnn62Lner0
DTYbsYmrsYeTW0v0ewMMtumAYi4e95fAQWyexj44lp7NCFTME50v3MgXwbwDYgZG
hxZKo9XJjDGQmLoivkSB0tahmGxpypxCcuuFpspLfl76Rsa42nS6UetWFtmRjX5q
0Oa7rw87RvI4SNxHeTA24llyK91fxpjj5bO+yqV+Z7ByXUEWcPil6kO7+B30mqYe
uk5auYO7A53JnbI7yy5cZTkpHyynVV/gAeTXcXOX68zX0hxkn82SpMCxIsV1qrMW
iRoiov+UQyI81RSODkduXLuLLL6Q3/HUtQOarleEyzwUBI/vkAZlpN7sMLjrkWDd
UPIlSdy+3csGHas1AF1znG512WV+du2sdr/okjfNA9TuCfxnl7wpGqHdCJdRXUM/
1b2izPVHiWi4E8mwhjtuSdFwkFNlLU3Nk+fOdB+pLpp7/uLPBA5PY32SB/5aV1I6
jJu5pymucSPqIpw8HMwk9LK7Xt8Un0GiXJVBVWGzjcWcVVgObASqlOzByTPUh7pu
OO8hMtL/tXWBji7g/9SmxQGLlxPfjN8noNdSRrV7WxPrLVZGTZC1QfGhxRIZRIA5
/cVdb1hDDXGeTP/gJiIVJcc0tHrFCYFfUAolYyhsgHzaOeADsvZ/goMXVwDpUOcc
w+f6j8CS2EA6Qw4pZNXmjmjUb0D5nLsQkNCtIsdvfoxsEeqKFIb+HPaYP+qfVQ5f
plVs+Yx+cUjixF8c4gEZp9H6YnSJO2e5EQlMLm9Ha/NpN2RiSyQOU9rMh/YXTOLL
WUme6iDST2+QSz272ad1YxKbDaXqrJI9AFth3fNd9/kGPKiKUTdSTQGxS40GZDzk
8F1hZpeb078dHwYWUfkTLmcuwlc6Cephug7ZKzxZe7obfmL5H8fbxNG0S4eNMLRM
rI1AJN0W+pbWqCxIdYAo8R+FQ5WQ9b0Hco6K3BjG46CcqBtfo6NLvwb/r2rJeEN7
dT+QSKIwWT9zj8WabNBu4W43NZkabvqshFixeo7UrCN/SbrPllNqZB1U02XNSfWG
G5sghXx31gR+um+iDlgSrbr9EK4QLA1Mw+14prYUwJLwM22CUIriglQoSGGNZYRS
U+4iWcEpaoiIKKDJDtDb6pbQdFyFBHrw4Oyavj4nj6qodVyYB3WghfNp3Y4hEqsT
JKHtpqlpsb9pyP/2Zvp6Ym7MTMDKip8p79Pu0XJFlq3XoHPesCzZ3c6JU3min7O1
4OH885ueMs9JYwhntX0PYvvOdbiJ0kO4CEwQfJiMM5MDs0DBgaBdRL8RwDvdqhkN
j5XuWFjWoGFeo04XdBLO9ysqJGchJplKGqiWQCBh5X1Ksu1uEG6mydi/Ky5Taiob
rkExsiYHCdLTCHA1OuxkAGvI/qqlXY2cagKQ7nyid9gZH94mbyJ2kX9f1SNUQuEL
3PZjxOerIb1OMUTnZVp0tD2BVy8U9P49QY+RChQnfSCH5YIfPuZjm/9CIChQPwVH
9obeYyLKgLj/o/P+xOJ2aTk/j0X05GTPtJUbd4hMXXhIFvjbcRKkTpd17NRzgyJf
w80NdDYLHzvbUAPCYdYjy729l/LACUHHIHMRPxZpbSdcEyOWoyhraID1XXLs1MYA
FC4SeN5PCm3vecRxYZg/MEsJtsQI0mpy8UQNZeN2shQ1SGrjlTztnN0Riq7NMVei
fDE34pXp3i5FV0u86glPheMkb3eDg3B7jqSh9+G7DSDT3TZrlPNAGeuPi8H5OtwR
E3CJ5geLgLHphhLXyQourVNump0Doi+dOwifbFn1cfXwhYoM3bH0OOA6HcWFgC8t
vVwhjOZ3ellPAzEm3XM385AL8zgZli6BfCT7Tvf/yQtNT+9PAeuDwN/mHwq6S6s8
K/Jzgxm5X5U3QoFRjT9aV1ppjemLOk1VJJKTHTl5NqM4QCG+WvCA5vCOsSOV5Xf0
HynUtrdKih3xwp1jPq3zDrb2O6XZ2hdm9+53JqUc/f4hj85lu/hRdAX8eGZgKGWQ
S4PBB+BqDY9+bP3VFzSEyrg3qzTsHYh7WRX25belqiTESvrIFuUqND/Zv4hJ1Dp+
s/3dtDREF57oJ04WXkgU407cGETEmPVfaE0SL7vdXdd1sLIh8uIo3QuyV5OFdvRp
3TcYdV4/cdTun0LOoW4Ht6zHmP12VB912kL2xyYIh9xDuEMQPXn984cZbzKrO7Rv
wLz27FVIYgUg/qjavcVQDdEwELjeUefzo/L971aaaBvoo6jo0vZQappVxf3oaXn3
cM8GOThBzAsrZogbw7h+dHnqtrTkATsQRs/PReIwP7k2GjX0t0tMSllz7RUR9zH6
e+rK4v02591UZiKQIivStGK9JQeoeztH9Ql3Re3Z5V1CsdGsl8hLsDAbYGYZMTWn
oiVSdHHspxsKaRH0ZU6kWWDAe9ka4h361wa4ynMQjlM+x0yI4g8o0NpKPeWHdXad
2LlKXjNEm1lGw/VsSOdCJBDxltdMJd1d6paoIkC8imnXFkwlIVkpmlO/uvJDK8H5
NMhvsB/lpt9ZbhIwukNPORX+y2wyXoVgtjBjPzKXSd4k7ABWqiF1NOIzKUj+/bnb
eeQNp98ylLvRrpsvYLsYL5Vd4UuBF66K1JToirsB43Z8FgLvt48+nJQgRudB7otb
le6jsyJZchJhAj7HqLH9Rec2Cd9zTc0jNOl8CGcxOJT5G7LYYdofQ/pDeJkP+lxK
kqX2ZylhwKv8Gyw5ziTnaGTY3ItBC31lgp0uoqboaCOEzzpFCQZZ4xE3QSZxyL47
KuzPVMb6pUkHphu5YHyVns3mm3lWfHq5q1xE4ELGQUG4mR1jzxcz5S4JkRlKfNN0
rTp/4lplUIFbUBXTTlzG65881jFictEj1ybhZtnw5spbtOFK6FndvOyefh4KHbVh
r7aYfFaILlqXbaV6ChbFBCnWgD+as364bMRymwNxZzcesp0omA0P4r8VRrs2tZj8
7cWyJTCVDLE3ufrRK0C10bN0xPeObbiB5riSJRWyMLed5XoLQvcVadjyjk1c+c1G
i0L9XUmlcwTvj/b2mpzJkbEu7eke/QzIWxK1DyfnPOW74SikxZI0kUeW8K+9T4o4
ya5cjf0Gt/94MCsyjyyXSM+HBIEodvbb0bNBskA8MBY6C+g1o595FZnENUrvmJ7I
AH9kO1iy2KRPCY12S74sM8zjkJGLNBbxwgvVNfkvFXkz6WQ0G2ZLGghYIOKN0A/w
IgFb4HMo+G00/i9DVUt+7itmb3kMw/esb1IDb2xm0vJ7RjDQE1aYxZg/SBffQL0G
3OYjXaCkrUBDIQFE4uLm9ekxOJ/4cTuwE6FT6Z4YIXArXGDqLBMbKSmbzrOfMTeh
FWJCGQj4rfetSjYmBLrICg+FjL+6LVyY9sVbiOHxoKKgfnHrCqHJcTzMFhOu7R44
XzveIQFvmdlPWhv2tdnnxwdQKsgThWwb9v5LZkfSUcTSSeefanEEnXwnGC+KB+e2
IYzOsmgXSyr6e7Q7A7/I/dTYGWl3cfjmjnzCSuckYO2usRUGrxBQOdxui42eLIZX
NkZmwKhOxBc5PRxHj/9Hy3bu5wXe5aZqNRk8hApKCFhfEkVAP7D6MDzPfidqyS7c
oJ8nhGamGAWJKwLz72+9jZOeYoFq1EvPtP+Yk2kfsDXzjon+90aVEL/owdNOQL9x
gy8B01GXKdCiXBPWnq6Bc1IjDXRYqpwAxLbNrdgkV23KbNvoV3HaEkUmHee19xbI
zVtFup4oE/FbgqmKWEeun6ITLkfRqaTbyP2gBXEzHwtAZ4cHjhhgr+8XQ+2gbFRd
0nXy25HuIWuupM27JBHOUdjg6AQHFwYua3pAT0+b+hU38R2dgz2LeUhosiaKg0LN
3KsqLxuCztAH82uB6H7vmYu7Lry4CRPuKVQrvEPPltVzoUfyAvbvLF79q8YmBgRw
kb9iweCjWyUwy2QZhBRfAptdI2Rk/6bUXIVZ6grM4QFPNel/bzNk/QLuapxpDEd2
Y5MxZ0/TAX9bNz14bKHyXfvSraVzQedWPm/OAufqALNo7iWkvokl8hp1XbPh/UdA
Z/tfGGgy9cl0UqHrWNblX4OkeSWWZh9se8zAtufYjMz5+WgSm3d2mCTQ5PV9Wt5R
BxeY4Fyv6VU5e7xF1q6chkBTiG8dkqqGpJUiSb8Ox8EYcCSwDvLs+e2M70waAY9P
G2yqDxmllIiY6Pl/SdLwzA3cmlvWzDGlA9zXVOUggJnn1hItPAdiKwHROznMxzf9
C1VZT9l/EGl3kxZgIAPZvY2h0T4Z3lEe2dAmjgYvbWu6z7OLOCqEUI//U8Yp1pOR
026hZSsKUJNL4s8CTNqKPr64Wrxb9TcT5c2MWo30fxVpJhnUyAsToDH9uSJY9HDy
Qwt6OI40BA63paA6DO7SCWYv7nhgme+NZrMgH1oQTm6k+A0ctA9Mjwyq5W1ltUcN
3Zw4iN3Tt5aRo2SVwXQbvTnHkpuV6VbO6tFGDbkykFggN0Tezyw+s/l/nFQetmJI
cA9L7HRDpJVKT1+pNZ3ZaCYRw9owGziqhi7P/rDtQZg0zdduB1+ON8IZx9UpJhOG
8LSIw/0viBN164oKijP9RlDByzhxKzjIpd1uNqHhT4p+27a0Zg6lK6DZLqoux1Or
w2TAfBVNUY4a7u+RZU+dkTu9NQYJK3kRlLLuKNck6gQ3g+PIqrlMK/MIbwl1WpFJ
Mx28J/vL4b563wY1mcSgycXSw9HZLVCgqlj1YHpjgPt1LVA/Bar+/2+rWqYDLX/h
v5MmVHnUoEMlYD3Ev9yRAGh+sf0B6t/45rQexAKEIE+WqlD1PZEeNBhk0sbIU0TF
hFplrCvi3hHbWXhF3JA2FvLcq6EYU5ctr5S3N/Fn2LlnccPDcxiUqOG0+STc7K/3
ZTx2iLRIb2ODSHlAgPTaVYvKSDI43c7wRWOGrUHUiiLadf4MZ65jtCM7lE4BjTu1
7gSowYix9bhHoTiETQMPwm5gxqCkEIPFqCZgl4ESNUwDA/KQogZRGq1bUqfEmJ1j
VUReTni1u0xxXR6xpUsPeLCZSs2sHjsY91yZ0KdUr5CkWwGB7bAs+r8B48Y6mhQH
8t/gaXaTzk3+EJUpQF63Uc1fVU8h/hhZmlnFrPtMHA6+13CZYpBp9UMuPua4bp0z
JH+4W7AkeTKMfLi8eCcwZ9wyuG48dBEJdIPfCeuhU15qIxFpfH6VXJ7CtcV9AjWC
qLmssvZId6bkTFFMcngpLhT1BtltDUhK3hK0ZRTbN8AG5Yz0ZqqwWLTHbg+yOfWk
f7nSL7327RzCeeXehHkd05QLQ0kKKwW7xagiEqiLCT8GHMw4OrDi12vbI1YguZ16
v703UoOUdCuLm09U6tBT1invSJN97iLcBKdS7LaujXApZv+/K3gGITABYtsk8JgB
Lz6jWssLLrVWeiSxCc2lUF+VfyzkCIv98cTktaa8ZK7STsGTYlcF/oSZtfP6YnNl
cUGItCJx/o8AKn9nrnrOm/JTW5ob87x6/OH33Y77pXYGDPdSBmrk1NWzhAAgv0CZ
nmVVYJehBCrX1NRIF9VBzopd4ivuX90UhXxCTWAK1zpB/F51U6qp62xkhb/a3FyE
MTog3TRz5C14QXbBhSxY6AOPEmTbsIcWOMEpabLPxAdKi6GT6vgxmKSuj5b7ZoOR
2PFv4DWeijDw/G0Y1iFoozLIt5qnLUuNJU2wgN7cKvLFQBLprqLCHL0dE6ZIDz50
w3l1MZIIQu3SjkqOEb1xOozoONzoTypliQV4KhlsIvHgd6faZhLwLtGaetY9FPAc
sibm5rV0o7o4O/gLnegyRMA27030CW8V1qGyLMhvpsQ2rVekiEy523rRzyOhjTOa
I8Y9G1/IyGu7/7oQCkBLAkRNE6hesqFPY9bk7bsAjUOuWCmwVypI1ad89kSyXREx
i5NyirLO63hrgTbioOHLFq0bosD4tVb21C2Vd4JL/0NTA80G6HamYWypyLKXwhIB
Oii9FWLfiRS8MHs02nocbWDqTRgaT96NDNWC6INy7eEGQ2fsE7Io2dE2g+EIDavl
4a3hiuG0KYaP9Yi9mZT9q1or1wOJASvTlFj/Fb/B/3oKFe3t0yzrKYzXhCsVeYnl
FgQSikuqY20s1rmExnN/T1QflgkEWkDuO2eUUMhg7ccRmVZcngRY9akiEQY/Cmoo
k8lHbPnjno0JrLdtksHd41YcsGLdGfPyN0l/5dYgS8o+Z4HsZBdKq6Q4HEUDjXEV
xwTv2c4EgtcvlJI++NQlx2br+I1YFzXjNat677dDAM0+sMmKxfCyZ/tJl4fGCbpn
hd7tkxPja0DfHDRlFvbCIJ9w3x51ZRBzIR5HrjZjuN4JUL3fA0R0zxN51JFLUInH
yGX5qBY6PhLeYs4Ujm2o7S5HaJ+QEWThy6hCnp81ddt5eVnNu4Pm0ssfiI2XAmBl
etVJHYuo9RDhKTP+/cznv+U/firg6QckVMQW0POCCoZEAK0HPhvAIVVeFpGoL8+e
jRI2lZMc0HLgwg1m9bhWOKMPnA2PINSuB+/mC2b/9GO2Gm021o8TO7K3Csj/zqZW
cQL04H67urZHrypq6yVrXKazwyCd7708DL2aufnEkvgDCMXQEuVgSobZan70jByR
HMZPjt8BgPOTHiTYQlU0A2ldxI0yojAS0TBujXGoU8Ko8/I7QnBa5U6uC8rS3bwr
vf9E0K8INxNQFtsNLvsO6vmRH6suyDkHMFWQlCSnUXTullzE7VUVA0JuuWIW51Ym
bWURnuDWyyqssLfsEgbOFf3zO3YXsZcwycuIInggfYtG9Zddmrk0w2Dz2VBXCSPn
5KK3PRggrokjYWGfXIGn7h0KyV+3Dc03+mXWbqDZDNdMH+am/dUmrNaJPQzIjiEl
c7WlQQcfzi23qwHHWmUGj1kFO6ShYuPG+J4iGMnyfsns7Srh36tZ/1bbndaw85UO
2MHVka3WbulhahrdnbGT0aqYUvGoS4uWK36KtgfnZzkyzINrqhbK8jmwbZYKbo20
AJTx12ttnKnri/SEmrlVqaSJwont/4PKbBWjK91OzPgjJS0IkDxTg63xWf/CBNna
kIhCVYnfDilBEAlvoFKCk/a40N6pj5sTxdDRA5+2QWQzBIw1NvCks1t0HWW/BftS
6J0xaQLA+xrJFC5CuBYifsQTh7Sjku9lmPQke/e8CsK9IRI0W4E9Hei3BOrNSdUA
AgOfZOoqqckzhb4RjO3CjRZW2XppxQ+Mcsgm9E0yiFxASljHZFA63OF5N8fd9yw1
sYZuGVIbmCB0v9oW9dd7Y4UYewfAZb1NWRHcT+ZHzm5umzw8CFsZVVF+wakeKcqn
gd1rcfzCmtURJhPbAOWQ+8jzGizfe+uv4xi07dql9jN/5NFCGsYRRaXIr5ZQmMOF
97TiXy2U7Doh74AWNegyQc9gjGfLWYRiCklCtTTLA8LdwzoxAKxsgR0SmW+6Hz2o
tgdSBTVBgUYf9euB74/vE93VE5+QrtV8ewGj++cFgkaiopb+px/ccTCPwXWoxjSz
zpkNw3gL/GbwD1cLBEGXQPYwo7GFEScFim6+lwGyaSJLjWng52q51Zdpzkiylxf1
YkyDD41UZe8epcnmAUBn0KwafrqXnK6uhc2a1uchrPuAj2lOx29/9cBR5Aof2meq
f3Pgq5Ht3SUjvD9hKEPhYa7sLURwn31+wXmXI4zLutTcNMylCgO6d7D1RrF4VATq
tzldCnJ/FsEtntQGXfDAFjanjy0SWemNt0OiwgtDisox0VwjFeQEwQTHPidLUMP0
bRq7SH/gb4zRyGzUfBAqL0y4UCW4+2YdRrXrhZKFgrhd3CYji6duqEogiz2Q7MZ8
Yl0bzFNkojc7YSe7AEYrVzrFjfL6AjNMsT1c55SWDOyuOwQphLbG0ASPxoIm4olj
ufhsxVeIccLTJEQhVkyDS9pS30cOjZG99h4k4P1ao/1V2C3OEArTEsgqBp9ohUAM
ZS9Tvm5kwzYXBi3mQUeVhetJR4Gjspffx4Q4c/fFcVD9ZlNvVQl8I7w92Z+Iu43H
IsbLwVBbmue4QdopKURp25hOHNvQVFnsFKtI4barcdJffQ53Tm2M18JMdSxkX4Dn
nVouXWEMaXpn2wImanjeZCrQ6BIZmd6r4IiOExEUJZnofZGaWZwysExRWH+lQSsr
qD3UdpONtpNBXisQXmlFc6iNHD7SaRkPD3FYaIyWOhNtifOuYyD3ciZIPUYbWHsv
cpFSHGU3hEtxiY4rU7UzlFK5MwL691b+fBeuLTAXFG+SEEGxs7P07/Iq+By8YfHE
yCwSiApsICkwsVIjJ+RmwvzSlknreW71RWR54g165yVXN3QWSgm1BWL0AydLr1j1
4tIqnJLQgn8K1FXvetBM821ac3ypsb0Q+nIeHAxcvgGohkWSY+OVzR70fFrmwUZ+
kjCBY2ze40HlVVNJy+cIy02PiiPyjQiHRJS+Er5ZjFrlUPOi1XTzyn84ajiIXUqh
pxuOHK2P4HYaEnNaRFf/Pv1se4HPm/2vowxvV+vdfrt4Xsy1OChyKvGNmFG0FQe/
QB9ZiKWGkk/5yiHF4PKcoRz9JzysdG0LbNdo0O0nRTgOmuRZ8VqeTsg+NVhCOsZA
q/mNJePZehKSSD0IDK8fM4rRCM4noH1gs0cNCO7WJWiFRF1N1qIEq7afPkkDfYxe
p3ZE6a6aZ/y768kbHHv93suIufaJYuWYQ0hH7KwKDXlYXQL/+XdBj7vVgLloEp11
/t2m9B5ly3HP6HrInFZCXD2hsOcW+itBiNKP6P31isDmQbjmKzhMBWcbqHjwgNKO
onBTYTJg6Afam6k61wSsGGTpU2P5bqcbVfpA8kJZJQzyzeBcbAnt5x4fQV5+oItO
mPLF8TXMmcZvUbOAeTI2fb4N2fBWtpW4Xi/Cw5qPsw03ktLKKcWYN/gyZXzZ98/K
w9OY0N1hfXKqDclKQANEbOPR3u85RmUBb9P7HFq621QHkeCreeZBYNvQVghEaqUs
G+xgRnTg5gTuQhDHAYjLR+CRbCn8MDZ8sEt/8uRiwn+iY6iWwCdgEVKzhi7LTXsF
KWKImof7qdfOjkRY4hA19xoO8hqxNK1ZWEonAGLkO8XklSYOFdseqWHq9SpHFC5I
FblkMMpbBj7KqzDs5Cft/XhQcPlkRyG2FMFaw0qj42jmo1vTb+VXrttHE8xdOzBN
TXd/qDiLrDH+zn9sXucrE48Mb7c9FPNxRELtwaY1cPVlfLT9lReI6stnkVqnDoJ0
OvM1dpWWW1ssMo76iIvzyahWyYTsI8ccExv808mWFCp+kpq4Yh528SRhpoirs3RH
vlPV9vshqIrVAyAP2xS27RgkC575BFw8c8JPO+N3hH+/EJQMAAWjWVmBg9qBaMUQ
r+uJV9Z07/PIuqd1NOct6cwdY6YVKG23077zxVVyK7qq88tRkVy3UdEFXaD5O9z3
LymDjxap5wXywuNRuFAtOIOVf31XhGBZ1T4n1BSUqNMRjWfEF5egQQnpouU5ZZOW
gWxCapESxHL8zI1+1RHJh276K2jNaGLMWL+y8xgcTKr3eaaLOrQXWe3zDdhCuM8y
TYzEA7BpTVzSFFqvmRB2Tui+ZJzoREqnDL6Fz7ixt2Rqk7DlPZ0IVR6ZGgCmja5N
6/qgnLXRpVJE+lVLuox8+rzIMvAvo6rHbcCKHIlyUzy5sv3MgqcYq5fojUzwbK7v
kuhTKWLQcVSgHzj3s6mgUfONMW+g1oloSH/iNf0n0DH4aldxxFznWMXqBFPl+tbA
+Gg0jw1avtfGesKDf6KlXDKLw/g5gauXePzwSk5znNdK5TqhzXNWdUZdLeN54Nht
bYH/ZNDJj+bzEJjT8JMcF+pFuKBouBjNWbTFgnB5o3qHElTB50J2yJbnOrZCGDtk
Qop9baQkZYD7HbU84KaHAfiNao/DcqeaP8jCM1AJhTPHJRzVkfGbZHUDRGVPcnds
qexyui4v3loJFO//+lRVGP5nokSz2G1M5hMfajLpsbDGyVBt1BWbtQ+Il5+9ia64
f2XuOEVtnF03yBxpsXsyHK+cWHVs0pGrmQAuK/GqTFlQgd0XV/+OMBC2tN2f/4nh
qp9apIp9XgMG0FpKQIXPgjYQTsTgiZbUpsEexjj4zmtpVeUR58Qv36a23d7W69dq
l8UwEJTypG3QQOV1Bp4FRD07yeeHC6qWPq/EEdV1PRCQMzxYk7E+/HVcoMTQcve+
0uX2rzGQ3yEpbYQxz3vlq+242N9dmxaXTDKKlOPeOcA+7TBpnp4siDiLju9zyY1q
OY/qyg919DmUmZW9yMshlYuhkfQZ1m4ko2BaJiNqrl/M+0DP6AOwiwCj3Dfd/2Uz
mP73rTfoMK7JHgqn2iPAylETFwEUDdLL/cPx2BfDzggGov3mbrfg2ujvpfgvvS6J
qvOft2ABiAyc7ed60xSTOJ9ZXDqM1RR/S0KASI+s84RLwSvNDmPznZBdY9T3yUIa
GCzzTWO+s0tFli8UtXbqNyTrsAiY9TWr6eeHaQcUCb8i3C1VqiwplWdep1D2hLAH
XwTsg9RkU9Q5ylZA2QGjWEQZN+frzA9FLDMzstbJ636394NfsUQ3hMnFW3JtI/h8
Z+zVeeo4glVKBgbexG2TbJ6ZQA3HZxZwistH2zRhTF1qXP1qSUjL60QI6n3s4So2
dn6i0T5dN/JTj+BE/ug/eCHBKrUV3GmLkHSHppssUwCLb6BOZ6nEMbKqyAe3v75K
HjjpR9plp7SvoGB/S2ac8MIfaA7Y1eqMufDm3whXZj+AcEQPZADcuoBEnsoPe0Je
tngNn+X9qU+UZK+c+2ai/FjiCSTPXrHlmc6PVSGEBN08GeiwHfpBPRpqIRAgOIl1
/HPFVlWlRRFXZ7fuin3C1u+yod12duPhxDQB/khZQRfA9Pg0lOpK1Kpf5WTjtfoA
xUR6RzPXKrvccg8Cx/iKYOpdKXPs+U9UKSXTRd7wzl/Oe9nVRV937JDs0lHF5Ovt
9+6EmcQbRgdqT590d8T0GWYSHps/gWO2wLmB1u0BEqS4Rz0Jnf8d7ykV6Y+hcGvQ
5agmpG2HyEaI4JQmLjjEgup0Kl0h3H5dPSSG6s1KTgXSVYjhAyxVFniPKejXvdhP
jXjo772oV0ge6fJb2G8LofiMe/Qkwuu2SX7LXlKo0K1F4wiYxwEZLh93RQp48+SH
mctaFlZ9VBxkdVzT1WHamrtLbm3UCzWGjB+lA6SKnwO174b6zcwzncO0v3svDqT3
DIsk1y2QY/I+xZyOZ29skSsyBVidKt5llgZGBOkX1jTeBXGVv+BZTqg6swa82aOd
vjylNWS3It1TTLv0C71aBAg/qBW+Z+vLoKJVSodt+LIjYjX1sKf4F8BJNmS5ULEA
G4F/ooJTA2jJOcr73JKSxyj4tupMnK5w18ke0T/74sDJ/lnKOheLL5twty5cv/+1
tmfEvKc5vHOWL0tjgd4rLKmSk7Cufh8XTqw9igHW5Hx9tDuT8ISS1/AgNwMLK5uY
gCFgYKj+aTMmBCmR0AxcDq/s2wEof1svxledeQFnMzb/98/DCGStzncRQkEJdKcX
IHt77WNx9Df4z6HqUDnBLy5he0Yt8qeCcwmji22aGQR2ijBa18iOUKwBFaBRCMKk
8R1zIMMUMqk40XPATNTIBCDU/vmOwK9bcY/W8KH0ZE6INVnu5YZJbfKQgxIEau4+
YuxnjdFGZBs7tfRpevwxtr5n2RjtS0x3SdQ96pSToeGHBk3D3TkJVUO9Vqs1tsk1
x0+mnanCdnW7sH3sj8t27Hc08GH8QsLCJj6QN6BVpWZLE/TeTLRmbRiJRnrxP/I3
wrwlbW/1zUd584+mLKEsVxT+6BCkvPz2HBVOL+fsvZ6BZqnfF6I/hlLeNXdZcUb7
CDcaZqoCH6dm5it4ezhntQi6+3466gwfTW1E30IGF/GRTh5NzHB88Hz++JjcRg0i
xuWsnzK5RL9qs6RdELksYDWe6QKl2l1XyUJ49iSbm5vHtfVBNVA9qHwI7i8UBht8
Wl8JxnVr08yjFwiuA8NI7SZOvoA5oNy3gX5CutVKSvutV/jcyI+F0s4HVLNKuCpT
L0PC1Pv0c4qRpTCap8MuKGH+PN8T30dWsiAYxIk9Kj/awERTfB7PVtmCfNvOQohX
DfrVFZuN7/zFuYxSe9kuDOS/dckHWamRG7WGBZav7BDJ689zkONJ60FRHGrpLyai
hrL1UWfMPxNHlLD9kHS5hVIKuUQQxnwkSS5APokSSD9ICpMl0SMF43iG/ZHSkOu8
Eh5KqwMUe4L9fTaS8DZBZpoq90Pp+sOr8b2dpt5d1d2RY247SluzjdNpqb5suZSx
5bm1+Ua+RU9TXE7Y7wQvR9H9TYe0XKeFFpjFzlDeAPsTw2+OwZvo08Mo2OvZwrEm
Mey8QALarnVkrOE2tyn9WH8F18jZDEZ3ww/9hO/fwpQsdBX4Dlxy+FqWViLeZNNw
1z7Uc2FD3IPNvT8dmPLKuuVmxUDGf35CjG0w7PV03lx+rUI0US2JY4UhHYQtjMLO
i1OuEObL31YL+slbkUrJlUK+8NfBEQzveSvLKe8hZDWNU2VGRoQ1v8M7ok/MDP/C
o2r38meVYwJXlMaCNqAdj0FW26VCGltXKNDOLEKonsl1El92U9msqiHmzSE3R2ul
8skVYRwBYxzbr+HENT0sqhSKU4ZrG59yyRTAk/kv9tH6ppQ15+jjMEm7yhHt3xg/
2EeBTTD1YROiJgdUc3v2+rXeBdKZaNhqPUcLeBlvkXsuPWHS2f2zZkjUtfZRdsut
iWW5FsGCx51qJ7gA4IfGOEr+SiYpuEZD46/uGZ5euEaHlw0KCCMYb5xjCDHtxi3L
nl+Q/F501RD/7YNq3fpYcCRAhFNkv7OsuvYOq7W1HcmIvmm1Dxza/+Eth1IovJY2
DlX9jdHsK0ZANHn02C2bvr7u2QLM7RAeR6Z7Nxgi2jqcf43KaAPOEB2o1xVs4K+K
uhDi21PgCRrAYWMbdxpE/rkgD8XkzkfiPkVK/FctxeDivc4r28EX93GTVX2f4K6z
tanLF4c1RsdJFlT5+KdXSHJQlN9RAfRGysQYCqQU2hWNsVBVzYwlMwyILYltsKGV
zxKS5wPL9ri2Zcjac8vVrOeKfTB/2jlxFk95wfXY9VU8Tn7u0NOx+Nzh9laBMYYi
idCMJeUTUDL7yj8wIgCqq2zyMb0duBJg3k/sCSHsaF8B6LUe/2GtyeB/3sSkTlXl
ykRPiY2NHEa2RBajOwkzvkkZA4+Ty6BK3hAIjvpcsJd/BxyOroS/LC1SJW1rCeWA
SD7Afyz/pkSrlrO0/v0C6rWXWMh2w/MFblGF54BDZVaf8eb54L6/1POiV/spCINW
lSod6lk9TxyslY0NAFPbq0hbyNEkbGBXGppn+qfyBkRq6uwKSbK9YsSecHryLteq
OqGAWtKuP3U/CvpMoQQwEtUPVFbm94DehTDaxw9yS82o+05xl7vYM0++4triLMaQ
ufj2g2Qc68HjsYw7iWLB0EisdGtL1/2ulkaC45VtNG9t9XXhs6/S3tooErBXqGoW
1bHImHCJGiM6y89xSzpvK71d3OWeYqsiXKEsyZjwv9V2J89IHD9w3ZRi65+mleFo
xM/D3Fl8Y04/ewm9X1ncIovfQ0ldpVk0AdwDUTlWt39Fl46ax4hbQzUwQPaHj+uL
HLNHrWdvkOt+3YDu5LuDZhsBZI0kypL3RkzEAgBlqmF5VaMP5yMf91oi+zxTT7a7
cn34kENo6QmKjRvef7fN4lZ/hqzhkZQW6U7Ca20GBApqG0fcXocprcCBBev97FG9
VARb98b0yHpkFV6oUBBtlv2Oyr1SC3eOi6Z4DoEyYYnmHX0EGLesyXW6s+l/lur1
IBZPAMxWN2NF8DClZ3QsfQOqexhXLHMfjNCHfg/YJAZjiyVhbAfnuv+OZ1fI8r3e
lOD0kwkTA00gUAyZuOEqwFOHJSEJgAmGePaT2HhVvahsTIdOd23Yc1m5HIqm5UgO
Fci+8XC42FSzRhmVlCpTRQKi3AY1MgQw920yASXcTbuQ2Tex8Rpo3vGKAlGvmouB
60xn9AeF5VvBKaHE/1/rHBZUlqsQUeW0ROoWjaUPTxkfbDoXooMSw2QlDkCynU+k
T0QfXQ+jP0MxazjnTCleYzcCKChays9JiVI1ONYW2/3W86eMYw1Op0MVw3wrST+K
BRl3VI2qtx/M5JUfwtq9bvGEY+eUSLVDJ62+jUZ4lktjIFOvFNGnxTH3OYMcXoi6
zIHRLCNeLV/caGIpz84G+jW0TUSlp6YtK3cpdRRXLCufaxcDGJqnRx1qBxO4bbgx
EXuF5zZc2SsVR7OmzbbhFUL9+b6u2IR0id3eT/Yci4S7H18TGDZv1YVDULXb16v9
jQ4gxNvh+Pqt0eRlinez48ozX+30tFsuZeVOs+xez7QFM/1RTahB2aqTq4UZJHCW
jhumVCCRuKRRKkCvZ3tNuxgO7ZDtbns81TwpoxDVLkOWoNhQG6Wjuh3ZYxknC5OT
eKdj/vP54c/EfYjnRAUrqL3jBMMmC/NB3eB/4FdkgoMDI8Qhnz2FTISV0l0ET59B
PLEDX8AUwlmW6Lh9e2rnaZDwtpRc+PaOtY2pKQZFOJQHCRYlCpNMY9mDSNLs6U5J
KJYNYMhg8K9e69sw0zU19aiDSq2BZjZY1v0saeHT+Cxw6lhvFUuRdG72TCseq+Az
fV4+l4XjCWEcXzm0Zb4Oj/1Utt1j3z7rRitosc2cjSOErE3Ao9iLhcP4gCZf9rMl
4V6ox1+yrfAx54StkoXJZErCQNJeZWr8zfplSI+gPSbpmlByWsdarnlhLCpRq54O
+HC9SzcOILGJx7GSIJwSGr1zkIes0NetZNhv0byZs5rncZSt0CDzc2Ui/e49DJ7o
vX6nePYKTzVvPTo6ylwJPMuPk6W0auRLJ6Mz6Y+oEvYq7pNbmr/WjqoosGPxWucw
WZQ3uMuaeqOHqW/1CkBwyyfcCoxZJuG+i+VBYYRGTlHZf12Q04WOA6K1eH4Mxs3m
GAAq07YjPClzbYpt5sQP2RZ/RgKY4Po/UArFrET+eG/BvZcgKCknErx8gWaW3fa3
MuBmfMOSXZBBsyMspTu49bEV09/S43h+8EjHWqUFusDplMs65fhBP5Vm4yx5t6Rj
qvWD8ZTQsvVA8LlMt5tZ7ZD2PQWVJ9IrG7NjLPkk95Gwz+AdBkE3XptUuRqvlZ01
DJTEDomWRp5gDE3la90pM6MsWV/rIiVKUvbNKpsmzAcYBU80p9eOoQ9eUVnJ4qVM
ws/TDfaliK5WQ0msPKql341cdj9pihT1GTnXx+XbKZ9PEtvCQLCSroiaCB02iapk
2xh6icUYljf5mDp4MJ06YF8+V59xRUzlu9yH7QrgwWpQUMU8T825kGHtjJ2fUasN
gPih5fkGvQopFAbtrjGTKzt5gokzzOC8Gbhevf+RvHzAOkydI6Fib5wWAdH5/5EF
dhOrMiQawQshsbI00IcxL6YgLGZTKnyc4O/TvtwaeZ12/YOLA/PTWQlMdp8z+0al
suHf066PG1ipZhgnYGoMPQV7D/jW9LrNc2g1g+HJtXR0A4GBNWTHYg8HyEd5E3EX
3D/y1HIWCbFkKezujvgrEAAPyJvWftvbTmPBvWB9de3v1+EjeFLDep9VbQ7dictJ
aHVD0t3XqVX0hBnn3/0jj5pK7KagyvIz9Gel6QdLkY7FbRNgKeQnYipelK6Bs1Rd
BkkpzdUdewMNddEjn0qpN9TmY4csBb2GUHCO9EuGKT8balQrCnVG79H6StYf/Zol
Oqmq9a8+omfe02xXo8TmKHYGOVu1tIM99VkHtfd1ZGei2UGWvthxkClDmR25qIPk
92rFYyTtYz/fYsLf262Z7KJOQ1LJ4qaWOWPZbVM1NbghyYTvhNzbsew1OGAx1ukG
gFfAyZ1ojo7ZPnNJBVJ7QTJhkPpU/DnlH9vPOf70W6ymDVN3Z2HtdPxZg+6fdbln
L66tPfFcGy9yuBZgON1JWOv2USk52BzBm53GhtjZof2jzaAEXkvvOJj234IQ+8e7
5/Z1aDkYCBDBaSOah9tSOITmYOpRcIgbIBrzGR3eVt9gfIiqDrgCtzng6uTPTEUz
8GjM7fOxti9MnzskRPFJwpYxZbaiSJhtOK622zBQ02EoR2dxHhPGZF4B70+5m32O
tCbC8AGTZotfZZjHN7+cf3uf02mI/dpsnZbb9DKER7D5c5/0r+Td+zREfeEcDXFj
OXDQg6Rw2gvfkAu238lvP9DLmu9HBKchbmxr9snaY4HWjP4S1Y/g8xQWOF5khJFw
uyME8tDJBaonkhZNPdBJEs99OTUekb1TesJyqgNNgXiDUjjyxFs9f4+MqAj/rwoB
diTSA/xfiicaGZadsHGd33JZLk/ifcZkDPf6kIatAws+ua5+9LLN+wBTMEk6bSc0
DHqHh2Hk2EoWx3oH3wC8NrBsKRRwXEu6dw9T3q3g9PQOm2azMKn+LZIA4m5SgFyi
y+vvadiZZYexDZNGOUDua4CWBLJnOzbIjbxM9VDHF0vS/+MvlyF2q7ZVeMaNQEZz
KITESMJACMm8CvEuVmG7oJzi/BtxWgAGLR1LVVtCPWgTz6TEoezJmtQu43Wrt8Zt
af9qYAi784axbxVNkvJ9D/ncjS4aMvAABN8zk7KYUwjxVxM4ByffPbna9TuXRgN0
I8wLFdVg5CUNLTI6dStTJ4nbLK0ch0sjbV6RTF//HSw/rqX7dRbo6gmGL0J9qoGv
wt8PIZ25Fqx3PZRqQB4jyd7hPGqlw1aZTD+pQdsZy/w/sb6DKQpNsrNSVSzfarjt
4y9estJWrreSJoiL83Kll0xcttDLiNIupUVCE093JYVQ00/unn4cgNuOqsTE+esF
ieAQOqAF3MVSfrcAVd3qFzwJU+0xppbOv+g+yj9cy816avQcbtRlU5YX3BMk7rk0
PM4/cq7GxDEqIJUM2B3FK1xVFDh5NLN81Q1vyX2NYlEdJeULnmqBPETGhiyFDyJt
Ve1ZBJHKBKSTUcWMfmu7xEG+kg3lyU0jgLFZnIcvbOgmlxAd06db2e/NTFWZ8h0x
tVUpSFh9bItEtgYe94/HLsUBUmJUL3guXGxOMjFj28/q3FrYFxqG7puq8u00ZDRR
Et1ISfZiZP0Eq8S1Yv+WR15VYZyXyi0RVQleog0lGQ85guo1ZJFgcRMomnbj7L1Z
OLmXSxEKDzNwc5NoNXoodGHuE5F3mJ9mszzaX+27rhfQlBimzXYjbLGX8fEy0LLW
G1oFjcn4y6PCAwege3DA0D3K+1/ywqAcovr+whBDwnUlr9MI+fVZgc7yYZPGPf2I
aOeoF1hB/o35zU1njnFO7cZynewoPjnZvljBkXhmLu/hF2gRVWZOc6cZMf2THsv3
VFnVP0d7KhHOu8H4SGufoNBOL/5s0jX01VffnQN7KcReasFbDONh0no0OD0m7DiV
x70PLAJEnGkL/Es7nYuyr9oYf7r6cbl9jCXpTsgdy8x/pPdPD3abk3aO8/ydJ0Vj
P+7fC5/sChnD/qdNI3zme89QA32TzlxiKuAb0xBLrMT7mwYw0eyy+TNc8C9bCget
DpiHR8UsLt23mfg9el6IFNsn1E0yi8+N9ZBaeIJ8bJcO85j+GnPEoPVXCas4Ac6W
r2eyCUWyiqLO0A6Kdx8U56QT0kQxVvBQI78RTFdiM3CeKjmkWlJ58Phl8rpTXN9R
ZEq5lDh7AIF3BfhTFnq3V4h+4EQ9+0eLYR44FBB5VTcX/nZvg2m9//DaUEpIMfNB
hhhTPkhl6s+J5Twj5XdytBp0yCsr8evUSfexvakz+1Cqd6WwAT9bEnFrYut4vGuG
XPxiN4kLx4mzMZ+jwD+zj3ZXGwrJj0epSVX+9Htwv8Zy6TToFL9yE2JC9Mc80Pud
QftXuzjNdYjd6x4cBNRs2aFbYqEirG6Lnm+14eOlHNzVHxPI4PJtXZS+Rl2HGfnk
NFOJLZ6xR97OCUuVilW/fqumZI3vnSdvFL1+7wbWAVmZMxF1AAfqiSXyACX4OW8V
hbE05wIbooF4neukbEqYo6nvtKFuqnGCuiL9XFN4HDZ+mRmpQ/n6GqaNSSv3k7YV
82T5qkuNVaHBJF32y9HlRNPXX8GB7dabR2CkdSm1Dfl3a33sg7PNhVPtftlPyYIL
JJkQDuOzRPOW9x9oJMvSWQfbdpnAB/xA2Ww5umDRHQqnEP3wO7JVHbmbAuSLm6ey
sEWNUtOghOMVU7tnClx23NPh1fyvRw5nEAE92C9b3jv3h8fB58Anld8KI3UvPOGT
+2gaS5pOnhZ2U3MK1QDgV+0G5UnQ9yULxSvBkmSNLfrzBLCjOfpjXPF8cdsIddsH
rV0fgRU0IzgY/dgUsHiH3TY6xPcCykil2EMfvQMmfk8EhlmZO4QYdz/q3OKqVIvL
gkOE5+GRVtqeqLIvj757XQ6ECpSVTdVekFbpdl90gDoKL59JubDBlav3ivuLW45d
sah1uPHyTgvw7oNxAaDAEjNvCKw12G1XuJiQIIpdPkGUQfdz5qo0JQIe+DOsiUJr
4esK5DSO0KbQpVRGtxT7sl5PceKe80VQDQr9pxAgpPEEqF6L4t3Hdc4HOp0Ffm26
uenopNPIKQiIRXFhjuvHp4kHDniE7P2Q9kocbd01V0/rDyq97eC+ChNfugkSuz2r
5hYVPUSwXQtnXeEzR+GmMxE8nY0glJqjg42IWHVqSS3unq3iZYx7uoebMwBh6tVu
Mfp+TGdBBEiyd8vxb9wZt0Nkv6mO65gYq6oGSDHJAUZUkXlUPemsyJ9XUqlaNlOx
yYy4HSvzOxN4/et1pUlhvNSDtFCc09sk3s+2WpIeGecP8kyI7ldp/mH71Cayksu+
+yGov7FXpG+8ri4BMFZCdE0HvtE47PkhaDQO2DCvScpp1aGqqozRAn5rxZ1/lE4g
VmAjvwgu8UnoEFnldvqmF2QpuUmRUjD/c9ciY/WpHVxQFPMXIZQ1GzSmAmnNtksQ
qsK9Y5rAe8W7+AictnlquGj8iXpjJzApnsMmSynaqQi2mYWYxFXAOtBnun+5Wjsl
bNFcujpa4D6UmFENf/aQ0CEsu6W0HvH8LWnopxGmGWo5Rwh0YUYsKSlpqOYTZ4St
i8OtYXRaCM5ayndZmHZJcrWUV+ldKIgacj4n78qyQAsnJjVmVv66Hus3dwxHh2Bs
uS0kwWiVPD5Coz6gyB0cbUU2m2jOU4n0qDa/njegoS0WeUTAbznG75c1AcdUPphY
VtYk8vdSxC4uiXluARsq2XlpO0qWMHbHWlS7wFEkAk7CAc6dpzNVb9jSzzeVpAU4
Gx3LMTFZ9h9VAYl/0FCvUZPYPk9i9E0xcBTVn17k94P51kehfE0NzOvbRddbCEvf
KsQWdwVRV8W0ZckZSmjR0Pg4Krkza1dkZpuHKyLMFt27xiTXyWprrKjzKO+cIAGq
2ENA9ZT9Eq0NOi0b2oyd/duS0933QkT9En2/i3PVimr2QntOzM4FPfH3QS7EuxnW
4uGrA1kfGJ9SvNfARlY+h6BgnyakO7m3v/R2L5L7SBYhzousCqrR16F8rRORZg1T
TQ11cWyPHZHpyFeAq/CSbHFI6QJGSilpfra91eY8xG+PW9GHcCugh+t/zXDSo7mc
XS9YcZuJumEE99kdOD51RR1EGyioAd77CstZROYILstmbRJqkpVD6Fc33xGPK4dJ
qWLJeUjvcf5x5p7l79HyVzz7gAztRJXrBYyNs0avr5GH+5e5T1yggGEKilYSBRYX
YyBwhjo5Z+ic9bOjHbjn0spGNWK29XcYI9oIG7WOjMnTFRLn5EX6FGMhb+E1fTXk
AQRE84xC5/2QXtrYfwCXQ/jvobjCPNke34uhTjTRJM6ZTKwvn7rhnG6JDtNXPoBI
kRZAwOxwRAMoHvJlaFfbKqZ21iofOqcduljjUv1M1iyOe3OXu483OjIbn3sDH1Zs
bZFMOYkOMw/7Xtb8mXjQkCUH6GUoi0dFNL3UnaPCqYLJZHoVPiXvdjfMb8rSaVM6
TDNDHdiEmsrzPZPevikLBgISWZ/TrOHrEoDv3lIzVLshayNENGqljBeULjTwYe79
/QPPKRyropiq48P1mgD93/4bFLG2MR/kEzfzQ0/76aFUGvVjr75JgNaUFpl3gTau
9MWP1ahA+Uz/+Q8IJhQsvGdyu07a1wr9VKo7kbhe9QET94pRiZtEHbda+iWx4Dpo
ZDja0A4kkpSJfTIo172xgws6WOM5eJFORBIUilO+oLEGqK2mElG3HdKaI/28aumI
0Lm8ovKaFgrKT+PMuI1ZRWa4+eU5MgtC47Mcqbr+7KR+wpcHwOKk3+2mWKsazW5M
G7qF+kpSS3s+gg7WFU3RyZTrFamrlcMJBv/lDALOfNaP6pchPlgaXLNj0FrgK01X
9FHNs1LTNkR8wYQTxyFJwitnDekS3tUl/QYQxAo7+XbAq5ff1UplNg3QYelW31dc
VUDsaSpueJEbHFHrnifMpcHxgORdJ7mVlFWNTcsEzKvZKqYOCjmLE+uicktl6eL3
U0LgZFQ/8WqhxCsotaU1LsM4u83qdRXSKe4maKVtWryh0XF1/S+5velZOLkTqUen
x6d7Fx/rSfTJpHE4ppygaHIjE+k8RcjWxBh7JVXsk0Bn4TA+kztZOb8UTQw4GNBg
4Qa5BaJ0yQfOWWG8FBqHt0JiDOlwgjfanzy+bOdsLuowKmhhmt5mtqT6HeeYlsiG
53ItunT1M7OCI5RHXGL0fOmROuMiyIadbKScUNwYXXv15l3cQ7BGsbeD8bVNE7Uz
c30vV/lHQYErTjWdQlwDKHJ/SrzoRZLhYhJbQXm8VtWZeLqY6lS8Q9z77T1td+dc
z/sg/zq+68Z4rmUJTko3buo5SoKkfwVz80oyNm2d0zURzHD8Zptt5Tqow/1+pEKS
3hQlfETms47AfMdXblo3h6+jqnSijUcKaTBqFVTdKYFd4xo+HArROqE9DWdzibkA
NOvcRzTZEDQ5Mm2Lr+TNUH5KXqhrq1jmhOo/2KlsKaiqgbkgymmwQNa5DFo/U1xX
IFhRd4+hubJRKADr6TigRY1RrGWGeG18SFwz5iApM1d2H6ir90bnNd6dLweiPB4P
dRhY7ZqFROg/0LtGogTdpm3VyB+LHKaFClZp/8fI2akrRPhnuVeE/3aaBtAGNPOZ
8gpuJe18d3caeUBqZ6bQvocoRyr3YgcmhLXEZVIThV16adtD2M3qFUJLkaTcA+qt
HA9l8uJHbUISNR9SeSRnQvhlHucEXAfDfKtqWmJwm13YGQTVsvzFlqDkONiNZnmH
iwcsb0hTbsfbBBV9xLKPmnHlb0wdXx6CeasmysuOkbUVAYLhAzvJm6QB1IR17pTL
j+3XvnHsIHDjGa2g+ex0mkjV+jQWVLO5Yp/Lcq4rfR25Z8+JBEcD7dxtGOSLVcgi
y6BuePGCHc2oyAzNS3Jr9cB0bOlwg40qhejAdc6I3KR7Zzw+5tXpriSML2n3vL8Z
t8OZBs3ZnDYvn8T+yJF5McP0gGMS35H8nkK04EdLWXHdTde2jhvy3U82G/c0Hiyk
oVbo32RsXlSeqX7znBQpoF2bVWW2Q1A2lU2Eynj7sfQGq50qnKpIzgmioGNZmqKU
HF1hl/OiVd5/MCGRi3H4OThPgBCuPB4sNuP6Pzxj1PA=
`pragma protect end_protected
