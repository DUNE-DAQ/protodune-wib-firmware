// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WF+kh6ZZ7sJPDuXliXBgWbs+YSAxmJvlBrvfAG+vLjNDw0EkiQ5c6q8Opwi2gciz
7XcKPJ1aaYQRpSOOLIje3FGXmlxpSOFgDlfQ1I8FrCcIBZlxI/GnB9iUWbyyRcJ6
bWqQONhCa1GGmLvBqEg+j/0E2HOZKIZZmhyZmz6/HuQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 123920)
mGmQw/EkDM9GFl8g8Nk3pOdW+biU+qLZwkO9Mqx5naJCIeqrnWddnIOTSKtma0/3
wpcfZnILc5Wq+8t5Qvz7XQ1+044FZhvSXyjHbVQKyfzpDSmrxZOw+G25dtGWqjTj
HQUChJk9ZdCqox+ucG3gyo4sAk3apvwmD3pmNHac3pjFccI3PNOLwGjIZ52m/L2R
1eCglxHkhdmu7jZF1ydTxjDgeBm/dK8+6GBMtN+IdLKC0jksK/iBMFf47VPliC49
ivcLIQ/P1uwmJ55YhvcjycK5tzeweyy9wkEdm3yOBZStfMSQk5kCh9W0KzQXMVwc
uH334WeBzGTFFSFEfHoN1QGgHhnmkk1D3kbYtZBej0182Wid1AeJ9MJykE001DHz
MHFqwiRw9aiWUYOBZisGZy3uvPgqvACS1CTK1ztMcbeSRw2lh89gPbNZ+ggXNxMl
8z+QzWlZu5fqxvou/Ep9O7sHbqBTeofItpWhaO1vKqaV1u/lyPgqqBhw5hldOAB9
k1/UHiX/ThPeXy+frVV1oW3VRUORIcuEN0QdhvHrBEVnk1Cxrb9L/YzyomEhEDX3
MsJRDHqbxz7796pfjuQdjWDvX1+SV17BFhM0MXq4euWWTb0r/uHzDOBWTEm8pYx7
tqD4PJ4aYRUp3tPkl6ODf/jqXHFu+uVYlPQemRjEUt8E9SguOrX9EPg5PDkEYZIm
U11okiKr9dzuDpsZ/zz52tYyEPUnIwAUnIWXk2493oUo91BWc4Ge+ZZ5cV9eBNzX
Esb3SqdRyFKSVLU+xaECQnvXYsJSFiZ0SuHbSxJJhcrWU7CwbkskG+aLOnYpwGPl
v8HW3BLwfeccrL3gtuCzUWpm7PNB6EwnNcrYgNkEMmGdAQI7Up8g6LEuBmqn55EU
5+i6lxCdDhjK97o6DvHU0AMAHX1yqIqS4LzR02o4ds4C4KVWKsN1HNIBOMmPkc+P
KVsBzaXVSLhnb0jLlz2s7BlJlgT3NJSseNCu7pOJoAEvxDDfz2V5xCBUbOQ9PXQ5
g9NFdGvT3TbwblPhn8aYrZIFgpKpuD4598BOd8u4zGqMj4HLAty3iWHgsWhk8o4E
7RIZs4HoZyX3C6QhGUK8jZnR26UeRc/aLd8lEP/diTq+fIAgOIWWKk83adEPphNE
MgTkcu5baV+xw6bDbCmkfb5BdG4PgXuQYVrd29UJiyS5taHU35SyfF+zgmm19lyN
Bzy5Hd8EYf/n2PnKOIKxF8UKor+mLDbLEgRRocp2J8rYDv+/s5++d2GL/7KL8kHJ
hhd1QUNxEiZ/c3yP5tMP+jNofzDeh0xtv1xJDTITKsP8xs7pJfTLJIR3giAxvZk6
y2hozmPlboDjATe1vnd99Cs3mGclJT+7tSIWDGLN7svftD/f64okDaHk6cByju8g
M37JpyH26j9Lio5G2YkNnD+nOMzRvMTE8FS8cI9s8rofN5FGUFoMhog1t++2uxLz
3EhT+xwTGg8L/w9i/0y3pmSFPA+Gd6myZKVhLC7wnefytLUO0Q9fS2bwKacM5365
l8m4AoY7D6Dzap/EHvBY6slrHlnN0YoM9z/dVR9ktssc912PCd+VPgEmEDrB3NBf
T4fEQ/Hryut/LCXKxNde3lUlmIPcria4TsJkfaTGJmkDHZ8WjD4oPDcwyxi94dK+
5232SSan8CT2akLtWr/hYH4txcZe6p41rK3U8ATD96vR9oGUi/GQv6ORta0mcZkL
e1QB126Ds99x+rVXb9/p+OzFWGVaNWHdac/EP/tVw1yxMOAMSUl6K2xOXIV0pARL
oRt0vXXj8tz0AJEM8OoRTNYWB47mO+i0OYZKUr6SoFYUcwwhWOZyHzVFU9WXCOjE
KiypP/f+tvaPjn48SHpeCOogLlevJMCkajdCFzWWkJIxxa1k3O/iK6lpNFbQncK+
AXfPjOxD+WVYk5r0iKUIMo3BYrOVifG9TEl36sXVS+F4lBdy90eC6goeTNSyJs6l
oKP0y7b09d8pUCTBT1mNnGqUqzcFd8PMb03QPVagSKwwYXjTFh8/7sHl2fSZ79q3
2z10fLYJUab6oh7O7/HcUNN4XLIIIo8fnDDrESTqmCZpriX9nlqf9wiYj6N4hY0C
xPCAjazGxJVdBK0ARCnGcJ3Mm5OsUEnU1OAjg4sghAEOxB5wA12dI0IRERFqDP+f
fD3dW9/qNRp+Hl3taZZ4GkAsfRCQeHi6iZV4ZgLI4AbILT1N7URvgkNKY7C06/yC
rsZD+EMI7BhPH+/wnNCSU4Lpg8zEo6RI00YdrD26f5dY12gebj5vn6J3Rl1X4oFp
RuJ5edPo1ZSZrGuHwe802lAGnwX1NVAn2NzKDB3YM8MZDQUc2Gy/lluLVUFelcO+
VOIbEN5deCXLro7ukSOJeFaM/AeDjFzTtLuEPTOCWzBa6t0mNSK+gtWzWbXu/WH3
ZodCh7L7vdQWdfOrqMpDm4EBZQ37hO/T2uZnF3j3Qj5ELVrxPvDmdVbngqfcws/8
LMPdBYNgNdagdCaRNhbux6+zsZ+19Xtygz5olRc9mLD/BnRIbuvc/Fsg+C9lB8w8
HcyL8uJB2KjBDFLq1UIh8tJXq+W+N3MSobowBVRXVAOfCO922hY7+p8D60ojDI8U
bMSlViS7P5ra5PgDh1ooRf01bXN7vde7c7/9IM8GJM1nkaT7RE+XJYWGBeAUYcO5
MBHT1+FDSfBEQE686hxESfGc5eVun40pwwz3HUckfXW2JbI/NAJ2dbPGNZMxvzrj
b+F2PH8Qqx/RutlQ1ejLI0LtuI1nUPgJh+mEw49eipDT8YcY1O4IPE7Qe9/mUhsw
nDB7yndVrHXX3vDBsvB3OFp9en9lMfVVTv9rZSd9bJP+MCQiEs0l7KiyLARcu2JW
YV+EpxTVTiKbhvYHM2ueQ3Qx1EY9eX//xIveVvD5aUcXB1k7qtt3ucT70BtiGqWt
IuVZIfrefPx0pcHiW1GV/BIprBiRatuOlXUTFHwqPuHoIoYN/oXmQ93qy8xGjDmH
aBvOsFg+xH/QQb2Gz3lGEEcny2YKgP1Gy1ErwvTOK5cy0BSZFhvIitJMR1C+3LLA
oj3X+lXPclWo0DzZMojyzXNUcfeiQTp2/A6kKrxr7IvUaaUp4aSSoy28GT8ZT28L
Avo1v2Ld3S+RxfGlfdaz55QRret4DjdQmPHE84QpAiJa0EjemAdrXWOjKJoqJhoW
gJ88inf8I1HzlUbNSJ45Tu3DRAz4kFkiM/i8NMVmIFjifvy54FFJ1nDh4sPxa2YI
6SKzdMBIzN0m9ONn2knIS7EyHbgvE5xz9CdwZElJ0OYGUVrb+l155L1/loip1Be3
hOB3nkuwnfJSbVRcItVMr3qw0iqOM9kLI6TmD8An3VkF3JuqczZT7Xwd1OUjt8wO
8OVIbZF7IxA6m0SbrilX6MgiUY5oxW8eKWArnCGzc94YME8oJygmZLPrE65xAZiR
ioBOZ/R3iy4EECDYF5utmIQJeEqKVmxpuJSq5xcgfMZNRr53njU+fnX1DSRfJJ5v
KxaKwQIHzdnUlWcMXFLh4MWSs6YeCO12xELej5O02VCGN9kbPUcLYH6lQYCniR4/
nM5mtSAMcS9utxKLrUEY5nbjtd5RZarJ/ZZYk8eskyM4fbKip3x2HF2v1SIuNA2q
TKr7wy2km0aApHlaPj5qwwounxHkrOJnzjz0XnGyAZxO/sHnP0ChXgPXnPzy9QuC
/nM+mZ7lCxXPJTFrMpOVH2H77XQsP/CLqAKbC08x1CGgfRf9A44wWlA56X4HCdfd
mhJH08Je0R+vnMPi1kmzU2/VqqqiipBpFXIBHVm9jeKuoY4hmQ2HXITJ9RnEpK7j
u7U+mizCqQ89Wjnh3GUQz2bNARwrYN35CFZ936U0VxAj+sMUMBKjjUnDb7tyOe+1
ycuCwJS6WAdd0Is4lBX+CmHYudpDFhyjbTLIYaEim69ezi/KpRewW3UBWjfordzw
GrFiUiuGSJ/K0MbmijfHOlNhK5+UEhsu+oeFHe5EvMU1gtqhpLE11oNz/bys+5HG
8kD3T01ILB8Zd68QCJASHLV+X0miOfTGJFhqHbGPbGFPcYDVap4TVxkY9d6I91ah
P7DpudeOSZRjbDcW079OVxFQ564etRMA/GNsFKHdg0lR71QI5RFRTb3FC9rJDxTF
5lrlCjMp7xnUKoT/OkH53nGgeB+R8ZI2wMfie97jIbctawKfazItrpc9/hqH8+Bq
qnWo5slDjOMWldPs3m+Q+BYiLbEf1nO4mTLraCK6m1ONU7jmJU9w12xuKH+hilMU
p5xDUEpSMwZO5x8GQHwTtDx0JPp1zvBOxg2fTWlgR4lTn598lBwuOECEVHF4Jb9q
cf3N8Yt8FXFUYCnZUA6CISaaNGLSpDEdiMt2gI+UnVRtevQONs0u5Y/PfDgdpmht
paB0FDEwLW3a/bu4F0HRfg2dn240CcjXmrIMIfZD96p951Pjv6a67Btu34y8fYjB
IosUuG+gLj+y35+W24g7OrS3zqxvri4LMoYz3zmnQUrgi7GCBomv8ECwSb89KH1X
orGOgA13qSAGPYyCiOb2tgHuBcwQTZ4XzitXOpVooUkqK/ZC1TLLhFR1+IHHuB74
/LsaV4mKSYjq7AgWLxp34eyyt+ZfmQFpDHExced/enKt/KuVB/wbP8YJoST8kbG9
3R1/9z9ezFJWF3R6k10p3MRXWFa/nC3bxLybl9DxAEE/8BCWnzBdjidVwVbgDR5o
IC+i17k7rOgamF/BkNdZAY2ZWZVGOVGJK4+9EHQSQOb9hFN8ZjgD5hRSgNOQi8eQ
YjNHPaeFgjlMGMYKDgypnvir04+vU1M8LaJVjc2TxiFTI+jFtXHZtpDz43fBu1UG
Uqq4J+MvQ/F1xivY6Te7OKm7JHZJcGH/XeM5/y8ZjTRtBQWogVohjLuHspWyen13
mqkhixVq68ooCbQakOpozC6TBKT3EaBmRSWWhGF2ggCg1UuBGHNvGacWOtssahxM
UtYVJN0EeY3ajZo2lI3UT/CPmG3oVyViRP6ffdXf0xAL2dY4w3btwGt1EihLxJVc
tSzKF+Z3xWbISvwmJJBQlpRPDFvkusBj0rxKZFjlxkQWReqVkHdb3Y8ihSuqgV/f
bArcJeBhkxGrGnURv4edyOael3o546EwBVsTNrnPOaGJkdNJt/5FkNRgrefXln8S
p3yFa/iKhEiCcQsYWkWcQ1WIYIbFEJR/fSH5MZuLOyLb4GB4jDPk2bWFIHKErRnN
DUkLc3pSbXRdeGdCtImhgcHB6ETaodGzjrJLyNlfYdjAbr9zmPkSg648hL4+ay0j
2MXNWVvyaxwm9yvUniOkQmzX1xPG33x1XCfJfCvYDFdFZfMYbR+nPZUVgr3RVCrJ
YF9UGMeyIvmGOZbfI6m7dK7kfGAAedeeIcuIMoJWqvMGa6mObBAc4zLwzk/Dlx9W
XX6IZTFD2JYFeSZluWyUh2WCksgRVtMxNfG2mH91DwtvdaBplh4QSxePykoeIs+3
L5FYdaz85DcIN4y9ZE780h04X+v4i9pd3CHpXE1/JeekXBPYoseP8SdR/VBdB2sz
Mla6iVgc26qoWtufTB3olSG7AoPspKS3z+GfcI4YHRQXXVEXj/CXwffKebwgkgCn
q4TTCjkjPmOZZdMiPJWWTJQ9VAw+npgravTnAEXG8dIiW9htUkTfDxLep/bGwNNL
b/ul23uLm3Ca8TpNlVk6yI4C9Z5MxPwvrXESH4OjbzIlvKUXv6z1DNJv9lGNSotz
ys7EJT8lUk9ss45KPqAvGt48LD34rrpN5Y3majkZW+0QjuGXxCXG86P+DLFwYPhs
FxH61v1J01rVw0IJr/Kx5ENeJC5uLTAYazzeY7LVdSVjh+CI26gSzvY1E7qUa2r1
pbRoT8ID+34mH3eBMoHLcwzAO0xvnJHjqMhExaaMpa6kNCoPWq+VK4QnMZsvIV3Y
Ot/ksqV5e5kaTMhU8FZnIK3HRYrJrlP6G+aI9XTQJFvmSYtPrk90qMAA+wjmqqOq
eLS77vTYc56KOvD+vm4PR9zGgMqwTJnTrnN/iDHqrGCw5uKlb6X2g22HB6K9XPTu
oiTqrJvnaUjVqgL8CZ5WWdQQyGqc1Dlg6DAWvCoev3s/aWg5e+9YRyte9bg6PVAE
xWDiTswuL8pBISxghDIyAv6F4Il+SKDET4HR7V0OWbcAWE8TuSjL9t8ZB9bGYhtL
goMbXjL3KD1AuSpM7QC6APxU7e24YoBc1+KEU/SNqFWjp8lGIXuhshr/CXluHCxU
ZUCZi/nat8WxfgOOvOrnF0nSRUY/G1c9r05X7UGbyw+7NjkWsZtm6F6TlfKJZzha
iaBGT3+lkKSyPmmrszgY//jNNSK+Cf7XV4QzoQqrYT58nPa8l4oa+2K/+c0S7mkt
A/AMWHC4K8YyhPcBbzB8kQBWcxDZmXGh17pdvsuL4jL1QbNw17EjFJ9T7t2/brTs
ITaoL7+uU6Id3FlMPCCIy/ibsKmaj1dOTn+zveHbyPqMu9J1oHXnZgryiPvXZsAV
55g1IhRr4fLRp632keyzc+iIXImrHpzkpzZdZXb2BnuzvAwpfc6svWztD+PQVyX0
KOhu+waMZ2dQLOX0fUCiu6k047hm7z6xi68RL5td+jsSw2WnyXuwi9+B4ME/BT2i
FmIlINZjDj8UhxZOqwLys+EAi+3Uh/Jgtl2P7rydm6iNMS4w7YxF12y/4ai9XvrM
iLVuuCRTY1hE5ZOq5yvE8yJ1hJk2UGHPiGuEH/UGFSWN8XZIiVQwPcBPRCCXBVXN
JayHcGXUpkGEAAOzbY2hggPajRqyeG9kiQydTOOYAKU0VLHLSI/cSJ1qp7wUrWEZ
4ISzI5dAYnQyQwIofG+yJQOTmIkJpZCWFSDGDHAYaJJro+cSCNuJcKUgubHt/51I
c760OhkfXny/UtJXdmrCYMEu7PT1YDPX9VKA7o6U4EckkEuQriB8MMdFDj1CG427
ssNwPX48PQdEvgcpsQomDqwBO/zN50jim6FOYavJIFigpR/K1tn0yGjoo7QxX03s
jOl0l1qIKEq8ZKc9j52zNYLdnCQGX/lT8pnVmmXb1vmJC+fxczfgC4xJKJZJ1B1i
4JbgrKf6QudL2EfuyaQx6MFrcIPKYa6UgihE0thFOCnv70JRGZo17GswW60eo3EW
oTxZZmJ2BkNzBZeMWMktcOl/fvYGYFmC6l12iIQs4g3sCiIR+4kLoCSFhoXOA8E+
w2/fwZcwKAfI8N2+YFjPxCyIWMwIDwN+bplIXhmKBKBlsYYMITM3MOVPUAa1C11Z
xFvQ79iTyZ0RW1sOQ7MNADMDe/MWfra86kTm/c/frrX99AgnDb/vetC9OXUUIkam
jbj7/a7nrhpmj+stq43h1oDvhs8kspOillKo21BN1gYznl6v0Jcy4kNwwZVWw3UW
Q2SvCQNNHJKgOQE86mVscqe6vvQDFy2xPtl0DpXPT7T6zjHUE6EN7LIZY9NoS0RR
7u0paehR5JWohHrltsFb1h64C+2awLlF2anwG3cVvN3jdyHVAX9Lm3/kTKxYo99C
L3S/DyPnVr1HE4ThM20O283rtf7S9WdjC0G/H6Z8gSlzdpXJMb+FvBE9tMbjUOYh
P/xu/bqb55Xdxx57foaUm541VF0P23HAM9cejySu6P/O9tgsGSw3wm71AXbbY2J0
ihJGFMivKogzNrodcTM4q467iKnlbS2G6ErLgNdme1XE99SNZz6JiYkHLqvPDfSo
aiM/6LFBjIlYQaEZyRYIR8Z9PahEZZosJMHrH+jOtk+WuOvCKaaUJKRjO1dSojpP
fuTA1BdPnAq7r87HULocPPoDek0ewZ/cPw7TEegnag+xhtd1WJxwHN2754WEKPVz
ijH/yn3aH4xs+npsOSaSFnxra6pevR6De/9MoRQFyB5dUDd0EnoeIx7n/kxPPuf+
jDn7aeE42V0RvZV36quvaOqCs8e+kFJt2zLNWvTakS3J5iaWm97slbmgS6z4huh2
N6LgeZ1Ok5CxAHUjtCcIDBB813tQ387kU5eKRpZbFG7xsY4ks580Kc+Kak58f8dS
aQa1Jbag7oj8xlsmoEFjjsuaj74naE1iavSTTUfIWsP94SJ86D1nihzqy1IiEHAG
0DvwGONKK2spVrM8vBA15ORbI6I91PDlt0w0C2Kyyw9Nyw/kafRpibVkFgHaVOWD
oiwVo9moshipHt3gakOJ5/QuAJxMjYoreFxFXEFQEgj5MLNBabpxFELW42i8bpX9
7Uj9N4lBnhnlRnlQmWfpcefk0kcaMFPybuiJyJrbUIaVqZccjIssE/aMCSZlSu1S
tWzmWAe7rKaccGE+U092hM2S4haD1VEZ0Vy/DUyxcBXD65N/6xRdslCtIwN6PUoh
AnQ8WtCkSOtLRpQTEvoJJkAwv3HpDiaMBmqnYv1zKmhLAQL7LSjH/hDQN66UHdJh
4uovvW0U0b7rUI00UhY6CEpyn7v9yZ8RC5Fh7wASKNGMAmcMerupJujsBiuQiPGF
bj4nOVNQoz6STwTFrasi/16SaJkb7Z1wUQRt3nqUMeoEntY4E5ILaXvU4bGMDr3l
vbXaNvwILCsuP5sTIJB8HZtF5sf/aY6xcg9pJDEbA4I+wSTbs22q9JQxtwgpgeMU
bkTIMd9OKm+apGcMWLbpZ0zvgIO8Hd8GTbGvd3U92xTnlcZ9YgM9AwZCxzlS4TZH
YCCNiM3b/yP9wetSTjvvOhEsIGtIAYmgr1BE4ZtoCmVaeVB+RKwVUfMjC7HdPH+b
EnNDWxH0AqcUpE3uZFBh7l6E/6VdZYmvsh0O8JT9IQPsss2qWSdaZmiB3u4yXLK8
wCHhrpCN95o2SNA+l59ySdfIpV5j6IVNbYZIrf3D2SwTIgrXqj80DC8iR/4uI/yK
XumYDsqcEjJaLsCPMLthJYZWydjsexPTqZXyYse70pd8ShdISe8wy4upLfzztgNj
ubZJk4osTgvJtgfBcytdL3C1MjXsWCj468ot35I0WjbNJXdbZ5HmtcsIvgDc1hVd
UUYa7zk7sOFHjxfWp3dB6pDiEnX/6xL6lTo00NhyPl3jUCH/aAXlR/i8x5/8UGSq
FfoQXxib0P6x2JclUmYiBEWcPz/RBzoT9zx6lby99zP6+D6KwLWhTjF+gm3ZrEDe
EMT7jmF+EZnXvVxoPU5vtk0Kg00XtYJKXK9NeI/SM0MbqtRLLzwkVod9rGPooxmZ
VfHbNTo7ZpCfhGcQkVilTXrPz7lMrOvwCRWT61THrEQZLRdQfyiGJvBt3wmuya7E
VIpe+Hz33rVS2KJhwKCIsL8WtGW0UqsGaYlUerNNfALrHzKagkDVvF+thr8mvCbg
PjJPIsaObsbEi0RXKmG7WJ+4gYKOP19Op4hGmNCE7C3kd5PEterIULv/AUy30Iak
YNgmBUo2D2bUG9sJyt9+IbikqHtDaJHeNatCbtAHEW5hQc5dlQhsmqzHeqqP/plW
V5giAX6YT2ZtmPxYlBMa8Xa9TcF55i+YxttTXdqTn7Rg1IwnsLYeRVHDUHu/jH6l
JZ8HIDwzhouPYWSmVdHZCd5tWqU8QeVaUGrYxIElWxT7euQYBMVscvsxId4qlhSl
U5qL1+H+KSA98fB0wwvD2U9yxPr4V+Zr253+7/t9S8peimqD/1YeGvx1Dt4xa2Fq
sEOcMJ3rKYk+gBhI4VazSsmuPQ2NO274PjE4Cl9NBckGz+f1egNs0NawvEw2K8my
RI5EYyJ6O0kR/OJ87wp/EPZh3fZSLn3xhhtIClymDPLFvHklCeF7d53b0qTfuruN
h/GZLnT37+aoP/YIlSMdO8N+FdhYy8SJh8kyy/dQAdTy2u+29udmZUitliPmpmSB
Ztd5J1PbwDOFLgnprsH3LI9kpy120vFh8sfNnh0iQqFlp8KzC+ical1oSCq1vfX4
c5JOTA0vH3WQPxtQJ9jLg1NdBXU6yeTm69Uo+8wt19/2WgoLQBX1esFhBT80Cu0n
SYJi7kHBNTAtpUjBMK0us6ZVTqUqFJOMaPe85cZ3p3GVIfdAArEMuK2e6tDqnB2H
a5JRvbkrTiVcEg4tO5H3nv48ZMQUC08dIRSKV3jLxHlDUmmAvRasxEHyQhs4tj8l
H/2jvx2qMQrCfrOzWLqjBPX5QSpglneC78wRTDas6UWAx3nY/YJ4G8GqINYLeuIr
BxrS+yYiKu6sQZ969KKfYsaoRP6QpMGIf7ScCHDyUdN4vfsu3Q81p5L72ThhRK/G
TMHIiT43pHK3umz6so9OuJbuCbH4wfuAoZOtxvv+mexaCXZt3GZV2N+xft784LbC
oovB2U/y4Ky8aZKyJ2Aye8a0Z3K2gfZwnZ9m03QF+fOtR6J6qcjts18X5GtACAa+
kViCWh5rYcjedMpv4/AJRMMOTauG6qVQenTQGowASC29ciPSZrWmGxN0TKrO3I1W
VjfXBCNiGJYln4aokrFABFbPvLOTxSO5Jn4nZphz4ne8hyrv/C/wnkgOhFOwWwdJ
8yo2/+ON010l+DBbKNoBdPwVsWvuB3khYk4JOh+DcI3Kfnok4Z6B1l+UZEvL8D3U
BekOanTT95H8ez0cHP8ws4gH7rWmZnV5Ws/OzHLHN2al28roCYcBSKM3ib/4uQYT
wTqJ/NGy+6lVWnvSVS4t7Kx5sGtSrwMHFfwMmiouJkWRJhmDtBeolWl+h85ksy/f
IMHOD48kOLDCA7eMppsCosF77VKRIRaDs/cOc3MYaJXG5tS7+dw7bm225dHcW7C4
KfjD+M/eGF2lQS56IpM79flqUXiXOckdXcKkbimPR3z2WMwW2sHGHsZvnfPck4Om
2Zjy/cTEDk0bmUKvWalwQ/TtNYsXl8CVDV7pX60pLZa5hmVRn89krPsHsKHf2YBo
Ar//HibwaAca7LR5vYJCLeeOjzfYqqBA4lzIL7VOeZyFQenUxK+Xfe0dzOGeyCxI
mnfmRI4PscjKTLbHl4xXIOwrU6d9ouC+6MZ7qCKb42AVafzriPyF5FaL2jjKiWxV
6iXG2gbOL1XWkq6tuFVMd01rciix/SS0jXkxXXe4ylq6NJnJJ9rn4QafPOI3FxUv
T2pwYEyeEalDOQ2UEaNTrnAzW2ml7ayN1WtNSkQqv/bsUlwHHJilGtdSNlApJZ5i
Ba4koK/aeSzwhQzP7IjIDW2NZuT6sPJ2sJ60wB2fTWnDnOGiDem7OtrCt1e88yUy
B4HNKxffgAnUGyDIhuDdx+jd/+54dua/+xhOGEmgx05bJhVJ5cWzJ+omw5Md6df3
jrfCzZwWK109v1OvJ5RlXftq5gz7mRUwFwRzF7uyoY75U23oh/9Okqhi8fHAC0Pb
nMStITa9Ew4B+RMF3X9v/HgO2JkZ8sxthvNq3pbpkR56FqNsnZhOTCtTq38QKzdf
IOMOOXYF0LBu91vom97Q4xbAVd0mD0DR10AJHpvMuhfubX2HRAwEJD+4lHoQ5V30
e12tY4b45FLI8XX/3jDOJxy9S1tvICXhwWsDtmNTC+gLwg8kWqdICtNIlWwcaHsL
6elHqyidUKxbuP6hCjYsuOV0VuhfhCF4lq7dIv0SFNbPyH19xmN7H5+sxAUO4vM1
RxoTI1IlftSvBWbP8MU2BnTeO1vQMgYRs/RCUbuySRqUQZaQ8t0ueTt6TGaowuho
av1jUUkMBCJ/++WQ9nXbu5Co4cGrzxWhcO2HGQBi1xs14uc7KRKhatbVRoFGCB55
sM47ItGoMu6JSFrgVCScJjoETPnrNbKm5AVvsLlwQt7VdvO0D6a/+4oxvvDuhiyP
y2DsqIGuzcJFDXaqDB4uWbYpexAtGVsWYFlhpaE4if0DZPMKbh6ZGaWJ1KpRPkK5
4nb7OMx9sRpf0TyJUIjuutrnwf3DvvG6YnM/aFTcKj6r4HPwnglQ8jfwsGhTxcZ7
vZD94MBfrjHbgINPhAGJQD0e0wlcGtVmfiTW81NYj47gx9tmLMd56lMoDfIp17Gu
mr4pFnpSYUdVxYIypVPZ9n38KwuOuK1P732frEAmrzORqVCtOZFe8Q4j+5wPNFcE
K18PrY7msYL76f1CiNWbfgqu/4UZw3ohuKgV6O7KPPkvRI8xx+62nMA4OyJjk6u/
pXYuBgbkQRcCVUPByAu4sDkX1Zik/pc41+50lzneRB9uFBdpR+gOXHdei1Gx+Aq+
MRxyMWfA9B6fcGhKWJGANgocU8mzbKrzLtCj2NgFPrPtQav0XyvHxwvwU+yaY0/9
H4zE4f3fT3W8nNObzmIEkHmAe10/gLGHIEPkJOzzQZ+t0V8rDscjQhomR+21ptB9
6RyRKwCk8epfCbkGka2bioYsWG2rOEuXRfmUqJn9LX/gBxHjqQF+HhBfLnp9I0Es
86e8McIq8F7KxQG7SHa2sbK15lneKGBGjkBwWnO9huj1ZL36Tyk57hlBoRMcKLHl
O8PmykIdzY5YvVLaTGkstimJBqdkRiZArCyZsGCM4f2ip1Famyl9ZDx7IWDb3/Ul
diYwQZy/+PJDnJo4melXktBkdhTN3F/pax5x67lori1Aoz07OITDpfuC+GDy6VSv
7lb/lFch9VWhqd6Ek930vPX0qgxmFbiOfD9MphAos3X/lFzpirpaIOiHVqFYodbs
of6/+KFjc/JpXf0kghmSUPUxJMTHADLEC252MgN7dLTp5pNMkjAjqpnDDfvD6SZZ
JutGxElbW0VJRuftfOX0rGI1Puzer6C1d+C6M1STLYlSCp/VZOdCqJh0Sbtd6Mwa
7nFe2um8UDTRE/nlm6ngy81uKCRY/9JxfKqkEqGQUrasg9yMvFFqgNjpmBZ7ZJmq
VEfqMl/y6qHkhs0ioPW2pxs7kxmQ8p8TfOE8Pl7PX0kjAmr4TfG2O1ltd8tEuk2k
VOq6TnTF9Yn2MOpEPlgHQps+2Rv9DZhf+KpieaYiePsDdXMYYF8iHDlj1IYgUdxn
k1q0iiZBMB9TbZsGRWT0xy+R9oP0wL2wwwC9ncH3jtmkQ1XAwh4iBVCmimklsxsg
SHAt0pRFM2BfEpV2YCkVko6v+P7cXTmuho39BwMqYw77ujPEHJquV/cn8/hs2ryj
GY7RZIKeyD/GnTBjlwSeFeibsUdWpPH/xV+NHvk2TwLKawU+491r985TMi226uWH
0RjDhTT/Qzgt71QRPKB//yO4rUDxFFAbpKsfv1IMUJZeNHNrTPqy9TzD16Svwvnk
C5/5DgJUilfoHp3afFSylL35dyxPaqL/NKB6i5zblHUD8TOGtiApkWO+u+rvLJK/
93iYmMKxXhuIGTgKLyzp7+lr0dZj9jDNtXKBAAxNHwcm9koxSZxeC3jAVscfa9Xr
axCBTw1DpT0LkmxgQofV5eGti0UgVU1qbYymQhqpAfrb/oG3V9tlQGGUyZCplxrA
ggz1NmoXO9e4tPgeI8gQUUXtDqEwIkita1YqSZcz6GOm5hv/NmTYjS2MYiJSx9LV
urB2yP7I1YJDeMz/Xh+eFZaUIVcmRugJ0VCtSYU7uco0A61kp7uUvnELw5kgb/5L
Dcb73VqxejtRiHrrU75gdDwkYOjI4gnXj4ldGMEmVlPhtLtYTOKDDfOpTbWswLsw
CpVwoAm2hf7BmfZrKnJBROdT79MzxO9lcKyjGeoWicEh+XIjPna2VG5UGFJ+Mfsg
6WBBnCJIcIPIVs8zGCCqNueuGybQ8vbUuCu1gM9nnbuqreIXy9GyjjeCmXUwAauW
LSLkLlRrlzJFvnJ4bEu7FdMPysQgIJt2NdHct2rGXDaBmal7QlTfGpiYQeT28M1g
HfX8Ch69naK9bMtK3xKsKlbI0LEaENb5X25EdQqBYY8QqEmGYTT8XGgDmekJ2rcN
ZVUbSkXixiQ4HWCNfk4zp4Q5dhkP45MkJ7VrzxgclLC/mzptikxDeMpjZrCfCf8p
FYg0C4KrozvKczt7UtgFR8HGl03PAm+7ZhUPj3NfOrolaPvK8PG9aslFKSvFbt2H
u5k79fqi/CIn3CKTOH1S3EkhaiD6HG3Oz/Lhf0MR4TCQluiWvXK1+8WjsfEjOIM7
jT1wuRAyLSWAsjEcS3WbTAGKq3VYsPQhgn45dhjvC3tFK4OJoN+n5JzseFgfd2Cu
tmkAlmV09XjyOx1BCCn/jFsqVu2yWlpppPVeRC9ZgEb4oCwF+kcufRc8t5cKqOCa
kD8cnRH6cZbRzSJCVoPWCqhgCxlR5XoIO087WaQg1s/575PXa61YBj7e3chReOl6
sn9hl02Ob8TeUWtTOWo79iwQ79QMrQsefH6uzi/DBSud+RP0iPuiR/LdRoVrgUbv
IH6iF37M293VOXhIrHcukURYbxAVIC6JNCLKzFdLFAlSKB0b2O9fS/Avi3Q6iMmG
h+e0Z8rzvd2jCzcND7/aeC/HrvOvSeAbKe6DLDeWgbfl2bsDbjxhXFxNou/glhX5
S1u0YEvOVE5GvNYEcUtdXotqqPDSD+LyRu+1vSdQFTECkoaUNHigxCkX1jFVGlJv
/mAW3rUSnR594TjwrQ67GGce56pKY9gvTgULEHtmCJ/aAq7GC9vwlI6g1vBC7BB5
885LBuTuYwANIzvFh21MaitCT9bE0vD3kviCVE05kx5yF/aznD9d9mbGsWycXD4c
006lpJgKreBFooHeML0Pjeib1WEugzVvOb17omHO5ZCVZPT6eOC/QRb0tBgDfS/W
OVjpnxeNTxTdFSMOsyh5WSjesYBbTErN82uNQv33zPAOLMs9p/ko1/wO5U20SJpf
IHhqtU7msBVdowViXLnP9BynT+KGisOxv+iF+LTejnSF2yqHQOx/BKWQSJhacG7m
cchV2dQsf77mpLCwMwi28nIeJ8u75XzBGRX+rIJjUvqKeuWMLtcJAQ5OkVXBY5q5
3x7aDBvMleCb3KJdEm6CBgEOlAsSX+HzHe4+BxIhsa+zdwU3EiIOlzpxbrbjmUz3
qC3oXmifQvPYLtofJ7qlQtvVnhiq5LFBddO3rnjs34Sr8zlF5adu08onG7ysRvRn
1WeXwxTVPJqB1OreZ5ONPJvfgFlkw8e/D6PdnFkTd+9qCTLv8y8XLi8RrvqrON6p
u2TkRwYifGnIcrCXjDQSvS8lD18o6WQb0udZ6VlbkHI+Abj2ug7SHCY5T+zV4KIV
TpB0FCk5OXQMQpQ/d7tDcVhGQ788qitV8p5cRYBy5fTIXMGI45hSR6KP8ga7OJjw
mVOI6dlbsbQ9tqGuVWRMc1PAoxGQiWGMA4hwZQHCo2iBqhsGEfNcspVW/1cCH5l3
f8RZfLXymM+xSyo5Vt6W0gYgF+B8oDU7UiX2chJNabUpyeY1hvy3e/KQ6apg/jBv
2fBvYM3alpY76M/hGTCtw/ASTOhWVSfQapnEuN8oy+uBJRv3TnELeY5DYJut7LCP
uhCnrVi+MzbP/Fe/KITFUT/6zq4FbQxjUQCV4XW81XK5nNnFpzKqQzcxUoW4z3+v
41V0wga2wnOLIfKNpjKV/zZEuVveUwzU1NoAQlktmbDC5DhqnH1Q94APty3Smmyl
NMLfhu79iQ8Rr4rhVy/LGzrLMXCWcg6Z9Kq7oFWD3TE8jp1KgShRmJssX7zpp+Dl
cVLnux8LdyixD4uWXWU/bPT3JTdXApvomA4YkynJXKRfahJj4rhVQSFQP1BjcvjD
WOQtZeI8fN+q9XQoaAxp44dRQgY/2ab8qeeA1ggZlBx4L2wq+KqP1LOAAc8YDh8i
guAIkAThZ+Lf2C+A8BDWQ4YL0MV+JhbpAnhlDkGF5Aytqq7QdrWt4Ofhd004Xp5O
bnMQZrZN1Zaz2ryGX6ORc59ic4/aEmSxqLjPK4AxIk0sy6rvPVxZ0sn3ZPskONyW
ho8wvlwIDtihoDLWnPHyU5pzNViLP0lPIaiBO130Tj103geieO36lu36l3LeEhpu
JaD1l1Sk9FFw51il6mqF5DYFLc/rpCMkVgTaiIgFVQ5gEqwgll3dL2W+jSqS2JTN
aZ2CWSW/zEEAmw+fENrXA8UIBw6roa0kJJOGBaGbnjqyhWB1SPUnIO+ve2A75mnX
enwHewAAeYR1r+meAXJAr3MbTePTP1sU0IooDLFnTT9SQKQLaMspjgWL+2xk7IF8
yJWSflc+rJg+DVpACJcIb7LRyZhREqZQ+1acHS34H3iurD/jurZyLfKOvytp6y9u
BJud+F4J9MstQPPEzCNgSHU6Ssp9xkcHXeitgtLubEyG38Vj/KO3zhA7wkbwMbzX
gtbIAwosrbBr8O7m3FwVtcMemyXjACUY39HzNGj0Npbt3bNChvID4ToFvyKARmM5
BEjZuVX7Y9/+0pIIz8JhTSTL7dTP4aYNBhM/xx4u1TAvwZ2jb0KxUJK4pD4TJhdE
kQ3troVrreth7v5avNPF8tGni3QBvWDRGSIWUwM2q/4bP1l66HvxgcKHnlvhMtaJ
eiCCvI2OIkWhPRBzEVpqb/4NBlmHfjEu7l7i8AEhnwqMbwETpI+gbBT+kxhYb975
JdQHidZ8veFSkV52opa6BDnpci8NXg2uT2ys+1YrPXwOd6FbGlYzGZ5pBCcEtLXN
ECuFl8opShT4AUrsjpOsqTHgLB1hqnBHp9HJBEjdqBG3DhQfSuJ/XAVbmipGSsrT
aWEdwAFFhqn6Ns9eBtMfzF60VucGfaa442+G2df00WvAFtk59dYn+9nvYvfWtCZR
6HH753hjdTl8kxYGir8ntFIr/k0C2bkWa1pUnfUklt2LLbWndEBXZByXWQo73fhz
wurbiKjUh4Jsq1oKYzS/sUJi1PPLWcY4SH/IbIjQ9tRLMfbi8ss/HSBVcdsaJiT9
RkRUvXMk7pOVpRSYcjF7QBaJN0ffBRuhuyMpz3V6TlB+U3IsAg0Y1lf1KGNpnYcr
akEmG2sQUnUVfDiE1EaAkWNEAx/HW+kycd5PEAlxrxn6Z5QnnCaulBX7Sf74vqkf
o8p864m4+TYNH4Str35m/sxQLpQQIyVPjA1L33piRCtan4go5qSTSRRNTAtuLPLK
WGuxgWhgCrQwUMI5Al9vCQ5OZ0vP/3vEJmd9b9aSZhrY5sqwZJHnsOSWIyHISCiX
Acnh4NKiQM3/+VbFxNzEoC8YhHoIjto1dF1s8rG2W9tUJSHSNMJZL17tN+RF3xf5
cImQQKFip4UxiKGlr1ciZfgIkko/d/oDl4Ubcij42UIDJbCaa7NOfNshbJBswtiS
SQ+QafVxzbOivwcy+LgvzAQjFcHIRPtO4CykQqF9WdpFt1Wf5Zz9eXYThs/oHH2W
vMO4PM6iVkWAzA77nEC2esQ5zwpr8IKRty0h3tsWX9AXgzaTj/Z3EyzGsCqZYp1z
ORZRlH7kvCXDr2mHJLsMbS+WvDonUIS/Ttu6GLgSCCLK2VvrkR6dnz9fWu7jZ6d+
cIzyvcOdT9cuOz0vzcjWUKJQv3u1AhEWXbJKhFGp7mqDolXnpBzuQp4BsW28OdCV
wFtLsC2eqrxdfD+mZGN7/k9vUY5sYMKMCp4YZtvnBqJN/lndLR/OCCbKFFW6dCgt
Cr/EqZuHH4F8LDG9ohMBIC981RCKnt+dcd9HqfxCjX3uOTRuEI1jKrlkaTo4G9+x
JHbon6J873qsSEy5plV34OAOyCzgV3E84uRW5qTJ0h2Gsc/qrGRMS41Cd+7tP4g7
+rZTrQ7PzqMfwUFurzfAvcVjQeqwtkxtxITDgUINw8PNzQ7QtfQetCavky7sTR8b
sV9W/c1za24NZHlGe9mp9zkbEyBw7J9AQgUV+XXpS0+3395TUHFE4E0cAoCDCA4X
8SSqSpQFYbXaNldicpIAJ/kGci+/8PKf2Lf6eGRlPOUHtecapuWmvt9eEjhxYRC3
xvka2c84hR1ex0PoJMcxwJ9RKMi2x/IklW4XeieiuLMcIvF0NAtT+Zq/hUpztPSw
GS1h+iM6dFRiQtesUoQuiY/HDxu07enHQ5/vPXdOIvDcdO1YtvOIU0IAHMNETpqa
4cB6DGacBD0wjge8YKf1oPriPEI08J7lOmKycCGpgzJAqMQugoCVL4PEiKNrdBX6
V70s1ogql1F64d0erVW8gNXDhhNENBDyMmWggdgbRJ0mI0ADpe/KYGdBUbM56Z7a
iL+4qUQ50QraR+s87JD6744cePZaMl+H0c2SwtM/KjOkquxXleR3dXyCxapYlqyz
JgOBwS9fJx/FAdTgT3fZHJwU44194HdVF99moO618x+fvAndG9vmg3z8Lt/exRvY
vL1yN5AENcxEhNh4rYiJvhUKUEjf6Wlkap+tByNRUlYFuqwstTmFy4Lrg4cQMqCz
IxaCgjw2mJm7ea3/93dq25qZVweabpUJWVqZwXWKPdPjRHi4Ptzr2iWzFlUtTyQT
fmbLbiNUIA2HC2DKh4lyCFQZiEtQ6hN6QWENnINd3PJoTTd30sXwgsUW9D0sVCT6
8/gAFqZVPuWp9yVDTlqHw3dbnThKO/wxnX8qFUk/ogZvz/bG5gF24jpV8UvychZo
s8BBmiaQ3Axg0x2R5ZQNtbwX3hnKTd5WUNwRyGTbmcAGpS3uUfLNJvWFqrqINeBn
d5s3iJo96i1lNzcnMBjf7JN/EHK375aNwNXBdtpxSF+0aSjqimxgGmL6KLuoUOwG
YPluEOgp+Ql/LWtzwzG9cd77dwpDYBg22x2+XdXpSUQP0KW/7tQv4l//LnAFjOpH
3poqfolACTC/WyOo67xcCP6NLLBA+5Ij8EZmcpZTDXl8uZyaQBBvLNX1nxPPSRfJ
yoBvaCWxqL5pGMADcWw9W0Jvbxg1fuJPe4RK1b8we/DyzJ76H8nfMT/gCMyU+kq9
VZPZfSZtQ8EYVGY+rRLbeBsKOWuDZ4c9aRGpPWFhTuX9qqYmNuN0JCRrtBx27ItT
YLV6siG1ND1alQeq1t4bb3vilGYsqw5M5QhlBuAFQSkXmfX5fQb6xiizJZyivYAV
uRO1csnKMvZLIuuD77eeLarOj6VguLh49wjg0pXa2ImYeQCt50JcEbgL9B6FHzXM
QFTgPlb0gww+w5JY2AC6iYBBpS8B5cW8+F0sv+wAI2Jr6dP/PLGkVhtkbROSqq49
W/BcEziClqMW/ALGj2lzIlZ7htV3wbvqxtOShXWz56Ph2uwAGg4tBAQYFdzB6Bu8
TpugdUZll/OWBiasxm6gxEZDV00/z5dshDaIoV6F17bAGWk+cN9aIPKGTgSG5DrK
DhN++e+s8rvPi300pNtZSp03kpjgvIdUbtdZGuqxVI1zIbHXptgHp9Jzw2uaEGhY
CYamVm0TNDdvYdo5Q6R9JuxTGT+6E3spkEFljMydi0OVJKQhfSHg4trTGevvTyrG
80806uvhJGb/L0a5aZr1td+ih0yZ+6r65aA+x8B2tTAnhhlj6EYOIextkmkYw3Cd
55H7CZTo0OKvvSEZIO/bTEWXOPcW54T71CNjOcwFoec3C/p158FvgbrzFXZFirAT
7U80DYh+opD2AocH+NoIf+Au5hxzxXsMevaaR+GLo34Y/5zwExmaXGhiU1TFz8kZ
bmpWPhaWF0/x0Ob8db0yj6hvUq0u954JQiPPLmwM33kQAzx5pHO6vVMuKS507LjD
lbIu9R1e3whI35F7Rc/0MKaBW7zkHVa5F0+nohKZvdqUMCqDINwRKus6MwgdCZTT
NgQE6J7L1V40REYFutqJbO1/J9+TxmvePpftOe8+4UbGMvMDO4LKG6LpLjPA9uBE
evB4NqRzrKMQMnowMO1ptxQrSl6SAnFQISzeSppF1N3QhubQMTouVbSXhOKRI15J
Lst1wLoRBltYnQa/Dn+egVST2+xX5Dbc85qvwMVrPCG8gecURnsQviDyifjG/6+P
0lmBJaXUuu8BNddIw52FGmDtbNhSnvIWRo67MUGsH0ANCHUoL8uFeVfSn/YKNpcs
8tbbhvYeGlkUL2TErHE/h9vzLBpvp6LcH/EWCQY9CRPW7eathLJAevOqNg0atve7
uHCfI4dWwhtlQbz2+5iweJhZdeaGomh+lK3wtSyRAdsNNwIX1tkSIRvVO4jhSoyb
qAls1Jjb2OWvgzW6kYSguNFWWQaOJJ8vehNpAHriSHtZbsVe3sbBIuBfJeXgplBb
o5ugYbyyMu+bk4RQrNysz0BL4vOMOMl9ANEGF3RKEUvusWuZ5GZZHirVrL4svHlJ
Hs705DbcuNX+6Aj4URg9puT/bsA2SmXGyk+Wu4sB2SMaL3jXO2k9ewciQOSmAGIK
zZ5NXl0wuGdVctGzgPc0Z3Y6nUnV3vnhU+rrrz3MDL37jUXScnpdkQN4ku5JitcY
QBg+Ax5WgqqzwbLhi5DDpuhU10C5nHBxRVBdpmCsiWGqM2zWL9ARSgGlNFNnJqOK
xA2HI8rqUNRJwr1pV4jLgCTRf34jW/0YSMuEhOxj/XlV07ji8o8bwld8D8vrRhXI
demGfcuF6uXnMXwrCLjl7CO9o2RSISXyW9fmJCdAmSlNd+sRtYIRGwWFAlLd5I6n
Y5OunUppNpwAdvPBK6Do0tlkc1vaDGYnceurb4PKGnC7tJ/2G047a66TrTHOqTmb
WojR0ZfZDecEp8GnP3tEt7Is8NCbcjst0s4VnJNt7nZbDvTOIfEmRxnfKppME3Tc
OIB0XoRvBqg10x+QSTK9i1BUylfbClp5QTHTATAihgVpgT5PB2M7eZ5uJV9z07y4
hnd/n7N0KerRgwJLCtLwLtM49+0Wl2zn5Jgxw0zEXWvSJD2BRRwM3XkOvlys3NVh
T1BoKWJqsmmuyF8klRU7Z4eyaai8mE1HB0NxbAvTEeeIp/Zn1RblkC10N2NIcTOQ
ABQaC5dGwS9cy1qtvluo7qeMGyTkXK2e5Uioc7iG7ArDy/VNgvi729tzucCt5kw8
uaGLXJatveov5PuVpTBGbdszXybOHmSSdod+vgjclDKtovD/oHI9Wd2VECoPwk/V
80R2Th+7A2CfHjvAcDq/TjzQqwihDFMrwHBaSI/jZE5Kv5qLTrv3hIoKzXjdZtD4
oTQq56Hkt142YIV0Y1wOfifq+6cXVpJCqHusWdbl/jEOPkuUyCVVEf+AWiohPuGi
lDKufwe3KJiR1TLSvdT/6wX8wtQGf/F4nvu13AluX3eRwCWxf/qllidYI2ylUmcQ
gMOK8wLlUM29hTbMyhnxf/QdoPDGEbu5d9CFxIsqXEZ00YSNLsMc5td6eDGPauhG
8++MIF/rLOSAzHl+Ab+9/K/0mIC1JMhyER3n6OPH79rz+1wIE4jSW73YGk83EJVe
fZ8kAYClP5iZC/YzeM4CjX3MracZaTVhCJ0hgNKQzlVyhgqqkBoDsArmbXeWXoDU
L0L8BWzmNnbrCFT180ES3toAcMXT5PoENwU3amB4aUGJGHYez9kxYKd7yX/JR+4y
snJ0xSzbJtilePC7c725Zs9bAN++bHlzUO+LSHRadoKPLb+QXeWtbCL7X1nIHBnw
Fbui/loRcX9NX8FoEXRFI9Ox8m+3R1n6MIiVDgNnxd8V1ULRB+HGofR/DNMc3qqV
bjeZ6s/AmT5g6u/Xp5bNHk9ahWc7LKKuFDOBJ206WKlzchYV9AwOkNQu5m0shwWI
7gWrwdOOjXJ+NtWxKDz7TXyj3ez6tmLbPuzIYXQ5Kqvr2qRHiT0YahEGkrd0pQxf
Hz4CabYgiM5JWI5gqS6Io7KZae/z9mVZMM2JclOeCKz5FbBvEhPfxcgCvbzkfcxK
UjuMAPAC+ZzbRkwEq16Xa9uFYdPqHfpKOakSq8WwOfcGBI3ZPPJ9YjbJlKFIW/tB
1KNix1q1IVTWvHzMF2SBg1lAniBTvO68dlv3cs3+3Qw5+Arr577oiVRykKmiDYfd
+I6gr1rutZdvlcz8XttcObE4+tkYylo+zQelALT0IPbPwmhqQPZ9j0lrWHeCYWNz
RQ0ZjAIsWT0cpy/ZptiE0UEBV4abG3FpJ2rWzxqM3nVIH6G8CEsxm/vGyiLzfEsX
9hubzsdsrOB8jXTeYHFIcBX8Am6k7xDzEj3qbkqhSaWBIGHwDWEy+qIFsRoduZK6
60xbddiDKVF19JaKo7E/qIwyzym9V8mpxp0qiLY+UNnO8s48IieT7B+2127lPCE6
yhkwvIe4mLpNDFHz36Z+7IQIzZWfYb0s5Cf63rxz0VxjMN8rbib/1oWKhVlwBvt3
Ow6kl5jp2TvdrRFl5FlA0w8HWyJ+3mWofZVu87X0LImyHZlBAgzXSByRBf84CEF6
GRjTwS4Xyu5KXpbpEtKecP3VORfbVdrdSYFa0l3yfYxaNxF3/f8Or5KQQatMeeCJ
tn0j9bMUueAazgkHSCiXKizxk08mF+RRpPjUCL1+9Ga5nFJCEg5fiU51hZqV46o1
4gl+tprmGQPTOWfbgeWi8iAoKmKdBfkM028vhawn3pmU2/HVjjMapqP2cHfNi+OW
pHGB46l5rISO1RtifL+loAezE4w/+Rxz2QqWu46D5yc/xoSIr/th8IlaKhwE0gdT
5KGLYacpg7X28eRuSkzE/jbZh7I1hTqV5lbu6dIZKEa9XDawqCdHpgZoojDuRx4d
40jaX1aYX/Bjdiy8vycAmY5QOhZ3K72+LTqkNk2+WEUf8FuuDSsYYwYREz1PYnbb
lIcdl4Vkcndbwdykdxtc4OnKHsqnMw1kAcf1J6Lb6WUGze8RgaFgfHw4daNxrnkJ
2i9dd2h3RRT+iVhKU/G+tqq5mzHICzdWrXtjX+MfRv+Lr14ef7izSyP0QfxMpk3C
535nt24aQrr8AUIS844HY/AMhAwUkdkk0q9YjXWswBox8/7r1zYtAf9C+d2VwEb+
2KnGn377SpsuGBdXTMCXnXy2WvHdQe7EzWTHAbErRl8qQtE99nVGXmXL8Yz/BSv1
3rhn3zgsIgMX3+Q3/ByVDgKcroOaVCELWtYc0hH2kzL4INpoxfXyRBDL8i+nGlqm
qBbH7p0awCa+8DcOTCbVMY/W3/0xakChmKD4O+8yPzqCa7dBxt+yzbdm+J7s0Bnf
7epXzsZvmopVSFgOagzdAKtKow7TzygIwJoaZL8J++Z3iDmljNPlrjVkXH6TQHRl
zRM3YbZ6ZKs+5iZqHVYtqCQdMK4UnO6WsR9uYZL7JkV8p/ikzuhqVpJAR2XQsiMt
zJF1ShalQGhaqUCIsQbL39Evv9ifhVys8ZpS0m/MT7oXETRWSi0c2YbT8gyNlhHi
CNJmEEaRYYgJZlCIkmcVKws3oOAFrlgX0BxNfnKp2sMMNzX10a7+H80vTTB/Oi5R
N17RN6Z8mdc/Tv5difI081a6q+h5NrTpf/N1KULDR42G3Zskkwx8wgdfAT5ucMbN
8aSaWTEyb59xx5Ao+os2DLOhUJdCnmGTJ55Kc1RERCZLEUSczS1RMWbhw2B2a9KA
nzxuw7rWUIhMQseufg18uMryTL7IILvkqFFZgBiAXBrN+q3LVG/8M3znOhjQjcMz
JcawSbzKOe1McoH5/lNp9RRVI2bRh5oIhErLqOlkfPaHspRKFAP6jWDO7BsFZmzB
tMRJWO/+l6uKXQ+raxnv/KePiMVEwOg/RLMqvOGuOae04Yj0O9HnztuBOOWeOJXW
aIEyEJqGjUuuA+GyjxVya6Et++nKjqDxdsGAXfQqVrYl2oh+GJ8NVvTll+f+6uzR
xfinL0jEax9P7Tb6Eb2FwE0pzruggbhjG4lbIh2CcfViRLr+bmMlp4edYN5FW9Hi
KYlwPXgQA7V5YzTkJ184ZPfJYmd4VWHymI+Bklj3qmQ4Kh+RqQ7SchBm0Py6AwXm
Agx+4ZIq7t1jEpM9Eu/Ef/5pEDrF8Tqtw8h9QdAeZJ7ymtgEkE5RU8i0S3NDk3Qw
VmIUE/irkb6draHEJ5lUfhWb7f7wJSR6jT66ZbZuPL+ift/+VNs5lJnKXkmQdAB1
QM6Ct0OCxQXd/qvJrrM9s1fuRE/FJ9C3YtIQOelr3SgXi6PInikhLWNmyyyptzFH
v4jeTF5E0eVBci39nUJ3RNe3hrvxZlt/u0kKvXc+EUAiSTEnp4QazzgfnrPbrPwC
yKubbACSqx3/+Q40IYouwqp+757G/RYbNH90d4ULuxCs6XGohbfimUCws0A5R4uB
iFjnxtVbQPUTxi9z5FYagg+E2rjwcLz6eMDhS2CJDAMPHJi5nFdmwyJj1N8VOGtu
gzut3E5AM10l8foY026uaUM4U82qrhOEprJBg/p1vejMidZEhJWpM/GxVTqvkwUR
1OzvEQrLcb7gI04nOXQE2vM68UZuzZrCJlaQMt5Zj/WyOKY0r/WWEVePiij33chU
NB/659llZsGMGvS5q0Zjrs/L3/LtiAR9rLF+HpoK/dib2m8xTu75N0GhkoJJ+amp
dT7i0Rq1M/FzQqU50ULadBkmBkgoAbqQriXPDl/iP0RK+8aVCBj8LPyw9OR+DB9C
E/4EUqX+F269StUQPLw2swOIfkHkZA4dyzL6NwwOJiEoagK9R3ifrjRI9cFOz+P0
SeuFNZ4wTP55V+XZQZNE1mZsxH76FA6R+yQlVYmEnDQmGMGJBDJQ3m/O22XK8mfi
ciByB4Jfc/sGmQ1+j15o9go7WrLuEHkNHK+vrLy6kJ+bAdwgs/GXA9Vej2ggSh4G
Mt4zh480KNxUqiXTbI8x3bk0dJ45GIKySMqZiH1a7WPT5AdNkHxkNse9YfeZqkjI
ndBf+LjcXfbU7FMEfBytFIbzNbfEGc4JeBjNRlLzun99c4+CvdnmMHKXudUamq19
Ytfvt9xjv7t5wrij7eBY40yEfKpCYUYSrVGjrzDPUXyFVPDBMJUPBIZTlQZUFNG7
cZkPtC3QErXYT7WnqMXR+D7nia1rYmu6Fl07l/YOYrxWszPYXFQjLYjlJHY4CmV7
M8k2X77EyRkNs5l4XVvcTy9faHaIzzc0idhU1Z4imdpTm+Ibkf1vu7m4zNqLA4R9
CZI6Pt+kcC3Ab2nQjuuIwBugNW5i7xt+r9A+TTRLvSS9PT29jNPCojSnIQ4aecDA
QoAO9tMsLHO8llAUfIO4y12gc6wHlWQl161bkBs0Xzdk9sKnwbef+XNMoaC3ZmTJ
UKqT6EHcZ+rRnTvandg6eNBlNyKS8fas4I45ejnxccWqfUEu4Pfn/x84Rrw3cO2W
ob/5QhdNzszvK2NgvXkXKAc/plXPewvxUFgbBBOEHL/LJRYVmt/fMb0BESLE7c/I
f/FAH13zytLg3u+AYUjQUGYBGFfwsIqYJwyamtG0Kyg0kAK0e1sJjZXM50ds25dc
a5UAE1Agsq/oGApZKyVxcuZcf6RfToKg8tcsCFX7QeRKVrLripHLO9bigLzaDuig
T0guds1VUMqxsYi39g23X9+8NVS55PIUSE0ZROG4MzLqSj9axPzYreRw+NOrET7v
7hxP4XHDJKtJek+VVijvp8tpylcI2mr71n6lLRIpIYuPXRqavAnc1KwHR5MU+tEy
0dqx9/cj1ABAJG0E6C7O9rFY1tZCoPlR63VsNtikjPgJsaHwgIJjHA/SWF9sFx31
RZkp3K78InLyGcOL7aybOnqj/oGNK8JZZZDsFVDrDKk9UHwrG83/zh7Oy05sfI+f
Ij/ZJzWhqpSyi2IorFHHb96H1qu7advbFzO1Sz2tG+4clTOUUeBwQzVrEhXSyCB2
n9DEg1IQkkKbvMDDZXITX6EXDOETjqiRuGf7khbBLfTrSv8R+3dFOMjXYEzLgrZG
hZogOtj71uKX5NB5CVQj1ijgbKRWN7Dstixh0bfVSAqJofaJPEisc3dUwjROEaKn
Dr60X8uwhuFZXFCJRfb4/w2gZBgdwfgd8uIxLS6e8n/B7Py9cgQGEkhXEKPGMr+k
r2JXHUdnDZdo1GibDc0GrBs8cPc9YlsPD8le6ggIgMDDKjdBXtFZqGo7IRFyrtPS
Oys3XkmMQFODnk+MA0PwD0MpoS1xHEo8fvHR6P3z5q7FnnPmlSYecewgk/QhmTmh
1W8kOMcruSF+3y+eYZWN6p1pNHhvdcZBALJS9fueauEuoA5kaZcxxgCKxjPJmX8s
fvp16AX4Or+J4V/g4rVnaCcmDol9tuWz+YsHI/GIZCgJuH+UNRD2olSZTn1Td04N
MbqfrqYTzXX0I2oEwwFZzdRbeanmm0lm/eN0i5lZdqkp/HjugPu7zvpgAAsqiebR
FzHHZLjBGA54scHhrdKukp4NgTKYfhMUWldZvlQ/bjU769sIaKGhtrlQVf7D6a6h
nI6M9MKjftTSZi4SUxqMYsmJ6yiIm0VGjCIf3TSXodbEbKWMADlY0MbDkLodsc5Z
WrG+el9+oprR5C1lErLQhyN2HIL+HD9MKo1CQ67YnKxzV5UAcDzEJGqa/09VFRkn
oPtUk5ggnrDb49OiArbExGVrN+5dCQhMadIQw9Yvi/IGom7OhUBPf7cfY7Vetdwz
h0Hbs97Ti6gH2RzNtYdBfHT6k1Ug1UmbokBuV0xqnpk4UQJ5Zz+vNg6sos8lgQ/k
MZJ1tDbDJD5Yy7Orezc/G04ic6KJ1IiuaBFTynYvX+T+E/96Pgg7yBuB/v0VPMQi
aTtZHGdWwEhHyaTytaGcxEj6g34x2OS+dj4MJ9OhjRVL0ZvadoehIVoFtH05IvZ8
T6Zv8beAIvHwAjZrmUxu05pGxzHj8YP6IegFJxTsuzSY3IJX/mKZ8jZpT5HexX+U
0xstoQAkWP7s18zUx5b+0cEuyD4oNJ6yrdOfKjGrjMQ7TcFl321K6/U4Rn5uJZ74
3GeTr8Q8XpB60vxZauvn1pEFEbYT3tYw5IYYkQU3q8E0Ve9ZxZgu2/3k6Gp36ciN
orxxcAyUlGZTWCy33052HKZXp4Cx+1wpjL+Mhg5/pJeu3QrG1PvwOYjHbLu+LL1P
ubLRdvd8k98tXf43jaOzBsZH7vP0uWiOIS0/1sN2GT+q1K96XqSmEmtJ5b9vT/Md
kWt8hp+V/ucOCV86iZPwj9wTYQTjbypKBuBRdh43T5AwX+VMafTiS9bThRSnEwex
He7PMIDAkI0JX1JxFgLaA5whbNp+fT2ysBP5goX9xNZGS0AA8KjwdJ1hZozQPxzE
wxa0pX0sm+4KeQExqBVhuj2KyBnWfopPcRFJ4PW2VVcOY3EPEadaTsknR1hb6WrX
oFllqSlkEzJ8D0sQx+zm8TTOgOdADJNQd57YEJkn1BDKUT7PNzZNVpuKIhW/3BUq
YPeUgjTSU+V/Ccsd03iDWN47wOad7M6F8sQ4JvgjU6sxbWHAh3pZsmmC/mn+Ezyn
Rkix5vOUdZOUE9jfM2+d98J94jdCZ4xXrJR7NNN3a9ZB32pxeLrcTi5a5P/2N109
g6j4SYUEprny+plSHOzNTLgRzCL8bKzOCdvC0t+2HLop8yqHkTQaO6SMA7B+Ne4q
XJDI68i0n2f+M0MKOH4RIJO0r+ZHb9osofLDQtDuGwGEDPkTrwyIE/6CxX86kAkG
X4bfKo4gS2RqozDNe6BRUPGj6aWQbNpUVotYc2B+M9HBfrVY8ILk9rAJ7L6X2TDk
DVw0wArrWoH6NLHvbAcilMXvKP4q/0MpQzQ3ueNWjIoSk+hVivr6X/T0hf2T0k0c
/yKkskt0go0Vu7HvbltT/dvo9F5ccQDPWS1S1YwL7tcK/Br+dgGqoPnxcZ3VZTIE
tyRNG9n6AJytJD69exVn5tGjWMeFUxACs0GyzzedULQP7hzkzo5grPCBRqYbScfY
mSAExxfnMMxG1ouUsuOFaGbtYtSCLmaMzcLn2J1R2tgAEH2GNmy5cdrF13GSNGhW
FO4YAjATSdJS95jzUdcNaZnjjNpkZ2gJCX4oW2a2xa/gQW+aYPYe5qmnKg1wTUQ9
Ebh8O07cgGEOXv6PECTZKoH4uLdC06tlgQcjsqxZpDZHOUtc3tF8gznN7gs9MCxg
kW6MJMtMjJxLsQuwDUDDg4M3qj8ISCOfHoazV0nG72D7CAnZeqwYeVSx12ikuneG
581VlGk4nJhY+a7DxCCL0ovT4xNYQGXYFllgOwSvySOPPcIZm/GrgikmHEehG6eV
dsltLm8d1A76ZdbwlTAQeAsuMiNg558EtPfJuvKlczMWGDrRbpS4eJX8ZCrRaGrU
kag8CVykAAz0UHWhFMqpZXWHaf14e/NVQGqM6oCd47V5E2aPA4bEn5y+cZoatZaT
jbYHth8lQ5UMNrrDLGFtDNDtDYWMlU9NJBu/i9QBqCniobqQ2aufGfDE2e2H/veb
6q7uNHI72wuTKIWl4RUhKFOHAi6CRQhZdiy4MWTV/OvYucpJUQWZFPZIr2KKkkYW
uTh9fQ+txayimEmmB22GVLYE0QETCs8j2i0yj31lZYOB2Wjw8QEZM9guqYsob83C
W2WfKlsVC+QvXq9etQQT73LJ/3yynSQ8Vr7kOOm47sllYx5EwldUFIWOdiHV/nyx
hhbO1FxsfdGvurXAe7ILK996KMlnowhdvyhwVh+u6kdPkFRgcSkcLXFS8Kuj0tLd
AbkcL5RnPBKTxDFiKRLVnsfhgtyUC1tVzolnhoXrDU8pCGIybM2JXGycp3/86QKR
p3dyur5LEyuLq6TAo6AbmQbO2LygF/vJVRWoLYjR63JhUz1o8a33k5vpTBxfzzQX
rIVhtbfq7fFtFKCde/SRyJM1nvt4FU+fUi6C4HyrdlwIm2wrojszZSFXMt62bRbi
RLJ7NkuaY1u53caWmhJM3S51Z8ta+jGTNqFh1jqSDxx3NFf13CVeXowHADgYwhmT
lHVTLjfvhTn3qt12y/fPqHrXwOdS3XUMKfZJZAb7w84e9cFnIrA+E3C9Kwzb6wA5
flgd27AtTY29jMc7b7ACqidSdMC8wwx8R7Th0+WYG+aAl0jAEaUkRCeEDVNmbsmN
6Bfp58KQdJ01DgA8m4t4GyAd4PQ6dQcviG3AGfpZW/YIy+Ry6pG9BUPUOG+iZEPD
gYi9jvmEiMInJG5thQOYzPv+TAO30uQvdkqYXcrXkIz7UYlro8hDFpm44VmR3ys2
Bdc8BLnjMBzJm5sPf58+Lyqpn64sC7CkUgfCcBurlBlYoEBkLRx1qbqaB/Mvwdff
yP+4TVvoX5FGiVXn4czioBuFoDMXGgP1/gmUpBXsenWn1MzD1lxiVySrb6Qm9Rfl
T92iU2jxhcLm73holdrSh6wnLN5Zus+sZkDqoq4T5H9FNgNf36IUqwqB4qkYchdh
OtG3uHvL8lvaeH37D2d/2oV1GdYbeD8Te5aHBqd4HwewTARvQBYK7aPRjndqHV+q
VBB7227uEoVNL2D9KD/0T+oYDmpwYLrMDLEa0zhZshzZwyX526tLTo4+cS8aPX9A
Y6CxlOkOsVPKZK26eFb17gB+Ml3Rc+mVJAtK2whFOh4r2STkWsMsfDOmNOv98M8H
2TrD6BtuR+khJOitkeymBPM34qJ55wnHG6+QzyL5Cs+CdCRZzAvasn6v87qP/vEE
WXTsuUEeaKgNHjDUJcYQsvzMHSa87SBz+M95JXi+WFcsxeuDQlxS+t7z+kPyYCcU
5sXlhfX/k92i42v27+8lilvJcIs4a8+yZWswQoYpJr3vqBB/Krabberne6k9U79d
2BMjSSsKSwHXWxb1+lkN6EaPSLKzQsX0wdE4JFnRV9TcEM8thQ/fl9Y1hiJfu3xs
dpV0PE90YWVvTKzFIo8DBwEIx5HjcXuzcf5hubYPi+Qt+KeExfEew0zS86IzUEew
KyUpUSRSXVztQA6Tr6/jeYxq7BGgiyAIJYuhUkd0RJCtnmjFgSuyYXYCF2K5U3i9
W5IAgZU3d+wPmqFfLtDtYhrD8NyWbFtS3ry7wurwhBkh2i06TvFsTZxt7XKQXjX4
L9SMzUvyXlVK8AvyDQiWOnyLvfLIbQKuQ8vMKCndXPlYy/gFzXAAMV3D5fobStLh
Bt3WOk4C2UST10ZroyiwA9esPUHXMMCe2hMlwTAlP49jopqCAXrqs0SXNL5eqLDv
yI9JDOQStcA3hRre5BjO2/nwMU1OfGDJxkSQh44GcoqeUrSc+s249tYyCCl7bAcf
bhHghxccx8O+rUGQAKhBFaZfxMRYZGz3Rh6xXPsaEcDNhoQx2230ourxQnmhyn76
pTAtzFDD34IsiLgybvhDoHEL7TzRNhX1YMbmH3PRPA89OpTvVDR7KOJoDf5NarLE
ZVVr8m0L7gXh4S7lOu+rdxwyeI0JN3dRR+E9qNNQ9x4lckxcAS4r9IzIvRg2iKdk
MyeuFOaYc8T5R1VokffguzYTyZIr7L++kikjHkJzsT8XKnVR38kmJNtFlmD4oCP/
ZnB/XX1iqyBjc5R9tHll6o1TG0z/3ZSTL63w3waqb5PHK8gBk+Z2AuLuU601FtHc
TvT0JBThjyI+Hg3SpTvkSii7uS+0plKcGNcUvDqzj/fMhyKLNxil7rWGHiAmDjzP
2PBJzpuETl0k+jrEDi/4VKi2JG+QVgsWUvdjbkiwrzkfikSJvspJjDuF5gmiYmYu
RrCONvDnHvAW8UHQnCSgPpHhQ5WBxEX1VwMdXbNA6SrXlfF8Gt9e73SuAuVn/ePf
rYbGkP8Evw43e/12RFnSJ0hdiCyK+FiEbbNQWCr8T+vptgKeHDOgQI3xaum7j7TA
ALjwZ8FNdqFLUoBEWpEdpUYPe+lXo6lZha00N3jVIaH28W2iZ3of2dN4AS8Lede9
XZgZ2+hXSGQQXv96WrhPkuVr0Gp/XvvpGY6PJk92CMZH/SxNiGCSOMqavJCkhgvt
UwnxgMSNVbhb8r9fiQMX4AVeoCwU/X4HSvCJ91bxYC7mTfUY3SckmywY5d7yMTvg
uuip4s2F0Pam5mn8MuzeBQ88MD+YtVYuT3DWIFwxv4iCP7n1ctdR13X4ec43I37l
zzZ5D5cyM5t5UmAyDKK/mj6DMRf+TIDdPk2f9IeZlE54oTG7DLGx+urE/DbpBHpO
9yVxV0Vrw/SfEogeRe2TPI8CHnfkOH08OJDAQQjKLXxpZr2j7RT5djZdPWPa4wpu
83aP1hgD+3QYVju5pg3yfIYf3uHO50XjMDxTG7vdor0PiMSock39V5+yRLAKWpQH
ULUoudXAVocOIiieZUIMdmJ+dkKZEtDbYrjvu7hbDqgN0e7HzqxpFhuLV2QdquaH
+JPdmmxw7cuPv9GZl9mOrIyG+Jv+3eOb1w1XrKjk4ufo4/miIo6X4UzI22anLqIc
RFeZtawiN9W2sUK//m1Hq42+/nCiQUL3/pTsNN3BhJieQX0nEmrYWPmO/UJFaepC
6uLXVM0mUcZEgzdEx1vAvXvN3OIyCcgxi/klhBLdOuR8RjRnEhvd2tqt7whG6AW/
U2wOYqZ6aTtG9t8uOOYuMAQTSGyCfefv1u4G+hl+qIxCJbUSwm3+Jrn27ANiyBdc
7K0V5YTVBP9PdV4VZh0M6YZH0e9HDZLlBssGeol+iRJvUFFq3EPh7ODgtANnklk9
tjpS+FnOzw4rxxdKWJbsZKnek+S15mz1buC64bOqaydL065Cxhr2DuVtnYP6Jjw6
CFkp0rOLyAo9fQNW8PTYquTm5jNI0ydB+sAHq7P1rvyGUHHmxR4TLoXQEc186gI+
zo7R/j51awueYEJYKEuGySemhf5riFiF+WQFId2yYwfijMFSXbFjYswd3MswY8j3
Km9kCQsSBSMAXSYS6haGg73Q7aX7iQBZQF5VxYGmqp/eUduNKW0kilBArYZXQF8K
wI8LzG5cN/MKyuQvDYlHB8H7s1SVLRoXyfOjlXXDpuqwFuAnEEfRxk/tEmEX9JaP
3+d7J87IzlMdYAwvcqZWLTnGtUY6fGqELYiPr/+a+pp1eD7E9/BizjirJcCAUcy7
z3Ai660g+ZC5v/i266P1GcCPQRNtfrMIy93NPirTcAv64w9Fdp/ojjVS3HXFNFYc
sWSsJ2D/7VXbGe2MGu01oCv6CCEgHN1HvgZ4BxzuGvi+D2Do76uqjIlhMzwTwOeP
r6GYAZQYm41YD3M8QW4RcA1sr0PnH7kI4xvwB9XKMLABp72gEIni+aeBzzogVqnL
+y7YhzjZXaRAdYjKzSUw7S41c2ApP8WerO/uAqZrorkOJA6fWoyzNdFm8w28wsmd
AHcgrAD6qLaP1uLMyZq+IWBKvgzZ6FHTXBTAvqrV6swMvJH+aCsJdleJpaVuTwnr
z3ngpGZ1aVfMShSudE7/GGes6kFbWsP4NLI2cY/Z3sFWhd/gnox1MthrQRzc+cfu
LcadJqcO9zs+d/J8wdJuufel5jpZaJ2FOzk04LvK+Be64Q+Gv1jn8WDTQHcQevMZ
HalxxVXXv/PNiSOvupuUo2Sgca6HSE7EDKG1MrVjAOdX3Pkf7yP8cEiB2obSCdzc
6MRhaeroHitFFFrA+8bc0kTXzzbznzFKNqdtDl0KnE2dAVRM2yP+WCf5TiFAWUGI
Ard/qFU4om13qqWorR3EYB5W6u1YUiN8p4aKrVDRJWlqGUqOffEg0Bxg6z++Y2oE
EesD9vZaFKT4T0zEkzEJk0KIn2rRJZHoT0LVmps1yrpfPhAAX11y2B4r/ZhQ291L
iNBJmePPiu5q0nLme5sUfAACBvWWiSto7sYp606JSjVkLPBR+/68iYYFWb5kMWGQ
N92KEqP/JvHitDZFnuFRapIEUVudzmMjkPBaSPOBMbXErStGPHHlZHySa/oWCpKO
e5dock/zIQ/cEtlDJtSFevz/bjxK8E7y5rlTpHH6F443FxLiD1g6R1wiFOoLxRRk
+5gQYVdXJ7MjazmIcwRfcKH6ghJs2L8SqAV3K7lrl2aSzAJGJiHbDtHdRMLtZXwF
QpC/qUcmSV0hdZqMMYQYxjV6/67hS1cYjxS9ffMOWhsMXo7Vm3xf5OmsLyXHCJMB
N3vH7EzN8OywDC6EnTgRBUvuDb6RhCfSnlE3mcjB3PqhGZy9I+rnyddk4xgeGTmh
R5hLFkBNyFXuQvyaAbWfHDGZZXQLEhZB0HBzmNcqhu6YsjHXCV135cuOxGk1wUfP
zhD/jkGG0AU2l0kc6PA9BFByl1gcUzkPdxGGsQaztCVm5ZTBtHDYoN1HNmlhT0l5
/8teYgGWg0AGxQdEydFaJbPpBHU8boMWDMuKmCqpov6y6pAq7v7sZXXutJP7ecm8
I5clO//uuAX//BAjVOLRaQ1ngSe2gsezlZaXTNWzsd+SE0Tnz7BDkcYQmU7GRmRz
a3jo8vmB2fyEEOxlu6D/GVDO1PerXu4veQUFovCFzustOdbjWZe09uYRTcj/Zafg
DbH5OvI+qxISi18IQkbcMLITdYzYE+FSzmpU4u1RlvoE8jVRp1BGKV22Iy+PZH1A
FqOSm6kOIVXXkPGI87x2TSEIcao8q5ghGV/wKOsm7gs3uvRACCR/H2XRfWUInZko
sitIa/HAQ+vAFRynoGsHkfpjQF/9KMZDyF8LucC1M/X3cR7xXaN7Jo86W05hAaGq
w7/1m8ILAecMGcJ2PW3byR9Zz4E6QHGQ1LS6lyPmhQmcGSNIVydGvtrjjOhzfRiS
xvNsEytr4rCM6UogNRlZkKwdpZDZz2WWhDhouJaw5dC/JQnC9eQ+CC1mO6Gr+2af
6l+MV+I77rA5JoAHtM5mWJWyQ/JzkxT7DCtoyLY1rC3t421dA0JiokHVIl6GRKcT
TIZuFtQR9bpjS2tDh5P1ywjlJR5P49po0v9vZZ2yNVst7o8LOefVPuf1TPwesH1L
hP9p0Cqne6BeNTD80hvVjvIoHRohjdSYElPPOHz+S3q0h78X7Kczdh6QelmjJ8ev
i8UkfQaq8+Jbq5v+H4UJST5tszks2Ahu6TrKR/itjCKE8+5XrY4u0OiPkMr6NioY
K8azAdNo9s0m8pyJqLybs4tYUGOdVU0qoqff33hHU6jszCBlY5T12wvGRqZQX1MO
Iqz1UnI5B5ZID4KWsW9fFVi2EzM10dZJitwBPmnuwGzVaDHyUeJ7PEBTEvDQG1ck
bQ2rIb2dL7sQDjzd1pGZv+lIxqRzeTWAPVMQ4QJom65867dhVMD2+oBlDPev/OVu
SqvBuzwKtUEPd3xkTr/+Eaj9YXltBFHm+uRqxOZdbvjWRGN60QVAxyYSuVEssTBT
fCn04fFTp+fPkvzTRKYYNU4w4R5kzx+Arfr23bXDsQI+fZWJcN7rW1jRPXrnjEfl
hsgJnk9NObZBXsK0gk3zcT+28a7B5bVjTRvZRJiQu9LHWGTN8xxMF11g2AHHjN0Y
rpJW6YWYc0dRTg7kcBsEGF+PLm7ute7gLqwv6na8TZ8NQDjWtYv7vEs8qVz/ZXx3
a4EujGTa1FimsbrIpripe+9MVJAHgyNOYGQwoivu2KHQ4920qsz+P3FRER/6cJ+w
mTSQ1J9AjpenXnXCNT7RzICJs5A/WTbTVFr+V1miSixviz2ATKZbE5LLUV8G5Qpd
Y1Vk3iI8GaM3ky8nwKLqu3WR2KETJdopETXLj8pNt5Nc+iYE98y7BKmzMGc1LxRb
WfMOFt98YPJEXIiYSJ9bvtSgTkmUlUrKBlZmYuZP+YEXLwIKBRg65bUnKSu1/cm4
4/wEwLKhRMtB37T8a6y+w7DSNjvEmXKIOu/cqgnsvAZ3xy4haALQ4lhiztmsFANJ
8pXOB9LXXPiHqdQersiTiMEYPabXvwumtTyZOULvtPZYfIjR3FzdI/BspDAhFXD0
bHwedqwp5SdsxiSX8YR50SeCCBPuC11clh+2SHeRTLBllBhCzqDox8OmPaHnAPQW
2IPRL1mBl/aOOFTk+xw7wYEN3sv8SYz138Iwa/Ua8znHdxG4AC6LuHlc1xsFY+UD
cYieLJCBy11sLvGE7xhoTrhpJHekORO4D4HsMZ9H5R7DINnHoH2TMtFLUpQ63vQz
3+HlYtADMWDMhe1ZSnvTyroTX5JzC5NPgYetfjuLQQShaavscBl2EujGyUltSsg3
s8wbxI7w4Cp1rl99v09CHdBnRTvgCvoPIgUPsjjc2mKOcUQeRmGn1GG5zR3RJnmX
DPXE1tNvnWeBRf8MQEoepbxNfs37Ku+3b5hDdwXZm5+7c4RTUCYhXQAG9PpNa+Cv
GCYNOeMPcasylELhmL9O6iHKcLWqVT/lZdmasYrDJgNIbmj81+X/SJhmEPAEa7gc
SrUSPBYoYzqLfi0LwG8hZVqeqmqp/ByVJWSYWGuMqAGVx9J6Df1hNL0vYik169LZ
rb/264qdnUjdRsjqyMQ9F34muE5+SiG4GgRZvAIQSL1CMIKAx+YkoRu8wDYoVnkx
jacf4VH+qKLs580FGIZVjDxCALv1WwejqGjqJwC/Mf+bekUbw/ZHtRzqkB60UUPq
XvQz2PpSM8XdA+1xQNqSLYME1E/N6XyKhrL1xPaivucrM2/RgH1ywsqSu1dQ6Lot
+Du51a3+TLnWiv3iDMOMLszH0ruHbzthhMtefxZFphazkaJ6OdSvcy/a7Bo4aD8D
EfavoIvdDfQ8h/1fTLwzmIO6BshONkB1VSNfj0xvc2qhRYYvgUv2MOgx4TZcOvGq
FDdQxLCrN8J0LKbuIARKhAMAm5ctuQbfrMZL7Sw+arj5PosWt2FEOucWvqPXvlkU
BLiq7/EQsFaBSDXXunYCgycy/MSr9AujCbl1kBHwfqYwdHpPgdFPTdvyYy7rYE7J
lzdD6+XIOlObxki0ZVs7jzCPFD1c0+OyHoL8L0byEPxJirCAOy8QEqk0fzg7VOJI
GJfMtEQcENkbyleNz0SCpkMoBhquZn7YP9FRPMyBLvc2nkbAri33hfd+ElI1dM41
9EkHlxG4HAMiqsLXLMayOE30BcDpAX+DdrBi2T/1KrAjK8tm6gAE2ln09Bn80JjP
FjerR7COJkRYbohi2abeItxhWiq0XIa3RNw4NTlQwZmA8s8Aw8/Hq9mxdk+iRYNN
YAeZUJfCqIeOeD2sWo7d/GsuJ+hvavuWNuPKqFI413MVZD7m1mSirYdtiq/UsEZp
rnkqs7h665JhsqCRRApS9fxwUHcX/CJWJRkE3iY42yi67n71hWrYxOAXZR0hyTjN
YqeT/6aL7b7lIuMeSh+cRe7eZR144Wpz6uImkFvbvgYVlVNATH/OaI3BE2V/iULh
GHVAZsCWW8cdflV+AnDbu5coH4Jusi8Scqa3c7kw95OoNUxvp9vFLxzQTrWuPjph
e3VakcimXuddNVlajsn/f2Er1DrATyv5rod4UTZKeW5BjoeaQZzaYTtiI7I0jZqw
4tIgNtAvUQdEcH+0aANjOSOYZ1tTYSvsFjGQcSrKY0GgUt0RELNFA/2am2ez2xmV
TyXvxrCGPThPaxGFPbDwMBMz68OpKsqJinlpl+WPW5T+AbQ2tmV+8eIW/W3zGM8F
CMzw6hnlSyffcHbmxkEcrIZamMvtwdOJPOfcRkFIine+Ews/q9BxiflKrCVE40jC
yZDRTh1pfAxGKNest8e3fNE0hzSS12TZEetSmveAE/T4U6JFRQ7wr43agc5s12wv
HKEAOwfFxSkrokAwp/MybYvBb/9CON4dj1/gXeDqWttIiJighRW+l4mep+Ykea4X
rLS0OW5JtZdsnEdjqpSFMwEhDL5y8mLgsyhZ0aDdgx14dQWNASxRxQXvI4zDHkiT
UMd7xVksvt5oZ7IFL0ZZ14HgiUH5PHH4ftyXo4VBJOh4w/450+/gZ5/5cVhTHX0M
c3jytvJloN6QpprGxEelRbcK0jeKL58KL8xG3h5/T+rQmOol5FX8MXNFEfd1ntRZ
lOEp+UFfimpPNEWjcRrj0oVsZlVWSD/xiZeS0NLpjEc45+YRK9IjgRQAcb/2PmI4
4KA9f22RvVEza0JS20VpoYh/Z2NZttxx55tMKy66APDNcsk8+aX5YxQ38bib4qLk
WqeCXGcAw2/vtZ+miqnCQlk6Yn6Glci/3vJwyQtICI8YdLuMlqSaBLWasGKUsfkE
MtbMcIVwjNQdk/CsXx0KNgiRgfG1re61d+Wwle3et+weeKqTpCfYgi9L29B3HRrj
F9/S9gK5Wd1q4qdxE03yZRinwzb3qPLF8UK+FWBX/zfyxDgsbEJMzUt6W4ZrAmqv
5NQ3ay2uhHfAqRCODsUeXZkoVXR3uJFv9ll/ys2BLM7bRR0lp3GVoOPy8qQEVP6G
bfOYtyYJPTMM27AFMQkBHPTQiIh7U8cOJszrucvQjRqXFs4AExovnMrDX2H1Tjfr
YL3CyGAo7nURtVfilg4PHcd3NlFZZfYdHeD8wSq/ojSj+G62I/dtXlTk/ZO950X4
CexB6q1U+0Oft7c+JQocqZGPd/iPEfOCsYE1a0HfOh7HPewQkfN+4KpwVjf2g35o
drGhwX4BS8AAZ7K8IJLHSe9Lr2sQM7d1uIGGRjOuHnPgmBZNwzk9Zj0RZs0sTU3x
NRswDojOs6C3OFNaPjGWwZ5FcEwPFjUVyNykHw4UgRB21WxmAWueZiZJr8LbQaFT
PrZtM8IB2y0Blu5op6LL6ugaRuFjBf0u+Thc7pV2CyDc/PQSfhpclGu2HP5Z411x
HgnTJc5FGCCvUOLoWY1lFhmz4z0fAQj/U7etdcToyfqNtwpp9ktkSlaD+091lc+b
1VXp3u4bV/r7e2+8YPLgsgzZY3rVaiwHq9XzXNPod/DUDVpmmxPMP+WAfJJfO0qG
uHB4VfASIQ2CO9xnJdv9Nm/2wYE1iZyFJEuM6Z4BLrjHAM41iX61XqZ8XoU6df6Q
ic9h0I0lNFVCiFTSty5yg2sYYGbv/D3Fmq38BsidT5/m73vrgW/r8hDD0pIfbFNM
JnD70rWhMtBLSsKfb0xfxp+AswLxFtzevLeX+6QkukmTVS+VmbZ8wjrkAbksf4nN
r2a3UX/Yc5RQ1Guryp05G72kySBjDAEqhcWl5sy2vCJPmWM7lJ76qR42W3fFAj9N
5paNaq+rNkKfKAb+4eP7GpFjadAbjLOABhwmJU5S065v2B3q+c/Ao3JtDCR9Ryx7
moEooZF78Qiqgyt/JENAqSVD9ltiJYqcSY1OpQlzKbR94xXTYuUkABvmCCUwCVKg
pjJL4clpBDx+oZb7hgcUtmh85royqdXugTKLlTnt4Y3tQmJH7pyaweCPRPsM/dMH
KAINqCJS8QGIfopWzAPpx9bvJAhgwfh1Kv/152L1Q19DpEXTCknpJSiX1B20tQgA
ClO2rTD5L+2zDrHB+UIaVmLhh1u+FEnA/t4ctrtz3r94p47inEZRjR1OI3wIxfi+
QrQ8dgSAs31sBehc/uO20FFrl+IgNBo7YvrwseMRpPR6/ymAAYHhaFH7Yxmr5ZRo
UIhVdjTAb4IgzpYo4YD/1e44PMZF8kWzrV5cvmM+jV6kbcJG22S6V9NkxAMI2v9S
HhY4tU1hECzalFOvWZ70G8/h4NTNtjTB5o+FSOLZnGjknAhMn88gtnHv6Oz53gpk
WUtf+ab8q1mpd+CJMLQ0eJRXQ55rtj2OXbCpROLnCi3lNcZ9DV4dok7oGmFf+Gsr
3ggAiB9e/YM+aCktZw2q7BTnsgbLsk3rCME3cGO2Pfyk28ul9Sd/LLP4X0qb9CtG
aYBrQNX6iuxkMUM+pn5mStWdgI5Xw072v9lZpd63I+GTp1vktoSIF5CqQ+lffEzR
3FFOHbPgtOzMjPd+/h8ee1dirYmCyx1sN075Ae1n7i2hu2PoN6G+CoqGVfr+hkAV
j+0p4hWvMBX6T96R1Yqudh8kD7pRd6sKIdTj9NMwKBgN4npfxJyNHreMyEJ6p1s0
TxFhFe+7Qcq0FbVlw9HMYTbn1UmbmDUvxFK01qPD9HVZ1ok7/HfonWd2du81H7va
tz3DEqYQl5aZYfHrRL5LWZvLnquFn20L91n4//x++DL/uYFWJVIUorlaf+lNYZ3R
PzBt7pJnwj4e+gzLAzoaXaYfBB1mWZSwx/QyELL4d2cSJVRxXpbKdF64kqgfib/j
91ixJzrH3YY5zVVYWfQeBbXVblFqLVPE70CydZIKAgxw2TuemqQM6abXAwQOr4xu
h7hyQdhszYM6Y8ARIBNYqf8GgBkQyLsBiMowgmgVUi2peIiPVgIwWcA7QcBi0Ywf
jLDdV5JAthhcmXmKTNsiE7gAV6+8wDJux7zoucLsrvDGV9WJKNAepkj8enjJBIp9
EtJ+WQ9KMs6OwqtSkfRz1C7eAudsLQcIrLJhdlOPliNxq431m6ltx1p8oPBF/lPU
R9YuQJAEQrxirh2p+Sf73o+81oGViguirzjE38CNxunOKvl9dtwgmxUe6Ae9LWlo
mpj1qrOWUGNfU9S1t532IeUFt48NR3hoxI8IHMNhfnBUcrBKxvFa12Gm5Ytqlvcg
EM1k4kk5uai82kfSMTmtDKAkA4YZMB/O1dGqCVWxfgWS2ccXb4b59Cwzk5jePinP
1lUqmshuYI1Iz0n2kSr1ejZd0B69lEvIwrFJzkH09zjMz8ZR7zfd0jGx1T+Pl5GK
IShmMnj3F+Be/cVKMT+kRNZH35s7JVr6t1cKemER18qxzajHozErYJEGGh/MPztI
m6lEzqm3z7qOoDE5y352s9K6kLVkj6Rqm4ehAeFXHdJOy25IZbo8zWxzmYkrG46R
DlUnIvphto798gHI1rktfLGnrrCWZkZOufGAj5odH3WyqLZLiDbgbHtd63I3JUXs
XqFDrwZDQD1HRGYhsPh+CZcT4xAH+UENe0W7b5FXSPHny1kPSmGPWvT3OPikCUqJ
uGEVF7HFMdGPp2YOp3WShjH8dgA2mZm33Em8ARtWcZjQxnqBFuxMAHDS/YdUKdOH
BADwhEyQVkXbUJbjINJsaZEmamr/ZvBIT40ArNtxqrVKtUrG5Mv6cOnWulm9ozm2
MnTQ+qRjWXwa9hnEWhPvzmmGPcFpy1mYT9KXnfF0r3LciU6DY1gA7KsCf8jHyff7
Pi9YLAedHypd6qTwM5SvhwpiimT6ksyqGTiz3iT5lbPngfVXTVP4aqeWp9o6uLZA
rY8ydx/yZT77bne4PeM/twyjy/aYd7YCTltICv0QX8TiFN5feeI8uNzO18vlyxJw
OQWiOV9SB4t2F5wF6CCInfXE3+g83cdjIs7Mpba6fQHWnIb3kdNnLrUfgomrdFVD
g6+t//+m24gpw/OTA+OlOWaLOS3k4FYiGHuPalb68RDw0D6hDFE09xNtWi7jZOKP
mp5kUgNdBQ49TbvpMMRAVC4KKFo+UueoEup49srBDEa49r/3F9Z1tF8dlkvPiu1e
x2PaNDsv2eFzqcwVz3ehNNogIPztHtSO1f3If8wQqq9xILYykGe0i/8JtbgQ+7/B
LgFgb1tScFaNgLXbwFt6GqiJS7+JSp2Z6KCadKzmrhGPyvtUkLG8JrovIgxBSI7S
DCzFiTdgQ1U6WAyZWHcKbZ/J/PZNgNZwYlH0ivxAzm6s55AFFrwSTSpPjfSVlisQ
VFXxuYAqI8dMHl+r+pYjnhymR6SCTg5casMG6e7eYp+kH1F/zRQVzhj7P2PYGyjf
BuzIc/mZyckLegbmuBi24sRQq1kuMqT6wcRISF+YWw9ywwxfngQ9tESzIUtGhV93
K3qg9GFdNwCQR/oCh2BLLkcefTp/Ne8M6Y9WgeEsBH9VQw0WgCVJUYvescjFRxIe
fgrb8NosSUPR9NZjDqelS/Bzfr4GIIofPNDD1tkZBZVdn1uaIs6fuwrqYmVdyZtT
aaweyZYT0UJTse61SNYqpjDIPNt6urPLgEK2LP8Y6sg8GSEXfYCuGDTivvNQxHrc
6E+JZji3xbZhluT8f2mQlGUJQBNsJZjI1kHZi7wKIqs1cuCtS9Cubj2a4HoLAao/
N6Qaxxq2TmbWIMOcEEnFBdaYYUSffnilIZHG3hrR+MNdXGC4451bKNZAK9wBSfNL
NTSsnNK/4dNnI8nXjuAA/YSJ2kjC3FTovUrxhW3kwIeX6Lfuz8DuWu33PcMDtaN9
NTyaj3yJhRLsKxIRp7+foVKXr+f5K04+k7q/sqRAPjRJiODdWyfSx/VukQKh4+g8
5yGw4xV5Sno9gqZAghHp3czpy6WwVUqFSkL0W6UHTaHShtiaeah8JOVxFobvh1zI
G0DHk71oGKFFl2CpOKqJVIN+9snl7VSRivOgNmvlg507qvam7oeA2pyts2jpNd4T
Swjme1BeqI0phc5lhHtgEzToigutufAwghl2C2pNipcsZJ1/JQuLmQgwnm+8rzRY
cCqhNv6je0dEpvMDgnM/p0frSDP1upUd+jTvXi7j5TuJ1g8zhXpTwrtVEJSasbDX
JmsjHYVcuEMuzZ7tTI+kA4l2/oxH004h2KSeehPup5MoEG8tX60DinMrOz26oHLa
mJqd3YdV800G8fKabtAQTMkkvjCDvfQrdEVz2mJAfW63OHMdanQtIaOYyAUFM/mQ
YPSxbLo9T6GIBAhQcBtKIpm7/bf6A/IzOo1ch3s1sH4yHu2sCzDHA3VjQrnUlYWW
MXtAOpFfGS2WeygphEgBhe2+Rn/Js9rDLXMpM0xJDw9SSWhg/b/z1+n6qGho4aUP
2/K5pbCO+Uc9l1yQ3ivQhFkKMu45AdcOvqeO+EbFcc6hTOo5gRoS16VaxyQllmzS
SZUFStAot5AGYDe9Dztg+iSsY1Q7U1sihzJTT1NBzm7YQxu1YhB/P4omjYEz89gu
RMj5Y5/62uTLdNvyXa5n22mlb11maOmdx6hGBKcE7AKiYWfZWncnV7QPAU+zl2/K
988hQkBDjcICljDi/pQyrQ7WRpLXamQuCdLdWCzE/r/VxW1r8XA2UCMJdPXQSKAo
hBap+FhbsfY/BKP6OAAoyo1z4torRttu9+4OHhdXGDxWmMu7biJCOnCxP/CQBI8f
R2G0V9W/pXgwsnm8s4nS750+V3kcp9OQ0t9gJGmTSrLhhPAlaMzHlWFaLHySTyQl
83zRrdV2antWylut2k5v3HVjDoUX+r4vnuRL058VEgQ9KJp41nP1aSxTiwsa+wFR
XGf1d8RP6p/N/M0f7LZ9naDzz+sbQy81jKix4KdxW9joUw+9B2lNAZnm4IbkZbzq
JFA2ZNJhrePpDK/aoHOWNm6QNSsHxNWjvy7awBv5J92M3XadecrOBiTPjxyxSNpa
ZImKTh5WVbq8DuRvFtIA7RRWYKAmhs3FP3LjVlyZk3v9V3r3bfKj/z92brOC13wZ
P2V7S7mENix5se5bDbD26KXoJm4YaAI01tgoR8tuGYWYdCehhMyVeqTrfxsywFYW
j3pEA2CJohWHJt6cD0RK7G9E/js2fZQHcbnw8EnwwPtmZT+riSm++ecAPvqsH32l
My24zf6wzz+7rR19I2YF3IskZW5NdGFNkVVEtCQszNUVXoG8KSgAbGmsZ86d+sy4
2sOnUOZXWjXmJ3X3VJM4aeFK+zjCVa/zBl1FG/3PArGvYCHWGMsc3z0AmBgT0NTX
JlXa8wqZqa13HRp6eLJ0uRtLk1+TV09RTDNgN/EVGLmsDeik/R3vx/w3HXN5Ie+9
Lb5WfENmnqs006e0qQ48yqsao1IuRg5Ut+nRVnhvXer2IpqAoKe+yKnNYOrVKR46
rz043QZD3sdsIS3YY8HT7+jXwVoBRpIg8RHTQPIxxAyM7d8VB9hDalpQtylancGj
LfQyZF/G/tfVSxXKk5suWy9EK4x4yz8WRYt8S4RJ9PlIJ1at6EjRxpHokb1GxWsh
VnIRC+Na0KF2SeY5m3hEXnCxxmStj8LB1/2G6WGT0DdOg1iw/Qoo9MC2xFfYP6cD
dLIR2TQALfp7FHb7CHr9VCFbS9nFqUgQzPWSjVyZc6oR77cVEBnUXuOvLK+MnZ/g
P8H9I1J/OSXDFQkEog3sCSejKeSUYokATEk3FAx/6YKDXDdLMfuPmzZHTNPWYT6D
wxLE/SwxH5cXGvtlw+Cz4aUOfcuS4btCaKHr1j1Oxr9aBejF5ctpClVSaRylCCWY
67ddpESJ2pSIsUP4Jr6ed3IcdSCypf1TWi6Txs8b+WU3DbhfnFKfnG+7b09bQTzX
CrebRTt3+nuRfkI2ZzB2r+mDFKgVThB2/g9WQrsgD5LmmhetQrczfPX74Yn43Nay
yMr8K9CVfWTNbUkUwRLJS2Cyv4HoAFAlTbQIJRbvRefdzA4J33tXbShlCsn88O3S
kiNDF5OJ0L515sFKnQwygOQZ8D2QEbEOP4+Gjg/11QJrrWdg3AZi/YXFSRG17ydE
czlYxHydQmi+HAxBlveUq7bYRamBIiwQygP/Fml4TXbPanCPxbteMawh3geNyPzQ
r5m8cQ2MeY1vQPQe0doX8thq79YzSp+rWREdQIhPiV4jNeyRJbV0Ht1EKoCJGfAY
t9KfPwcv89RVnWcE2t5GTPeoguSLA8xJ+SAjKeIuu2VFzd4Cq0GTNQ9FYX3cEpNn
iqkg0LUpzrdnVmqHPnERqCD3tZw3NkuZUncIhPxQaQOG7z0iSXCyFFyTu1Zh8NxA
EGsoTouierwLsZIiqwa7wegPAVn/nRFL3uEicYZXexeSMRx8P1sw9YmJwPGAiy7L
ugiGM7B5+T/zylS1upeTvRsTDwlESatzIUPNiBr8n/aSp0T31IDv59hLrAEgPGQJ
OlwgeJvpWCkAA5OGZX/qrG3535MbA9b4V3TKbXYIABYI5Zp5K+KT8lPdcfKkv5SK
x4wut6qfvAeCY9HhPoQUoez/1IFq7Zhisr7U9GPslSUQwyGp9fw26bceEdq7Aork
PJ96kqWD0umz7bLRPxCUzsG9l/24okXak/30W2YZmdc1ECjVuqjQ/couJrV8a0oi
RM2ltcSONItrrVFq86ttSa7YkPZbWWhQu+1Ojwn7/ad+sfDcLOW4/s+Ml7pcuKkR
CA8qk62qg8VV+5hoyePHgFEhUq9tZi3Kblan866ciOtO65GpObHDGtNLni0grjG9
bVSBKsTlocBkO+qcpOxJciC0a9TpHRagDqMkVBH42BpIrAfgggd3Ps9fUSWwMbk+
zqbt/xdPygcNF6r8n9Ax3JPqNPKLm6aA1XzH6lsEkKxR/Dn/3Ruy15aooO1OMz7h
fniBWUrqZl5WPQostc7b3Y/PfmPoowbVVQSEkDKUIsVdo2z7okZR1Dt1hB+5VOb7
OBVqSbt/MXC1eBoLPLMdGAiYhHuNF5CVq4tuwkpO1aB3W8NEp4A87rHm4/0pj61Q
g9HqiTDnpB1jtioYWkjUqTg/CjRoTg5JFrz+g6xpLenAMFUSq5Az5xLPubuFKQJR
EujGA6JkSZuKxY87vY8UPbQ1Ky+fToi9kMBiVyD1RvBcI+6jSW+kD39hYjZBKE03
RqTOB2b8v1wZa7AvHBMukk3O7zuwzEieJT7wvDsRAed2sBFZ6eKh+Yn/icWitPgg
i6owxOBk0pdcwBkDgOCiPBYO6kZr0uzI7Xj7o/FoOTHrH0CZbpM0zATeotHG/qju
H0gxmtjGsDJZ19On5jpwD5g7L7Zo59GrsFgK8OYuUy06NBgp4q0zZyYmL3M5U01O
FgM5QIKFzhyJ805dTXjbUUrn3WtQndBTbV5+1XAnr7NQCc+mz4t/Ux8vQv38IqLF
fVwsmY8cXuZP89eMDxcwSTmw4UzoDj/fUBo/QvBeuZ8gyypLnO3DNKiEge4IATUV
ducmNH8tCQ++tuBNQS7ozFRzzY9RVuCMUkMqXZcc+DT1F8vSb441E5Fd40vJd+DI
/FO/2JeUgTG/EZMlYLM5fGT+U+ZuamD4vFR6S00LfS97onRB2YChL4dEs9HxMMFB
GoM6CuwpK6ZUCi+sgY7PZ6dpWl7FcKOcrYIGIYw6WsSzsnt3pTUtcMEnlCbMORdL
ZFE78dx7ARSb0qe/269qZAZxIBvx4LE4uvK+U+qL5v7u9i8bc3FAWmkzPYEPIEjT
PzSWcIaH+xpabuwOOnOteJj5VguYBcjk0RIVEavzcxGGgPWS7yckEN8IBUep/9Uo
8iRTyCiP+1aKGVvZxsmZGz/I4yIJxVvaqr0wYPQfpfrFqfOiIFhZKklDawqWS9hp
rJ7sHpDZdEeC8HwVf+EAXKvtNUGQXWhMs9/Izf+m39dGDS6BAvFSCi2hbRsTMPa/
a9ZJAq3x09ria8EsjFGaxs47X0dcBKNb0PcWHF7vu0Bdh4Mtd0A3vs4fvC8Cj6+R
WXfkvfEUqUTG4ERKT8eqUbAVcxDYbAbvpsvlA/kVgFxgy6cxkb8hcMM1wrGvgfX4
sznI0YqHcvMEyLTF+LB0xtmpc+n2rLvx4dvVNtq4PKoSIlVToxtObOviIFlpdIg/
qnlsfUS/cVlb8MNsP/pwQBi8w7/MlNZRP5WacrkZaL5eIL7wYDYlF/N4I09Qd51w
P0M2CaNJOWcE9y7nOwmcqW7M+phK2cbh9ByduLbRC6NAVnPI0zUXXbjHWMHaLz/e
tX7xgThSHCtvpBZA4riR/l/kakZ4wSRqqek0y525uIVPhwVLnvA2KILnbkLOSMpH
usZTzZx618CQwqwkHXVBwZiiBvdn0j2mAxz0ZYccaBZfYcKpJanuJl3l7G4nHxVS
y1WIDiqHskCNEXQ7UkVfOIq20msbDhTXAMYt2eIIyEhIFbnaGsYG0jFATZ6+F53m
kAiDi8bnOVmfGdpwzbB1zRSt4+U2ATRJWCy42GUWL3g2evR5hPGgdCG5FSa51/GZ
H0UMm7spQO1irnO5PLWC6o85t9M4N86U9DpNZLRB47O+G/Rx7dguaEbKTPLzFy6h
uxQ7x5B4CphlEoEMpAQYNYs/UIsHGJCsurLsORPZodpl4awr7aqJnIcmYSIEFqGa
5BJnxn1W2sr9L1RLDVuLzYUx8B6Os3s6ZUQv0reJMhmfa/86pBZNxaCxEVmNRILc
mRfsC1usOhtDL9rnAfvGrz6Qi75JGK3BAXoSmGZZXmqpZ52xXt9i4faNvev8EFiR
fJLhwJ9/Lt/VhrCLwb/nfDV2lpPK8mEilYy3O6r5NIVRbpmxTQsG/g4RJ77PdP+o
JpOxGjL7lQXkvafjwlHy7oPipP4h/sFkOmgTnhnoR2Hki5/vnO04LQ+3N+j6cVxb
vFa/TEW630kzhxXq9pPfuriMIc4clP4+YaSnEQ0e/pVX8vAap7wCbFUEZDqrL5fq
pn18rsc75XShWk0lg6vamznAPJAiYKf9BOjBXjEFAyCQjNu+6ArnaHmiZlMk339v
3EWaOXoVUD4AipXwV74r4GKwH9LhMu7pOVwvaqnAzXXiOB1FdaH+0WDhKMPwO/Sq
5f4D8LuquFj1nBiInIFNSn3ql/r7PSaE/s1Iw9k0rQzCl2oQWVUINzME4NG41pqz
zup396ZvllO1Tmg4Pn3RuT8hZNkHz05JO+8Q0NeRbZ3XHnZMoMeStuyVSXOAHaBx
1zsNxzyumfmYQW27kP+9RVKJ102z05iLvlLTcP/o79IaaLUKn7V7DoIoJNaUc1zh
hP/BDSpRw6LIgdRY+oRdpZBpYoDw+hz+XRDfx+V7r1QYeuxfZVgC+bSX98RHHlpq
VNv7mugA9AYi5awbg90ROe6n1IES9gHqs02GIedW12xEkibKMZP1E9kkuw4H/Rq0
0Yjpj1zmPtVSyv2Zu+HX7LWF16SimteLAhvBNBBgdi1o6tLEN1aI12tq4/mYWrCp
yaGwh7hpeQDTWCrU8zztkhhh97/bev1p10wzfgh/h/yBYrbGbQXzuroM3uEDlTq7
J2sbCaXOpdVfsyWc2Lbaa0OlwmBajXJ4pXkYSkPp69j0qJ/yDVZ7II1/H9ljBT1k
HvL1rwDsWx1XJLvESr/SEMKPBYd2KE5mNmLH5XVOaE7bIBcCOhN6+G+AiPlQSZy5
cM5cpAbKnZDc2NMcCyjOP0uLsAly+7dLdvFQinSwYNyZu7DjqSktHP0GIXru0/qD
FFS1u9nAqsDZhPHl1rAkkzIK3OJnhAc9rGKpXs10VW97rWR4dQgqo9PWlaNdDCFQ
lPoWvQ1LmdWDzDSH4L5i9CLofzOi8mQz2ZEFkg/WWvhpW3hocJ3pMCjkMMe9SUE9
QtKiXxsdqCivwrf6ckR58R6AfmxLnt1+EXyMNZSpsdf/U4LR+FU2A891wCB9jHcn
rxX6Vqo9JbwPG5wbeGJc9TMgmuAmSjbACLPQskOuCNZH6IYGmBVqQGTnq2YtNmH9
7UK4KWnDCLYQM4vaT1ejFOxSoH2YUx79NL9b3UQm9gZeqKXnxtWB4TfHkMU6NTwX
mShCh/6uPKkZXs4kW4DWRDbYwWVVFS2DziyrGUUGDII3K6plQ+e7FQI63C0CE81m
aknEAODCNff+gO2tiRd9YvH0goVNivi5NrTMPGN49KDrb9cRPUG6dsxBsCDueEfM
TT92tcDS+ky+45ztKm2h3K36r/BJT2Xj3GU1CxW/nlLBZLL+xnXOy+9bbU46As3Y
GVCOllDH2WUo7F9j6N3PeV04oFkYHX+fnV7l2Dq71gJvOni6RhsWx1dexFgU0xQ3
W3quoskZHwkAd6Q34HqSeWgtB0PNH8U+QQEvJ+zwJPF/xJpIvAXYkl4YLVB/hvnM
wWESZ8CmfN5lpju8iSZi+B77cHds++pSq7J5O3Ry4thquohQpNg4CvR/ARnXjOsV
9nDxyOvs0w7Knu1K6B9Fh4QLUQlKkK14gZ/popaXI2y2b3hH2n9QY9sKI5I2O8Ij
5Z1i/0ZaLoRglxOzw3Hci2d3hPya7v0QeSt3vDYnqVXxLQ2RnXwha9/kl/zGy+zI
2xryKxxFu+0kAIORUz9heMtZyMwtH/oYmcFCy6sbGGFc4jiwg3kgWtxuYkUCfhnh
UWXk31vwuCdt82apURAFtiDZxHsmcqnq1RwpdgmzQbcjPoaM4xejuEU44vTFmg8l
pdSuQBmhrs20VbzxTCAeSqHltHNS8cDY5SMtMGADEtq6+XNCQ4XzHUT5Oo6cZEbQ
TJB8KD7xRbbtqZms7DZLrfl89OGwIS188U50nPqJV6bXiqyeytTfry71KkfRdgH9
s0y38msWw03LHci5U8ZS3/1dsoZBK+9u6Uai1XYv9+y0dUbxvv6D+bsIsI9Jdxfd
PdAsti4RNy0Zr8qvhz54/KtHWrx8f80ebT7hvt4RQRuX7DCcLbZVUQEGaE/IqMWq
KOdOqEi14+HhcWCDdZyyI9Qi7HZ6842pZ/ESzF5KGGZ4gVfap1Hhjq0sjHf9TLMo
SL3VH37PlAY0tb88Ms9FzVpl0jke5v/+NlbsnG8nuo281Cy1/rYyDHPKITv7w1kH
waaegd/rvphjND3FvD0hpCz3EdpnjVTd8oRC2nr9MzxRkjT6SVAa1vcXyJ/FRSVl
jmdoUOANvjkaugCxYQRuyQ6JWAc5GwLUrxn9+ZyMrEPogI0e0hvpweOeXIhbCVpV
VRZCtXgGj2MHBoF3ywA73ag1VWeJpdEq6xn4TVJAFpY8TOY+bfbe286yDbUT7YXm
WOuBRzIkAntn447zuBLwukexMHjpn8ubyXYg9eM1MheeyYQ4sQvfnfg3VOs9sK0C
em/O/21mPRoi7NPRanm5gd8GqgpHaKP0ipae5ZyXOe9GZOAYa6u1GjyLYsiGGRep
DCnNiwAO5e99ccgubQwtg+rVu1BVTeCXWNuiv7GZUhdTC3eu4SGitNjPpTDMEHfs
egg5WB0bv//yQhZ3Xc7+KUuyeHVRoPn3eO1GrGj7NSK21HqEc6ZbZXT/lBkXl+2D
DyGP/Mmrw6pkwrMkXm82dqlRXroPcJCpmP3cw7wHT0ZLKGEtLf0JuYCik1UXs66w
uCZB6ncMKSA5bVKqQR/sPHjqMXlTGN6w1+LV2UzbaODNhqbVqLqQ7zRWmbcPTlXc
TZg09sHFd9AfVy0S8zUu7jkAkKP7y0eh5TQBqiXoDZ2PHoB5KM7L3GUTheRoAI9u
EEhAOi3dh0l+CboWC/9AVs8KWbL5ixsq0VzuarXNId7KVoiqG8r64xFyfr2APE1J
B7nT1AgtZoaQ5k76NKC0GnKPvyy8A7/aKsF6lop3BmPFKiKwI8qBGq7W+JP866/8
V5j9k3+FunYbNMHebRi4GSML4mezXfdbRHCaQOTHpYHm14Dn9qjkr2VSmON/AtcI
3CQzATymwZ6bJT+e2UPs87re0slgMofsh1yuv5x9Gxj3i5N886zSA1TtgNrhOXiP
afjQfVTIOUwK8bJoJHS+YNJ639PqmMaykvn6w9eT/fPU5LZAtwAwNNWoqn9V2chG
zzL9dkbQ9Udsi4oZzfG2x5Kaq7rQl6A6HzAEsKSA3+NUKkMK5FfwLXxpCoAzfK+M
jnHCwNxTVc4q/q/cJ7fEkB/PUXfDa7Wu0C5KNvtV5r54AdxyoITq+6Uhp7nToj4Z
C+nOf5Zumu05YuAs+KpCwE2DXtPXQ2nh5S9aCJx/4X3/fCiTAiZnewEh/GGUs3Jj
NA0Q/fqEbgdSmVqkja8xhJLjsbY00H67rc8DgSrVJWsohxovfG1K+X4kB+KrMlw1
y3suFergDTW07ScBcXlIvMxgIBCcSYdlkJd2hJghsojwlFFs6gSOXItiiAkqi+XV
gC7ZpKFsvy0jQxc1KpaTzvxOd5o7dIk8KPcG234XjqEUXeE3LVQccGCvEX/HbxF0
KX/M8QaamBcAJlK0hHfL+vpU7pRmvF1RkWhBQFiiRSOSHuEl5aAc38t78UNypKeQ
PRrfGBEFcgk1vxpasIX516N/jU/py670GLbkMA5q/OBb/PyXDXtQzOyvZOarle1O
TN7COEBjiPVK3JHmtvAn9UhPakRRbLP+8SVIptBkVEuvBw6E9ytlEHbHPY+WLPHP
4CUya5//BLujI26yMBp8hhOfkBxDBpKERHWGf+bb46h5SDXIbBuxYQkBZ840ICGN
VGf06fcmJpPcwXeiDugHGrL+va9++PFLSqT03BBNx0S4wLbLj8o2OJFfu3Uwtx+9
Eli3Q361hIaq0mgP0ip4/C/Z+uGC6YHtFJy+YCX7VSPiVSsDGEiWR4KcYL8lUMIW
6lF9EeyIsVVwQn3bf26IZO7NEqwYo6Iq07hBSuHnAfuVZNhElKsS1995PNKrWoml
RTSYXt4204ZFf35FwZSUrjPI303TyQn86xnRzVDL2758UFhJFvOEOmuUDWTJdfNn
/Il7RdICQHWFuilSvTzeYVqYD2xC7JLdokOeHhefOyWeWO6h9+e8vlWEy7/R6tzk
1Z/+9j+qUOG7ejkIZGQUmCrI6/QPezZSCu+shk37NqjxQzRWzdmlqU/+Pfh1xMip
Rfw84uj+qwpWPZjX0PGdPW4xeFJW5SSXM1jc6CghW7zV/pS1xMN19yWCG+K6iEQz
511l+uR4N/ua1d8GmmSjko6TpucnIDdZg14hwF3bXiawWMR86Majkb0+fXfdkG7m
3KRmYohrovwoe06kSxPbF6y/fRs2WofwxmK6ROKy4A4QnmP3Cux9Ykx2pri09rw0
BhzUUWT7Z/sauJPPy8f169t+e6RTX99qrgkqzft5J3jZbE+HoKksSDbm/8+EY6Xn
XqrbSxJ67PJ4YQGNVXih0nvNBnQTRAB13j2h5JS0zQh9Ab7n7QBvaOWV5ZM+N9Vs
6Px63qEF5ICwVnlpYYSnSaA+kqn3f97PALfwrT7NDUCLSzazRgrSjO4Gh1zsS5zk
mWdYaMwthCSfPWZ93MnqQPXpb+ByODt4oDDQPmGigQogmFaPMJO6l2r4A/UUqk4n
9JxVDjK2DeSAbQdMvK5Z9jxJOcK//jMuLc75tg0qC+qJcNitQawNLpJX1k+x6Jms
1JopBCUkMYM1i3mETbD3hwhKfbn3j86BjDRYmEl52lhjFg0d2+XMIvzQDfhmsohV
IO8x2YOjm+rkscwerbbSaFYmLG1jDrf2mznhAMcrGC/jIut+gfTkwOmfwTKhYgfK
lfJqtuK99RVINVqbYIAGizSBfGYCicLKBACOLSwpAbIRl/yTMmTxySq0WmCLLWyi
we62qB2oYUow9zf/kK+BCar43bFRm+ro02/bO7xQutZ4OWbj+/pIwsA+wgTt7zkm
qMOowT6l0vwweX8+ejJ4K/GPfFzHYE5IrJpxhEnImyxRJxe9CZ2NeQIK7jn/j57c
f+vb3J+zEzSvJmcd8cOAaRlTzvVVzvV+EdAmFHPcEkipgHG2eqCgtBQxpmytiG+e
KQSMQmMD7zi7Pw9BRgCVr8z2DjRfVfdMaD8oZrZlLwuf9IyY32cMWwObQ6vmp7Vp
IApM4LMy1uftpXeEwyTEvau6GDpTjsOB6KVoq1dtoOwEoc2dr6qeSCcb9jXhE+J5
XRxBMz+hy9YEx4F4nt3/7+tEb6lDMXy49zWM6EWWvcSGuObg0RSXJrLoaEFybnaS
iJ3r1YD6to1KVsJ+nUtZi35CwQQW4txUuaBeBbqn5YlQN/Kd8qIWWCoDkKy2Bg61
gSzUxwDr/kOTbtLW3NhXl1xbE2Eu6s2vx+m56CUm7feAW5xUTfDVxV0MzbeAWy/b
UTvV/l9c6CIrHozFccTbQm1Axg3JJi7cuRDwbrvzEI3zE1IySvo1rW6VbeO8VPxN
sr4OInFJYO2GDNFVxiJ+c9Dsyd4nT6LncToGWDsUTvnKKPuHQqlzF7KzrjehG6QX
OMRaAQmAVVyr5fSybYM73Vir8tBjqpDH2oh1bubNLH//HC6+CrKe0jd/utv0LNeK
O0y/4as278gF1w29aOs2MEOa7j0v1iIBUHR9JAzhD5g1lergGcHkiSN0683ykpkE
Znkiai6pbiS8gyo3PryPvhHSEr5B/DFwxi2KjImvMzlEWTIJ3XBLVFDZM0zxU6F3
ILAPMK6Rbj/ZNqFVN3a3xodIn7P91UPDKlLY41hvr/sXvLKw59Mfe812ux5ZfQ50
Bhd51915VQP22pfjtXBUAw6yD+km8uNjKepjWPDknNgbRwEE7t9F7UulAlCZUXzT
QMlTHcOv+yXbHZ86lUgjwAmscfbwiXDnwduVFTeW3UELbe6LSu0wn1omQf1lY8+E
eD+CKgk5snlfVEebL6PjElkKwVsE9Sy5vcTOs02NcaoysnO4p4aEf7lJMeazuVof
Fl3ztHF1wlj6lNK3PE4JdObJORr642FBaKB+KfhzyoEz3Ii4i9kx/B7Qe5uYfHWs
wpMS/Ltb3sApzDEKVTxWsAdiJlHmPSiDr/aVQG0x5sHvJ2Ask1YtVAEAvj04mVnW
2VkxUhp7zr4sbVizW4YCS71OwyM5Vq8PSO8LNzpdJGtj4q2ke1Up84CnpztBRp9z
sTXngwnZI5/42KQCdztSwPCTJb2nv/pKhHgFEq/TxoEtzf8NJ5uAV5J7ZIsDCM+e
UKP5aK5UZRDTmuE8l472cJ4oPrmaI1A55SDtN6CQkpmjh3gY22ODSlm98lMUXUwO
fTD8dYoum1NpQtu2CjU5juKHgEk73OVI6iMkB/V3k2gvZBFoUAmvcvbsNm96ow/9
BsTTRU08MburR1VcY6D7yFha1M/yisLnW4y2dvJYkK56Vg2JyiitZGD7Ulr3ek8u
VTJynqId6PGDEjUSKoi4pS2534EtH2R439/bJZMzhpoz/k9XQ2MvmnBTKsnqx101
VCDw/qqHCKPhWgfa+Cu28ceWm+HzYr7e0y8Q7MwLDhByOGUffVjGqga9rwsE0jJi
0glIR3QLT/eOrvei8Jz1eiqzJLjvLQ9wmkbjA1eeF7t4XoOa2ku5KUe3YhyASzK9
gr/vSIOG87SKrNIkKmNimYsUrn+9XDtTUDh2PQx61Vn5s1Shr0uW1vKaN6KOohD5
Of30mMgaULCVBbIvID1gBEW23Ag0HQfrRXpGtO8UTmJqYIXMYxlnEm3K6cSHj0DJ
ekHzO5Zigttlo6OtiS8rQ06xq6OpjCsrIdgzcf42JzVQFwLFlfypwycePgpocmDu
+s0mb2GTfys4bGleUu6/YQv9woR9rkC3G2933aydNUICHWEZ6lNjlot3AC2TexrY
VZ0zhHCAAIvR5KxDibUYTK/u5KBqN9kTsxc2O5zoF+j49a7GOmJKNk5rX8DSLm0f
Rpgal+bV4RPyIYmNbqbyNjZxqqOe+5+iypE0fhW6p7fSkBWtU4JOltdczAftFEzD
AalJo3Xnki+oQQBDdpXcmAoFDZzPSCKjLluhjDqrTodhCoS4QEf0FXN94MynKN1z
8UzUEIA/NJry4gtXJh+o4s0wM7mQGxxYT5Y7A2iVD7XOzOf7mCZ8JxqW7Ea3EXOQ
bnLCu8bz6dxGFKA1WvaTH4Z7IFAHk3QYRBf725fafPJ/NV29kflW1KDdv9qy2T8L
CVhpaRl3sksvx6FpCZYX5ZWwYDI2Zfx97DMPWl0IHwFYQkLu1s6KJcxdL6plstvM
Dt9z0Fn5odTtn3k/wpwt9xgI2+VAOyGlioZNYspFAZUWJgHZpa2pcJ9ALlRnpSJN
3wDrcOhqS6HYJtxITE33FcWW6o7qxQjGbA5n5gb9B1Nlm4Z3Moifp2dYRxpmQvWT
Yq1YUXwa5J2gJcI6RERzhZ4eezlq6H6+FDYU2bDnAldprmd7o5++FSyyjZmRWB7v
X3l3NG62VnnRYZIQExan5y9htRoAaGMGZAhx7DDZWZj7fnRQGiMu2fISiCvPzcrf
s/QYGaSPT8LFK5P8+lTBHA/OxBMpIlpL+BZVhxUfLZ4FMdXCQCU5Kap0NStLgp15
rupGvGsfZZcy1ccoqoAVjGGMef4QsTuUpXzBi+A+kZ9o2QaIt5HFn+yK7J0RSnVc
rz71+jLR2NERgpLUcMZF0XWemdMRUUSs2rDe1XJxoMkK7yGTdNWmuImzCMTHJNRx
sLI5f0K6cNWaO8I/zhv8LJOEC92YAl7u8HQqEhE0KXsJSHb0h9qEb8DlQvH8G0P/
GUfeYBi4ZVWVnMRu9sqVP/S4/n55E1IIhfrpT7z/Syy+jSWk4w40j8oGk5QplmTI
Wb2N3V+a7iLnGzcIJ155vkJ8C74DYKenvFGlToMaJ1mjfvcvK4nO8U4gRrlUu5uE
vFbg6N6oogjvRVOLuhVfbqNDUTIDEvUEgtGOV1v/p+c4zZ5V6S+4nOG9Kg5k3YaO
KtFiwGfsGHAkc36GlNjLd7YMYZDmvopCPcZaUIHJBOHNCL43ort/Kr7vkbay/3Rg
z2+qOcJcAZxDbGJqEW4Tbh4wugsxmWeYnB+tIZAxkNUzkb2/h+ykz73MTFC7U1W2
4AkDFlNp5iIOk7PyB0Yr1wiKBtY71gqQN1uN+0ekso8PsBUras2EnQpUC4nkWeLm
KvEW+60748U/ViDprRbx2SrlWXtoIfYjOdD5UCJz8EFZaOXy7E3ddyBAGV/33BOt
4VoZnZSLe4iMGRbPBk0U2nvUBqPApsPikD/3r8Jbsek25fqk8l2K4sGpNb3DdIaD
PN/IaVDfyF7pX4nrSaqYPkWSzhlyBO9ze5G3VsooOENU9UJk1y9b6Ni9BRWdp6Z1
zG2dwt0SZhEIZbymsakkG+2x3vG0BytdEx5AbbtenHhoaIrVmpTii44gyYaGu4+w
XPmZ1KJfRfPo/MiqwUyTTEaVzPOV8LZhy2KSpfkW3WKv3CNWaTk+0nRameLlmw5j
Tbrpw6VD/8LUhGmXFJVBZPr5hMR/28leg0kpYAMeX0u4Jn6BJX4n3qSnbno7S5rz
8NHUz67991ZrMonUgIcp11ixjgHAvXohjqutHWfSRKumlVJGTWJ1vwI83vmF8fvx
Y2tFC0tBRgiTDQknPOpBJDgT+iHwHjNA6UxZ4z0oq5eUUe8WNdyWZLEDnbrVGY5U
SJdc/4hNu1dMX7VNvBGwGb1ZSyL02VjwbKyEQsvq8sRVE9/bkzcivomVpsVquw84
V+WGQ8vai2FtU/Ko7g+1IuaOg/Rg/DQDKVyO4vtGsmBbYiqDiqRPMcvm2DRAt1hv
uXA2Bt/6FDkaSWwOAbxgBaicBWnCty0oSgQE8E/KfUaC4xuPk7CxTdRjCKMfFebn
b5bEyGAyTBnxOHTzTiXhEcMkbngap4aDCCD32hyJzxrz6JRIOPAKz/GjtMGwM2WE
qPYhkOmbJgeqorp+oeLUmnwVwy8atrpRSAiHMVQy3aPy0KEA/PZEU1TGd6Lh0UL6
CanJxPZ8TmFY3MWHxFFeeJfEfcMuMfbANEfXjhOJJNgxCjydLOe73yVlENkwvpGS
R1E82pyNy726uEhssMWPLzwfuXq1RQ2z2QwSlcPLkpQo3mZihJM0xCYCdBOIag18
0Kpwsgt4ODg9+6hg9c53h+JD1mSTbWTjy8e5I3VlxUoRNo2tYenahAMJmQmIKa6I
8+FS5NvVKpu9103w9iBI8T2gkonRNI/Dsg97Pi11l/YHQ/PJI/koU7OqsJH3ZvWT
4rCNmyPsCIemjnDhRJMV5j10tM67GgRyLFtiqmQe+vKtcSNsr1kEz3ZB2yI9GaRh
j7+2g/uxvo5z1ovgpMStpJBPezeAGDlF8lleQCHGwPi+DJdSFSeVi0iw8qrlH6/S
SQtZMoelI/MFq2UPTc/cohOcrVnkq1HuIhVxpRpFD03q21uO/pwNvqmJ8HUWEAvu
pE/8/O+eZ6998sDF+ascsECjBjH2Nl3AJsY+9KUQ3AgMdLTKOKgnkJUmwONvxNrE
kskvCGhtVoZZwjOhqYUm+C+/Q0VMx0nTIvzkdshK6ilB9wrmzpADE2C3Tdp6yXoX
wAcGNPlezzKcAZWh4PLXzk9Hpvddfz4H4c6sLq/S2+pmIuVj0MmSWDow5u0qxC5m
Hhs2w40gydWyfdGTiMwr4rPtFu0hLlM99PiMVQTyUctkasYOo0hmsaSXEughd+Cr
bte9yZYahgSWQIRxGurivKj9vVFPq0u1gzp0llZLOwAU7w7cm0/3WdNnz4nlwVem
f6kmvrw34X3MnOTfORcRAsE/5+Gh/x2k3jAgUcdp8vPJOEBTWdUtZ4xGtMCG6SMo
5PRgePPyWgmdlP32AiC99aND2USd0jQuCtx9jbve2Fl2zof75TqeLL1ayny8WXpf
KFISE022Rl8A7gpGBWiau+gBu9nJv5OVBoroUBRnw6lMO9s09hnymUQouvqL8tT6
wdMk6new8dnSwesEeFMz9qZlRDe/uZOLKeTm0CnIi+w+oRyL0QKXPViExu3a6d7h
IV08FWWMUsc+JU91WdaWUCljN5aYfgwhHDoAliom9khMQHh718u6BO0GWhCkZAII
LBpIiZG9nrdhJIgp/AiEn7SfAw6WJoSNNIJunGvSxGmZsOnNkP1sDMYW/S1IgDK6
PYEPXeHuhbg9Nd2mgehJ3SgEMkmf4i7lqJVqhoEePCh3jG6LSrMFnKgZHEOQTyyf
I6+W8SUfacwcYkIN11b+mdBnA7QpnCwcoqjaqRBS8nxHUg67N8m6uoTAwkjTpp2s
HnuiRoqKYkz5pZnbC4F5myGsmxiwnqeJXvQrI8BoWyUH8kvvLug4RPA4KP74QRcE
7UQU6FSVKCWubd26woZA/ObvSKN+7/of2+2/2fcB0lD6P3wmqYyqVrhBfJUUCn4w
CbZyz8sTuzodiljv2S2eq9/ejwKdDgsUk6VI9u7anTC14a82mVJItR9i2ikDK7n8
2+SrOYuyLBqmaQ4L2ryF4M/rTo7MwSMYPMP+W+gEVTRqt/r+qUBjNmmJevinD2yK
Ni9f4ArA9y44sPsxSIndRpyb2hkSoMXej1q5kOY+1bshlbhO0W9J5q6sowNnrMK7
1kou4fkciwgciDjF93bCsFqmBm91gO6YQQZO9DOaEu1wwS4v88QIBxvY27nO3dzN
6DLZpiLNW6a/P/AAkgE2MvOEN9jpji0YtJgwSqC0prBFpzBDtcq/N2lJUTwc07EC
/BD7aLqqILKhHCCUVRqs/BLxc/vRIxhhq9Vo7EA8vPni8GX2yebIE8hZ5nZXA9Ja
UJy2h1NWliLy2TbWGgciS0v7YnuIjv6YJo1GIdF46agmbDaMBOAtnmibvtFaCW8A
Cya0Z7yuEHCU0zmhTMF1t8fKGXDlVy0fPsfD3MPsQTok4bC3f54QXX8xi/irmJqH
O82gyEuZbM19COhbfu1hOG8Cjg/Hzg+ScQFtJi278ntOuJ44r/1jy9SeBOaD1iQr
hO4NoB0+0ZNvKO9BNIKLSGHl7eOUL00PMoMjwR4pkliWomLLeTqIBQfwD6IIUBZe
nuMzJz4EwchTSJhPPnumQ/x7p7XP6b8BCzq3PvES6JiZxPOsL7Cu0h0XcBkXyPRK
Qv06/IyDASo7/nNoHseuGcpS2aDH8qCL9lFX8emJvuI8iNN+NjP6pvW/uA3j1tkj
YxZsDLYkIyIKwRcrNpDQoeTfu9jb+D6o4gcIboTIWoqFrCYxBqmyz7sI+Q1OMyTZ
Ien3cQi3xberkVHtjZiLXMRWaqmqJOg7/3QId+HTezxv9KXnxwuPegd6lBTRyqYk
rnqyoXB62s9ZoWUgQdZMxW8nSzK9XpRAmvE3z5tVPt3uT3P1a8mpnVNbyWZ6n/sc
n/x6ihrJvtMNWCPG+XUxkxTVAlfvIWu65jntvJvF27sNbrVVe/UvtkwWkqyMALQv
R7ohcXcioVMcOmA3DZNcBKjhPLDmwuMAqeT8xUHQw3sEI/XSunxPz7KXBBiewne3
IBM8nD+79JlH9+1nSCNXfxN8H2UHLpYb2vCG7jdECmbVtF3IhwCgTA2BtPwe0NK8
n4Ox7cBiJiNDKOuFccD2Jm4kzAxr2WFW5XhXd1WC5VIgZNfE+NvLbIpxB+nRffXh
Ncwi1Bcg0rMH9NR1NOvI5j+AtgGgw0gv4pqjIUV05y7RygBQaZCEFEx1lRugiUxk
CZyrj9cPBqySV33UsRx/g9DLo4s0ORgLRIANAzavKQsc4R5S1i6sRM+mulYezbYl
VBpkQwaRRrtxs/oYgkUprAlJXLk7A9HReI+8Cwaqdec4hyKFRnL5JWxpc7MIDHx2
YhHEjFPteOYMG8nTXutKSrOLinURlravz9hEDc0tb3xFBdx2oQebYxJCPh3Nqzux
PWL4rT9IigfFczkxIyLk48kKewr1wstSYuDashrHH5MA+oGieZ/c05lAIEimalH5
nLuWZ2la5GZhuUtvAlFf+pS2ivO8jkMAj/Wu8lpE0sLKowfqB7Hqm2BsSGHroTGl
Z3myk3tpga0pXS6fjN1hGXx7uAWLbux7JvK4A3wStE59vAWvHG9WMAJgyCdOymcf
+4yDeD6rcH5UrR6RQkoSq5ZtqNyeHTLAwfbPJNxqbqPJzQ7O5RrgktmV3hCkcQTN
FLL8MEyYXkGoNUoXIDoph1AoL+EqTLOMTA56cf2K34I0CISnr/v4DwWwF4fvutfm
5WguqWewNnpf7OBXQ6J9AWwm5AfYhQMdM1zOaFKPzwaBbv3sRhH8eluWXmFNqQH+
oZ9QKatWrETI8Hu2HSsc+D5IAss3BMV19+94vXid68CAf6Mf5YCRj72CeCRAzVz5
EpdKaOKoTsU3etAE+c5AMOy1QSOdcYRAbsro5tedeN3jf6Xr7fR9MFsOn5Kfny4z
kUmDRxR9P83/VyW7dUc8hyVhDDxlnje87URFNPCjW3lDunID6noqxQQRNh/yU9PG
Fs21iANNimeIvok3fKgh9PB+7PH0i6d8hFzTq3x+EqKk1tHDUF2fF3YW4pH+BMI5
cRzOg52nFhxIA0UFBykD5+RAVVcaUaJmsCjZVAdfP+aBwoYybhpxeveK7RCB/C27
T8QBiJppIHSOzJ6ZeS4bjMrUM6lV2KAlzjqbREvvm8vDKZ/Dc0dNScWCaaUFS42w
IJaVH8PL/VfBo1AEuTvD6+DHD9N5ftKFsVdI/aKFPe+FoaO7cutSVNv80KW9oRxd
uXZunUgYmt65jZgOFjuKuzmEeR8zZ7wMzH2VlNHFCJeBLwNQzq9j5tBbpxM7tj83
6w2KGClbG4NX3nwOwCfyr/roZQEwL79ECdaou0UAVwM3ItGUwZwF4o89N0mI44Bw
Aglzv5juuvodKyVVay2+wz61+VvLzJY96YblFlAYQAOVx8I0aKoTTpryJUdgsEPA
34P2rKl2VS2yJnMic5xYeOFhsuZ9WxwzkX6/79SiSJ+LYdMyulPx+OdZAt2tFLGd
Qc/NxQAvcuSCQQbZu0UWNk66tjYZXPi6IOqVU8ZcmhsH9ySYaJZriq54QpQHwIUf
FE/LRsT+XdEEi5HF/yEmoUkYqMLMFjkhfbUXFCWQFLM5GQSPxkiXhhZgovMZcRaL
GPYWnpKtbCqYWvq0/bdXwnp/jrRxQPHZBrEjP1QHLCxYc/JD5YiPQf8Weyuu1LXP
UDMzPEkK58qrn3LxheQxZp5CR6jINKzfh+WU901nYO52G0bzvkyUvazomB9ocDTZ
R3HGH4zr1L99G0ce6PZ2K5jx9fqJ6E/a6nfgJT6unlvqQoMrNFGoKOms3KEJFTFy
zz4s4MJtP2M5AY9kUrl1/Y7vQwwnxzz0rAvCtmLyhO8MwUb2BjBrI/vT8pWc2Nal
OCCA5naY2TV4ZfN0QYe3f7bG/Ikhwgi2mX1bvXlp8zpwLqhPhU4ue08WerjYlh/Q
9Jj92N/cvbh9e1zKMJ235raAYnemzyQE38sgPc2N/xotNKBblzzYKXbr7Q4ygW57
5MqgEIJx8+vKPD+v8c1gfCxGBruoVmRv9GNlD7gE3E5PMGRxeUmAlurljEXmEqL3
OZ9WGCHfB/t0eQjCLs8ccv2U3Yh7QKOR/wkjOKxVbR7gF22jk9YoJvWFH6iX1VhJ
HfaOlRvoR6b6+BJPiwJzWEhLiZ+Cm4Kh8e4gyc4Fe1zgoBwbcXJqZ0Xoj8Op7wNi
zO4ylHsQdjK15tRGwV/Uj59JYTeLjcSBq7DrhoxeYFcvcF6er9qfPILRTzzxFlns
Me1Hb6J5cYlCqdypIs7JxaM5DFFhWiwufbDKFPkh3+lKKNQIKbgSzuKl8zuf6dFY
ynLCmp7GpkaQ5yabNNMWvdSVR7FQwNGz6DViSgPbgqFn+icWIn9rMB2dNDx4Mn3x
+MQASVPBcpK8o250z1xh/tqNZyRKS3qJ/vWWtO5+OGWTGIhQ/zPkwklpm3LE2Unb
uZq/Q29gaAhXE3Tn2GbLm8BmYUwc4oMty3QJ0OCu8oWsy67ShzbAxsAj7TO4NijO
Zhgx5KsK+s24RvoBgGq1xBZSQYwf8HdZIqoTHq/s7YSkn747HWSUfccyEWKkUkWs
KO1y3pW2xkmxx/yPZ820GLf0yKNg6tKYVHb0vpfh4I2s1UuDbQ7/x3E5WT5TZQPe
PI51yvwjAA1wj1TQtf7DNgP+sktgczRLpJWmlGxq0w9tePVSbRRrzs1klpcbM+KE
GzKLofnbv/fS9yOJy8DUfxfOxWQy1cN2T+HKaY+07IP1NR678vTrI8AwLqRP3l1l
+lUT5cBEhuMrJbMUhiG58zQuSvosNUmeVGGjdi45SwZGai+Ri7Ho9f5/TjTfQTZX
ex90wEq0MtKoB+z5dYwlKlZQXGt1ONTek1X9Y7JXdtFSbx1nKSBoDTckEiG8Unlt
cTAKVxode6eVO3hUUPnLeqyvRfdUmKwthuNOF3cTJznDxmERUw339H1RNoxbAMTM
8/MqD6SIQ7JsCNgTzhlWqtGNDzsYRDu6oGt7VOGjOAWGrMqZB8IEm6ZY8S3Cisin
QHl9tisQGDAtefT+HAT2ONIqFDXMWDi5bO0YQnPp6zR2Ficg+Ajr+TQ2LQPLoKym
UzfUKiCunj8qYvXh4RvclLsYKnjjRqQoe96LLC8idBEhhwJacp7KTzZSmf+az/3n
hBejUGAGtCcCPwKbpgpsQ75dPWgXiFhejot+qA9MRVJkQ0pB8EUR/820iVafCT4w
Xq//lAphFeFurKN/0lX5qNM/WpstncVvAgWkJrCrL/LigT9wxU/rRRZjbLzK2KUA
mkQAZLNCQpXHRRXGmZeoCcA9/2FUmTbbvEmVxPUYSRRBuNoa9tinWgnb4jt5dHku
Qkfkjh99AAbgFuLLwFSHCfrdG6OlltElvuDW0sPwPuduli2N/ZM1y4kiKwVDQW+D
WK3HplN2re6lDHqiC0pRAWdxpkT+PbwSpp0T06rZwYGYKmhX0Lcd8qgFnH1iITdE
eHWfWrbmcYHfQoZA1XqPRtQNqN5sRieIE67Vd9zywmF7Yy+cF56QVDsq8/CuzqLW
ukQyhkR2DV0aUSCQEt6roee3xIU4hq4yU6wyMaBgAkhPymTIkay8TTdl5ScpQYwx
IS8FqQ0nvVflCfJpSiVY3kqVKVift5XH+DlGQki8/HOmzMH9tTd07fmGbuh6Q4vW
eLyoc2ccEM5TrUIhYCB9WBmflBlC9SMrvrNEijXVKC+oNTSelF9NFZS6zLSZUSkP
2hAnd8xdO5kGB6G+ZvZvNi92Add/NsMz+x8ZT4aPv3pwO/dEyPdOHtcZFa8I/fLN
nsIiBJXuF1lG6qLeG0cZSaKEwlKOvti2hJBTjh6KsZt4TyuRnuwVdb6b9juekGJF
3loBJzCjPRB4ne2hu8u7axkeyZY1QsPb45bBKyoOWWZtwmnrNyIbw638DphCd9Ze
lDfQJedazkHFIM4fKaEsVrvn7AujFkLIM1OfkVVVOG4a/h2cBDAb7ZGeCsn6jZmG
qSi6morG4pGUVahzLW0eb0ZhpSOa4n4lHkyjYt01R2337g16F8tZSE/HRJmyNmV2
YQ/CTtZClB6IEcJ7zSF4iprXur7gAVSy+MGisdhbdlJNftWP501DD6RaAxBNi8l0
KkcdZhpNwo8mXOJ6+k6W4UM56EyXco1rO73Buelo3og7Pdxx0QfCE8b50I0V4xk7
yUNcjkEZQwiVDbxrTUlswjwj8R4f1MSnOkDg63d7n6eSHirunzeC7OsnvBVOq01Z
+QA5QZZjUPIUroBt3IJJWEahqFsuCvH6FVE+Z2EMGEB/RT49RUkl87hpOCMLIPpF
u6yuj9OsgQ7Gaxnd8ptWXUaefK5gvyt4XvAv9PmOtW4ydecnvlRzyDh/cM6FqLsR
kVP4/D+OKujTmPJq6JyAHWLiDN3qjURcIJJ+7GEBbhAwHGWwsxW9sjIo1ZJbgFem
KJgG8gbO/NpuJrr59fJv6GMZ5R+HG16YCtLGcPzyhdTJmcZAZ9xvcwZO5Rk2xCuS
d0V9ItA4WTwHZk2M++AxezFi0X4YiNpQ8BEiLlEQpKMCQF09oUz6kG8Jh+HxCMIs
w+c+S4gsom/aAzyYgr01qnb1HpChLwwgW7dfMyws5R0L+9IOjCYn3eM9uUlXrVOu
K+L0lvTDgzEiA6vPo4bxxikk/gKU/SBenhSGXt1nTG2A4lxacS1sOkNhYQX+p/QQ
yMNbRrh5SizZ/XLJ65jyjACTHKiyOxrsjyrE4WvSgXvzDOYeGR1aZr3WwZRzH8bU
F7ooG3orQqLoGR/52g5mYXiS3jpzorBH6kJ/UJA1mxG1SIRqo3Qj+R7AbPb7uBUe
ngebrvCnWcNmWjNvedRFZCMOWUuZh1+yu5lnHTwmXf8fR9TS8Ils1ZsjM6fcyWTi
R3eqZ/Tv/gFvnmcG9V4PinmYAGPHJ7hsOZRD3NiqMIvMIZxu+lEQmoOPabDXYRQx
QQJCr5YTG2SdSiwz7IZmcSiGeOiFZtoiJng7p40qFCBevVp2YsMFD6zDbUDojE4A
LVOpThFfL/zfUbjkYvH+ISngoy9+5Ydx1SjS9wMLVdbmelncWBH1dSS6u1zKyiXt
Bua9VDoueECXCn9Pvo3qkVPSjaCUr6QxY9Fr4DmTYbOR8wIODo3mISGYp3tQBV9T
j3y3RAub037stht9A/1+fqB05v9bbKQnZJS5CR28CHPZERAv5qIzSeFdexngsqyh
xvLdG0qquO5EXSRhGoJk9SarSJXwDegXYqgK7gIlhDb0pMXtBioOtIKCSoX8E1tP
hmKeY2afMND8RFgzOoq2DvWMIQnoUeTKp8cvO9c1PMdFcp0YP9sXIM2aFWl2sWAP
CV0kMZvWDBBSvKglYwrgWZXq2ifpKQTWu8+y6XWLJIJJBEew/TqsnBpvki45d1Li
238Sf8EcBvck2hvsrhfEH9W7Ldr4p6AHejf3L0wxuSYWl3wS86HnLJNMF1WfyGKH
gZ/WpXfStO6w+qbfhXfUs33nhY8/cLTUYkKEmyU2TicNOQefDN38PithOkRoE/WB
XUDPWJq6OIjhC2WdNonY7C4zd+rdb1aW3h095nq4Dx81XgWDqIH0y+I5at9cCliv
2NjJ09TxENZjSkmGckmFnydicHKfcOU40xHMs5duIcAH6kwFWtCFa3uAwQYCpDVn
e/ctPKqmuL82HanGaMGGXp/D11BYhhJqsDn4pFyYsdUQWhPo8h0koR8bAwKb3NAh
4B4g7CU2jpm6QmiJBLUbusiZ46yVril6fxaNYpXpDDJ0hfMPzQsbWmgw0Ng4zQSa
hoEsp2EJ7VU6UNfuWFNbZcj40hAWb+cxNnM9h7ihcvtkyrRTkZQXqclbAS+D2H2c
0ArD5ti3jtqO0mcIo7eHrtX2ObqEQ33eeL3SQRyl0rjrQq+uRJm0ePqNJWM/Pegj
ygHay9FewrEtDxHLOb/i22GXLtDLqUt9z8WN+GYPA+d3yKq6K48HywYSPqHreeGO
RJvHlezN++P7PqimWmMOa/FqTNUnRXydqQ6o060fjebIuoP/Bju5VfrHSGDOrPqj
Kg8L7xZvruni7RsPVlWI9nHSkrifDiu+N3xcNq6t6SuTvrj/KL5NWKFbOVeZC7j+
r9r/pDJJhNPS2bLdTlKVcBuX+iSueZxtV3w+kcuHbblhz0occKV4sR2s5qS1HJFK
EgYEhxcNWZbwV7qSMYBlCEeQtwJm5tFHmFWuJNR2O4msw7Q9CHEQs/SgHQIqhDB6
uop28+9HTZDby7D/a02sbmkaALxi8EVKWhsxlV9XDuF79dmfkZymn531YcwcbwIZ
vMb9Oo4p+qivgkXh+5O4q5WPpVZwoqQENR1PTZNuIYlbM2onYPV95T95DWNY+FNJ
KfIKbrUDQ7ZdTGim+Fjkt9AhQlsNS1le8f46uQs3xRFTo9F58b+yyGoL+MI+lbw9
/BOxPTdKknpFrSbJc7xE2D461s29LucB9O5M1tdtAiRBzm+c9g6GW4w8yDRPi/vL
OQ9iWqsj1EYWS5rG3m/gmcbwh8uHcb6+NlYGUYPRQ+1ykBe8HlHWhT4mZAteKR8g
M8gIYPyoo50V78dyXM00JKIMaIlLWZukzgHexQsNv4R8h3td1siYafQsUatp/yVa
lxoU3aZI2dBSlLGLOyumUREcI18OG4h7L+xRkeLw5h4uzdqcfEFN4Xks5xyVWdt/
SPIzGJnUbg2UTqAjUsPMnS7wXsSHxhRzmzMtUJovgSDC7YceDgAYfyz7iPdbRURE
rfyrVYqyqIjTEHHpYv7C3S64FRDsTnAsijsvwDY7UBeM/BADMYX9FknBqjapSCes
HaufE7HonBzcja7ejwi5I+RNyjgAtQz0mo//rP9liutH6AJvKP0dPFvZBQ68zfbU
37u9367MesZwgDh7qtUODTsCu83TWSztmOEg8Gd3TSKxMTzhycILoi+chV0iWPCV
lwZpVR5N6wM+pl048HCpjG3piOE/IMVzIwXNAkUKsgGhCoIBjJFcIm0z44TBr5qy
KvwMpCotO9GmL9qV2SrAaALinprXfE6pZGZhtbeENDmY63/7Cee43ikuzHy5GK13
lOiTfCaMchwGhACJ2OPmo9O48TFuVogYI+zCH4IrDPtzUV+ErFQAym9+wqL7Izia
WFqW39HiITvkRGIZBUx7MyGONLF2RpjRmwLGkvVMyYjVQ9CIS5c+KkNQZylt/sl0
6pS78i6kU0gN9Sksw0s+WQikZHN6sey3mKgIsbG/GEg3ew3fMBypi1v89KDrJCs/
PhUCZAgVzHJg0wPc4NUBviNwd2DYIBlht4LSkAjqVApSMiFqX2YuSmZltG1kOQac
WmzHDyNysBWMCN88C/hY+urVog2/cMiIULufMsxsmpDzxzwmJw1GfSOz1ewGpf73
MFFZM2VnSjdXCxQdmNIAG9mnThg4KiHxKsQPLhjwERNrdyffh3tI/mfeQQfV1VuQ
clFLvt1xCvnSxZoioatiLaOMSUddIQjKln3kDYMewxXluzkSEOsQQF7JYUNFSj59
g3HBtXe44rsoyIVhRQbcAgTGIMxJInGC12JbowdM39IGr6a8Cn1SHG5ma7yU3wEu
Sb5fT3xUefMXFu5nIo1We8J/P9bX4YTPO/tHkAIRL2pziuMgwq+pUDikSDQp8cQ8
Sz8YYmcaF9ZDWUcOuU+F/JQqXugjhiaIoensq55ObzvSPUB3QEEf6dH4vBAuCicV
C+VGgpS1iBNxUJmkR4935N+GQ4IW2gT27dHfIP5LmG5C2ancejBDXBCsgQix9tws
E04K2a5mubjofeQ39fvJKEaOsqosafqjMjvrL2gxu3n69de3y3YLywRLZCb987Oa
MyRiAwote+Q77icbhcrf2Qvpc189Tb+06htoGfCHOkYIenYp/RdQ12JdgzSP9fqU
Z0Q9wXdcdFOz0wahkH5NO9KmN9lbkWi4uRuLzuPqYe97vYreLIktU/NETcotaZkZ
cJr1TVLUSroj7IyTmjtETFy9uaHnI/w08njClgUO2bnHSwmiCy7WQ/rZ75XM1828
WHk9gNPGdj6v7MAsGillnkt9jIrQBe+yGbdUOpETjgF3L1ZGdMMw93tB+c2f9lAR
6jQP1n+t2ya2Wn2/Fez268IhtVOy1DGPJtTRCycPOhUUyKo2shfJ5Y+a7BTmAFAB
tQf3RUGk8lCZOcnSiPSvbltoTDJ8vax74665SQgUXj6TFMR+pGYVpG4vCDDkR38l
sg00OMYpXTlG3NLOFTKHNBJppm/0S4ssNZ7r019WPWxNS/jGZBaLuJFM9vvwKNRx
/aZPDAfKRyufNekJtWJu1RjZAtcdydXQKZBly0QzyDvXSg7mH8Cdn+zp3QLrR+H2
OegJkoB4QStVdzrNkKB0gTH7Mv/OHhYkk1WXO30sWNYvyu3EKYRcQ1zq1yCPCgwy
nWVLP3O84005+wI1oBYcuJ+jfJydx7hgNfCtWCeEvmhff5PSqe4BZ7/7JMeFIDjx
aA260fBMZ+21ieguhXi0SmFtvpMjXCxBTAS4+g015j+Pk2u7L6Uj0xwzQB0gWEWb
1ZdWaBLzhHlqQQAw7FclEloaeEdVPd+p+GDkK+4DPXVz4b2J5lwRFpQeKDhUks/l
nmxh2B+Tzxieg2X24XLRn1h7K6zMfncOS8wrC8MksuSHdCL3vKmCrHj9h2s18rWG
HuFFjsTuXCgzTswgxdNwC3BQEBpLkhTfy0iMxZ4vJiEKQmPX0REpcfPTJ5QZ0hJu
E5qMBHaagdp3hrm/c+GFYkkSTloK7TNfpA8gUS+m4Ypn7mDfwA9L4Zq6PEs37jyg
n8V3+kbFfPaKUyt5PzyOSPLB1bTaHcLRQZtilZ1/EPrtY2Lx/cHnMfbwjAk75d/7
Be0rNZ/prKBtvW/h4sJaQylrMJGe4+OC+LqIAlOH0kbMC/v19WVEExOOxAuZlXXw
kaaQ1UryETLWUVS95xkZApcrBzyUDzlj84mJ0XbcHPyaYV+PtxAhIS6LMB7FSe7S
RTvinfFvBQ3uaTlYiCjJoc3LIzXDjhklpcGloFWRRK6g9uQVR2wFoQREeoBZui01
NiHptLbtPLh3IBrvDBRWN/eHhtudlUlre8Tc72lt7ccTgoN1ceFKHYV+DsD5ySOx
jl4NLufM+iaHqInFzjWIgOkFa636DQXf+skbQfq1d0oXc9ELCp0wYMPTeCHioT74
LOOwj/Xx44F1DeiCNSKV/L2EqU3MPVHe6a4Bz9nDAKwybhr8PAjBIf4sru41fdAQ
c6q4DXIyennh0a5PEpuDyt7oc4saDzd17zl86x3NNP7t2O6tItAHnfn2AatUCUb3
6hE4A7iQcSBm1D9/LXhh/FBaijrizlDSVshAiIDHrXb/4XZCUnKzepX2XCa3T3cq
etXKq2LwiaoFoAfRVefw/yIRJU8D2OFKqd9mKa+LaTfv+m33FXz6K8E/sq2wlwe1
x9bR61xSavC8foR78SQmjUzlrgrU4YgQ4V56l5KqqcuKOc3/aMR+V+tSf8ZJegHU
O+qrly+5wqRr0tDRqARACUQzYmwuag30ZqV+ysvP293qXxCW4+H0aWc9Vupzn+Mz
x7Lr+VUQEZKqbBZ8Yu2Uu1M+LC1Bkd2j+dyQsylUo1kW7RHuKZXxEqDBHPYAmLEi
0wEh5nyH23LevliNspIIy+tE9ao+7N/Bj4JbxtEA53lMKOLltiFJs78zo/H84nEQ
cxWmwCWb/uuPSqBSD+3fD+MbWuXD2304QvteFE6Qv9HXf/HUvqP7+7ytaqpSb084
GvwuuoROjfbIALCK8ZYt44amdONTojO1NaxLTjvAbnmdBAR9pEqWorAknabvzApM
RYuntJzAMFhcHgFPVgPmsT1xR8LrgtfHd53GFr++/KdYVdW99iJv0VcbpTONJMy5
gXUm6V3b0LFmE53klMC/bOb+XK6LtF7f5nH8TrTgP2b3SNFYn9MgAuaMUvm6mjwI
8cGOeG7bJkwCGIr6HfP+Jva4fSefk5lEKh7DK/h7u24vZVNyNHxCLoRImdNZnBqq
OT7rRoRJWM82/Pqv3lw9igHznKQu4TRP1kJlwwvyj61hFxaTC+RQCOeleL+fQqI8
dqsIxuBTlSpVWN0qYemu/1C1+RnwxtM2G1tdgDgrlOyrueu/Co2J5Ydq8ikQIXtJ
BYWY4jAgrRIhtO3UA0hlOEwWeCukHBU8GwWM2jBVXIP9vhkMygg2rS0S8J3yLRdP
mHQDBSR4M/HIJcqp9H1pY4MRuhaCqnbUWiqWZO8nGVpLKP++AwMivBv1eG13uzVw
guYnQlhBrGoIhewgXU9wl60M9hzauKogh0m750dawajTCSbAikCyjrPIweFhDGFr
A/aM6HEuZKhchELrBvGi2nkyt1OQyyp0IMLFMOYTCzx+H3I0OiG2cZHTenA0EetC
GGfZAm3n3W1KFJFdwMDN2PqX7KLwLIRQFQhIZupgoBByX+vPfINFhOpNnXSfKA5i
+IpLqoSREj3xuxqGzk1vxETI17HFKaWD4BER+W+O5AIcyrV9PJjVagAECWH5J8NR
l/c7T0SEOcJbpUBLeJmWNicfzfr/092kd17Gmv2O5OGrqW+a1DlBg9mIKbAiOv5n
jtdCUT6i+gN40Q64z30bibyIjDOQDimy5Xpvq6XF7gCUHEqbrsPbCDK95dpLfom0
aXmSt2UwaFzqUBD9dl2KzD9b4GtVTNJGtG9B/V2fLiQMRYe3Z0usq1ZV5hQU60Hh
th3QeeedXWwiGgMXdcWIygDMFPTmzr6bMCThV1x6JdWtHUoReqsoMuUeYaoBPbCH
N9st4jqCcq/vpA2sDPVMnSuZPIGxn/PcL7PceKxesYJd8fAWKE5AXpWwbIMhRdRF
UxtrSQUW3RxYJlQn+hWBMxfth+2lc2JcVpNhqeG/hh2Ajn0K6NmtqkHk6DW8e0ao
abxVTy/hWFbdjTAwvciYSSTK+cnndzlJqBaUnCXvbyact/GK9vRZLuuKALivPziT
jtY29KCuk2mjr2U1au4rvT5Ym61OxJVJKiGlHHUGXHcUEqonlxAOnaxSREu/9tmU
AnBJooVPk1fLstSOSeyl7nOvY/+ueV3SEQW0qwQ7s4/xHsYZZLTgRLW0gbjAyVJZ
SHDsn1fCv9lMlldbEHfbwd4MfbRXGEZrTTrIxwb0D+cfBEr9EoF0sO3YfWVHMCVl
6sMx3rx+tEA4VZxpyfDneBcc4GtP7PGRw2Qy10XQThSYOB5c9jvVYRWtcEdEPd6s
WKPpF/E4sdT/3y8c5VUgnV/NuISZgu4kv9G2dPelKFocg8jGwKBpT26dyBdsw6mr
8Q3F/mDYt7laIVm5heJK+7IcHkl4T2xQJAtP9m3Cmu7sGWdZ0Jj/xMsBLBDh7I6D
mzbPd4VNGyY+rvHgpMiTtssCuD/pAPS1O2RQ6CT66MU2Un58s48IlyflCZay0voU
fReMiGlS1RYUAQzpwDFLUi/xqz17ANJd3EljxMhMXlsLipkIw16tbVpHdneYG9dS
WhzLHnZ6e2ewucfSmgXgWWbv3pASNghQmIrGjx9sVGyPSRvBaVazJLdadh+s05cn
saJsHmjztXMQGRMlf0BIOJmGYf3OT4j+QrkETGEP1GiI2H6GWEn45weqh8NuK5bm
nwH2AhxarkOL7C5v/KS2U8xYsxOOtB4YW6A691lVkAqQ/FIo+5FDsWwm1DMJ5KJn
b289acQriTp1kum4HbK6+3i40Ro1eM5JKR/NA+r3hfXwuxZ3BC7viMCxlFE/IMIU
cOUz62mcISJavmeFkMhdc0NQ3fhyO3QSbBwnDES6xyBxc3Sm+EyKxxGSRHq5bYv7
okvBoeU8iqoaWkgpkvZCYD03mFuN4wWcjtJIGf7XK4MacW33dX2Ps9y6d7XW2pzP
38Ktox95WCySw8RKES5+t6ZDkHVqMKCXle+Gg1O2Tsdc1LxTPGnhhTJE/BxDgpFl
I2ZupoamskPeYoE7fiZTQioVDJzEPCxV7Kw3YPvf7/A71EJxbjF2DY/EcbnULSCZ
tj6R04u6cFsEMKBEVaehhk5IffynUQN4wSCgYUjfJxjzu66GFr7sjzhPhVtGfdYV
KL3hHVo0AswTTVVb7PaaT2KiO0OZyKdTsyjWRwUlyHTEJm+vnZBYDv+9nCJtzELi
sBoqsbtRUZINdPakdpxv6TH4PO5rem7d5nY5axHZjyawsyahFNgaHEhIOK8XrD/d
YGqL2u9UnEUd+7126lC5YS97hZetkUzwuJZ+FfbPIo2EJRk42JzI83MXfQr6gIDu
K7fDcZoGUSLnZluRrhq+Nx7E96OPqYHCvFsq+OwTE+hus1cAgZokaLENOIpf6lrz
UofHTs0omPGmJyLP0cytOaoApqvS67VTD6/YaiT/VT5lCOHbtrrqqXH0dR+381mm
DNliwxN1/OmqjpOQnwTrh0/NmEfeb0yhWo8NUFxrK0dk2y67KFvvxSKXxRAQwS/j
rE1seMshjW5JqazI+7/KrXa7+Xa97arPz4auxCXBt75JQFeR/+8NTZVm5L8JKfEu
LZa3iSOLb+E2Xpszxgh5XkhJ7OBGhftruIXxFj/Lj6UWeYoaQeFNTcCyIlmigTiZ
Utlg/2OFcoa9jXOghj4LN5ycAlC0wx7d188Yvcr/kAr3dGoV0SqjRdSdO7aW3glY
B6URcWO7NH0zzCSv3cmSxPZ/LVHgFbA14KAv9iU3W9f5XpuSY89pwI94ai8lNKGc
assD4HpFIL8olDNK1bPd4Zd2yF1pRyrEkmzl4jw3j/eq8OPu+gFzF9ybjd73v0F5
RHbcAssvYOFTEDBhJRGc4RgxyN2NsmNxG9SdF8vAjNw8WIGPiIDA6GAkul8u7eCB
Zo8XN4UARyt33lH8Emcja8Q2Kutu51iltVJN0r4zxUN55Hzp6ijN9PH+at4bOkAP
lBbLQbRCa6p4/R8ZpN3y/E6QwCKH326btmkwcoTZ2H14Zzxb/FfGdnxi+Dz3mva7
+PQJ7mFbDX8BJDxcoo2Xe4ren7zjKzbJPsPs66EjTWOq+JeX9LQ/cBmGSnIQm9QG
//ZS8R/0kQtEbuLUJ8Rvs1YH8XMIh66LhQyFeyZ4o0pe8mGldxBDjmXXnkDwnlJc
f4FOEh1l7t7aB2hHbNkehcogrolsRZdBVuwh3cTFauJE15e2lzH4ubhNhtGubew/
s+ibEUFO4IOSmx1bwkXPURmkjDcfW/ttMpVkYo0wJZY13wXRFiOB51TrBV+Skqgy
ntTQzbDRLHsUVvnHbClyn+MvLPKNQJgdDPx91YTDfOJT0NByQszotwwBcXhVrM3X
R+RzMigU0MUmdp+gu1D+qsfIRuiw4YA06p0raLBWH8WdaIyK2BN1Cu60EF8Ll2Lx
4QR7mOp9aainSnMVsauCKx03kNtJ/YFUi/aKZdlxRoy4CSIuYM10oELCEG5jIEtT
htqophdwNWM1opBVaTn0ROeKpafsFFySqq+ztar/VzP9mN3aACgmJuwER4EFVxqZ
YUF/suG4zodvCspQj290OVuzq/UQst2EY6NR/HELY6P08dB5odbKLz0YQtPFO/dd
srd9NpJvY+ClwLttq4VnOn+u1yHAtmh1Ig6neo5NcampPZZWZGjOW9U8sYVmCinA
ezBqViZC8czoS5HdZarRKlKqw7518j92S+UGQ0TFLoU63ir27xArprM6NBYgx+do
Jb5WYbP5d3pDeZORILdL5UtgEwvCoOY/1ZfYL6JRg8jF6x+xvElzZHNPAZ31zO3d
sQb/MVRfPbFCNOOaDWZ0MrwevYf6bE/qPy/JBNB4xyimbNmnt5QNoe+rmelPakVU
Pbshb9DIvdtiW/7B//YlHXF+jzmFuXxdB+adremxweG3kxSpS0JO42DRf5kryQOc
TZqQaneSsbE+5bztsbJ4m0wY5zLXilCjm/fpTQ6SRKvkfndjfG+oebtp8eWYz4Hx
aBfFiHxyDVXuW4B+FDtWUkmRj0K+3x8eE0dKHjcu4k2yIoyckl5lkqJLuuc6HCsG
bLDcKfpJoEPrDvuaR055/NHLl93Cyj9rLToJXYt6cs9Q+XIuHwx2Ami7wbN3Gjlv
ONkm9giEQS+MqxbpBuiiY2wpcA84HrvJO560mvoO9pF/MkoF97ksJEZOupgEE+0m
XPpIDvI3mhB3/J4a13pMFbl4bn+xbBko/Y/uySd8LqoOKvo2tnEST1cxb/HffRhp
lRILbb7UtRKdhGhbinF0S+xWipn0hTJCQdYdSU0LC/t9HQHWvcJifkpZ7qfayEwO
5wmrHyctN4VX4xsZ27BhxcZP+7ibOzFI+yLM7QxpbEOPnH6LMfzt4AtsYXrJxTA7
YAGUzU8rZWSJC0d5tJ2txLg7N+tn9wRaiLP5R+rv6lNkzRj3OEp/MoNNunTC3Nq2
gpFajSaof3lpDyD3JE/6yBDhqIgoGY0CJ8B4eobCFUvPdTWaCQkJsJst/+CiV9lO
35Hb1yszrPAJf5kNGikudmGYiB16RxH/TriTAphC/ZQavQ+1ir5OU5zcOzDO+9sk
zme8ZJPjRsC6e7lJlWyxbtqWQRPcD+rkMrqECLynUSiL/45bR5tZZMV/jBabznEP
m5TVFGfQlFQVmkvGetK7P426jpj9uczrDW+dS4Blj4q+wrvv7b3cldWDfytY/vWw
+FIKnnG8UrMAvzECLYpFY1TTKtSyQDwOvqCc7iMXGolBq1SEnSIlQG42wS0W5Nir
v+7vXOkGYm6eVwfJTHxMfOf1dFTZ+PONwih8Npe+wGfXr0ZNyefP87JEnrrGuHgc
0mdhNf6WcGZo+5GHrl2FVoeBtX+JbDoIu2D72YxU4Yjks3hjb5LUr1c1Dp8+3Iei
5ieIsO9Qj7/yMgxR0rznAZz2b+nHBgEqxj6ZtRu/t/cd+pcKBeufeaXrgqOclF4j
io4BN78CZKGbYqf2Z0E4SM10lsOVPv21XPr8PzkSPgCT7Z0c6sau36g2GFNVuKzT
f1OQ1BfcUfl6boOepSLWjyK10zmyjygqYrD9V3yEftJEo+flFMP7XwjJAAs8QOqe
DLVBi8sMMYeAllgzAfLuj5Zdn6+1V9QB5/per5Qm2SP/nFMAn0DpfxjbD/Jc4Vfd
GL+skkzSwVGspCu54RFJxWCkrOQQCGIT3HM+gxyXOR66U5Q5xVJ4NDY4j6QiXHNc
Td+eu/liAlUKmNbTrbfxb3g2rlduSGoq/kBkq/nfO5N7wxX05QvsXF2u7bXePtWa
7pkjE+S/k2KFZ27h3h4YuC9DuU9UrUuGEvJkpjTzrFYKVdue6znPBHAfB5oc02MO
FdgE/NaMt3tN7U0k3Zv4TRJgjtGmIOOzriTYNCiiypdTC73QIFsQ/J00yvtH3RLq
xGYLBwnAoG5alhsL3oQGGY69JVqBkhFs5QpA9dysoZs1E8xQXljoXcuMu1gzw/C6
rwUlhG1nfuFVvif0+3RE9ud7QihY3QVXVNv+/4DS00XAn3QIHmyVah3TOaWMrCml
UuDKpO+0E3fbfhaigLSF2Z5/HxNepIaJunoVaqEi72mUhFwhGcTu8LV8tJDadzF+
UEdp34pLDMMTjxdyq+aLA/qZ5GMqQ8ouwWXoW4kvexrWu/2DHBLjVkJqmSd2ziUD
yB+F5romEvMWd2HXTDYg3VYKLJRWGIPj0cuLVU3TjNLeiok9yC8fD+48UKyXeedQ
WPXzWwaoNsVDHOkVgxJiWGs955TMPGwavovzcWQigp85GIjgcX+yuSwqqWGF4o18
/riPETuIpsHK1NV2eB8el76+jl+IlAfqAb0/+XZ86vOI409rT4jfsA5wwxpmkT7g
OQl8aG66dVsWrVqQCrpmd8c32KqJnx5O4Y1wDBEg4Cl443wVY78EIWXgVagpX9uO
licY5maYsrjZkXivoJaenP3b7BymrzM2FGlmqg0I76T6DhDSz7wLVFmC74QA7AOg
AlbqwkYEQSPJWAN3D//zWBF0T17rgHh5WKyTObhrOpp81eV5phww2BwDp2u8glna
iLDiiSFz1tXNTXg/NPPcSthSY5ArTkXU0BeX8bNkICOK7STATyXJg/T5t3gb0J/5
t+p2/ZA6zfuoqxL+1+xD6vdk5MFXDSW+K/5SX4JfHPwcTHnmoZEctN8VtO0SXkTr
NaWmjkheVhAjdjYYknEAsEsdOv4gQW3b9QcTQGGF5W9E0ZknUgwWwHD1QCT2g4YT
P40ay8AkFT1npHuP3kCe+wyuGN0KEEtmKHgieRHlWSDdve1VtvHbXerMWSH89Dtv
YrRFMPI66dGpy6yxwEBBrJQX1fKkDqC0RDxJ/O+YFS9/ZybP8ukmoTJoM2uZwmCz
aiWTPBnkiH/s5pZ5jjlKOwTO/4YEyERHJ0DiUuiT6VPAQwctom6b65jvQgfwU3NT
C5pC7FjQ6IRJYly9HrWTXU0waiIm74tnTdSnbn9FsrrYgz7W2f1rEfKsj/nsY9MQ
7IeDQgraayiOTdZ1LPgMKpqY6LxqyEMRPLuPfTKorIsgb1u8HHWyu1eOSKiHaAfB
59Sz0w0HnLQRbclqRHbWJW4f03rw/ovbT+2kI0HDe3ySaT9HjOgXyhZf4B62dWvT
kRytZFFmwQUg2+FcgiTDBu6jEA1YRAOqYg9ENfK2HTqEn33TxE2MbkluiIDkkh78
az59Uj7E+ermLx0kSNL4iSjOtbVcMOTtAFG9W147T2c6LrGm6FuGtrTtAEWwiPsp
OAAPurVhKe4xUP1+Q0IDo3dKRrvZCcKodS7XdZYDvLIOIG3BH7JfKqkRpkD4cmeK
mCuy87yMN1EA7DR2ZljNwGrZbcDPdx8hScIHiDuC1NF2deOzpvcTAvsjxsfgXRlW
MRttYWFmKdKuvKLJfde2rmaL2I5quhMHcOGH/hA/YY3y94pcf9sqNDnedeXSJ8Hc
R3csoc6GOz3EEQVFAc1v7t9La8hFzAhuDJnrGBoia3cBmRa2qElhrQ9e5bO9xBZx
rjkHodygqoO30hSbJXzOIJxtdMcIUnka1pTSL/9pn5QGNZHy20N9Y24Za2JaQqFr
qjBYscIqUlSDjJB6n9Wde9PFZ2aFTRjgEDqu4GcdrsWeKBX8R+tn/WtfoOT4D5w1
2IzAtvAFAtLG/VQ0DxCyTpN5Vp8h8al149TbBbW55U/pHZNk7yTzVdhb8VwfTU6g
RyBHBwnZLvOJtzzEWf69h6fuqtgDuSQA4e8WOggxQzxGnQbQJy+N36FRGaer6Hpy
ChnGFxyAo+9Z2o6QTHEFSWJqY2tWtHzrCJ4/9oRWYDB9gK/JfciNWdOvLakQpZGO
K5Q2FI4VmzqPoFZXugI8hZ08omxAuwJIncgP1aN9BmSVTo/UbTlyteSAYBi0uYnX
bUDzWRZNkkeSRW6rXV1vFxbHUwe21h0H56gww7rcviTHy9aBJtShxsAb0v9DgsXR
iV5wIScFb3yEzsGr1LHZBt8KnqHBPlzYqCt4/pi0hdijsbjP9RDYZmAZJC/nDuy+
djOL6x9hs9lcM8luxVm01lnQRbU7tVrFLxz+/569hoID2qc5HYUAlTXLj3e44dYC
CNceCK6WeK6KfCgSYaE8il5MfOLJC3bYcnG7Uk2vi2SnxF+znotNONawzrc+2V+a
kn4QtSxTzTdEUgHU75owRJ/boHzq3/1TPjnWXVeuwvqCgy34QRJ/SGxvF3WAubV0
9GlwmxMPtMj1QADHBvlddV5HVnCxQnC0INHIEU9yBHYamp0mgcPjb9XXnKshVs2i
62T3zhAaYGFe8nsHjWF1dvt6C8mntv3uDVCEA/5t6U7ZJv8UoJMNhzyb2vRycCZ5
nku5DQoxUqCu4WKrvY9JhsgE+LxvfsNcMfdRVNjtpgZHT5r5UhPmHQRhGrGo7P5G
8lMC42izOItobSZ6BwvJn1oVSY64dSoz8neYub09hul2mZ0AYPm6GJOjPVPru9+c
fgxj+TmYnQGxKewvH9CIk9x9IAClYSu2aFdnrPf2/oAfu57juhcLShoeV1efGriX
pu+vnDYxXrabtZTXyCZ1NMyKrX0/hHkksMF9J5PGUUfHgxifHxbhqd1qY5WjhWG2
NtyL2F+Lk+ULXcbgcdOr4/31MSHg9mpUQhNjzvbgV78cnahgNZdRp0z2Gt0S50sF
gVHZzFVatOlHKnI4A64NsrfuMFH/dpKUsLR9aalrzja1x8wiUUxCvEYCW32tenCL
s9nbiWxH3+jwhjQSj9KSBCAhmQMnnswH0jJfwpx/G/6+0YrRBEfGn8uCifCTJF4Z
Q7SLx7R7Pj/J04mTFZDXctqhQ1moIov8SFwqhH8wOeTx+E5upPXLbm/iy0kBcL5p
Eu+og5EUNW12X5JkIRF6n9My7dyfa1trXbQw58ahw+Dz9gq7Ul3+wC7UGCkQq+RG
l4YKx6lTgNgYf+mLulHYqlyN8qWkV7XRPMC7Jf0hBDgjikj/255fvOb7uoA+Tfbp
p4QsHo+HPw4skXPXqPpdt/JSZAxh+WxC0Z0nkM/yE4lf1J7g7HNlPHnrQmdX6nEu
PB7KvAJV6IKnPxHxG4LyMzPElYiXOWb9aUtWBe9ecw730XJAdCaoiN8vxGugi80z
s4JjD0vrBUck/vgJWGnnTYaTlg1pTilohRJ1BYNlPVmt2SQ3ntr4iRkm3ai/XRcj
ZStX1TTakSxrnlDYqPYjFX8DDG4bqX9hIyGacfor+lvztQBIWKMx02JFulh4lHYx
0nDSmrJA8AFc/wFqgP8fijUkACIK4NKKbbZt9kgvaeUTTvLTnZPFBARYXI2xUR95
4MOX9EMb74XzFja9BMV+rNzVrNAcFvhuk8ntzOStFhNp6nz6e95JjgO9qnZpESL8
6e2esF2riWV8MLRxRDnw+pA8lp93wY64DXTLk+m/G9BJ5sYymK94BE4MFsZ+xFm7
tzY7MhxobrVyyoZFtJOpWOHEsyQ8uC9uJgoL3LvZWRK6VRxSXjARueLMfryKvDDX
Lx/iRBxZPJjD54ZaZUB1RwLehWVfG796mR3ELgvxO4FQ/G1EAmaMvVjhFBPqWBlB
PvxT9GGWHdX3wVqjlakOyM8M7A5drCmUk7LO1ikI2W+yRKp29HD1fRQnHLqcL+kf
yx8122dW8lvTgZfUM50v996eBzAdDPzPujf8cT5BRGfjW1j30vRnHaiR78jn1Wf+
xMUqa5mbfyiflAg+VFzAxm2zK72b8i/hcH3Bm/iCqYoy7SlZwIE5H6v1ezWGHQC0
VxrtzdWDrJnxZXX9GuvjiKrh5yNvcry3apKoc2NHCtWwzUBTb85RV5ItZ5J0j1hH
eIq/QBoAd4daQqkb7a64Orh3iWGuILvkZmxumyGBZ9nIDd24b5Ngg5uUXP3IKVEH
IkkgKbIys4Rgcl7rS/w8KY9mIYhJvA6aWAHzHGae4YLYAyMpEG4GuONNp8bU7umu
feMWbxpQRAzkoqLktENJ3T9zAhzRwaUgQ374xOu2Goe4F43ZMp2cY6aF9u45ZdFK
CFjOiO4K5dQaVK0pmNqIMe194R821prj8vxi+RiHpR65RGByc0AmU7p2Ty4Hx5Hq
QhM+kQqjWhfRJc3NlGq5jqLk9wSXz1c1o2f5gOb+RNBgCUxxQernJtVfROeXxvWN
+vLyVdFGrhTJ8hKz/APadZknKB4wa9I1GhD0t6qQg6/GZ26Ph3NvTyZh3NPEaYyo
W2zS6mOtdB16II7wAf6CiKiXd8vIYrbwPTY5W2NBx37GNzP1ZSrbv+AupAiVNUWN
rQnDbrQ7YA3zcUuVrmNhc9yQnsptTU6ceLuzkuFKWPDSkEb5tmO0CKZU9PLZhCid
P/cRTc/P0qNr7d2rYJfqakmG2fodkpAO3rEOAbt+zVOgZPfVNyf8M8lzT3qbTeAP
Jorv6hR8ApIG8H3/x7wgy7EROIYfu4ji3HA2Jl/sKWb3atSMcTrYuA0VmbH2yZ43
sr++JHUaDWPJjb+bGxoAO8X4nnPOITqHpmdIxgh1NPCBwEnRhbfluwd7MIFIT/oK
CgX+vMU581PoBkLHzGe9gxkiMybw7ps5TLEF8K/9oYUc+0HeOCEJ7nuqHZBtBdzo
tIdNctoDUds2nkfiFGd/T0HBVZH78fSzHTxxs1XnHkguSxNFA7g+nfED/1Ys2Lms
4/0vLsPY6jnrglGgvmP9Sog6FIYabd2NY8GTcYLe+7lnbqCv+KUvWOfFACdqQpaY
bYbHpqsNoz5tF48TyamfeJspverRJnEhfB9HNrtLVnlNQZVk9MS15Lg+J7tsmpi3
xPBbrXEQXyJ+9lZmwJnMSRAvep/WGaTgZcaAe5LGAvuzpPQqqXKXLjeX+PAOhL5i
wP9Fdxqijllym4qt7q3u7/Kos8Apleb0l0BynB1+M9dEiMUIJAKRlz7DIZm3HBQa
6GghHt7aV/32ShLhTWPlfi6U9+guXBcfAumvHIll24habYujswREnRLzvHa9CFhK
4/UagNoI9YjRMX7At/ss4dokJxgREE6TZhVXIEVPL0hVRvEcUYncy9lXVh6lJFiA
0Vhzg5cP2aqD525tqeGHNI4UYlSFiUBZTyQ41u/X5MuqblLSN6j36u9Am1bsr+gD
ZyEqjusOHgCaEN3AH8mJ12Vh12x5kBUTrYZQ8tOl9aXxnR4uiQBoiu7WrOEQMZrc
5FWx/3DAVBRCkJrmQuXmXdBHvf52HrZUQBdO3CVw4AY2bJizbvE2zdK3QdF0x/ot
k5uwUZ4NL14NzXJAB3ykbV7xEh2aoCCOredqmTxPxw64a42KnCUq83OauD72erQx
vuLfKXeQORz5uxxQED8O0kDwBnKvG7lHZpogPXMZYcdaqVenknGJpb7hE2unrj3u
AmTC/99rqZAYw29VdbHgiCEHgTbjSOygUzLF1nUSyvKFId6KPmSO+Pg55m71ee/6
Ea8NfwFaLedPh3mdOEiDrLiClu063U/mmqVZqm6lEyfHk5xHeTHyPDElAgQYzsbV
lE1kE2LjAW/hDp6bmXC1qgXNQ9+23+Ks4/zudESFGLiv0ZXtMIyzIk2AjlhBF5Fg
A6l/1YpreM1CbhrjE2OAGUdFGCblAdQOmQuszRIN0xWkfpsUaXyz6NWOfdRPJeUe
cO9FY1S+RYvpddpfCSplLbxIqAZPAAuL7hvy4MGB6Vc5ZS8wet+YjtY7cvpunzbp
ji8I1UqyKLtrvxFNk+NltQPoeWXd8WCtAZ86MsQDBP8sghcx+vptSK+DtVaDA2V0
z07f9JlJB7AYneqHZQRXF4vP76LqGlB3rtrJGgL16L990vET54gBtckc+ygFsL2A
8/S9kHXvAEvySJtQl6j0NfichCgUrdo4xV43jrhF3NYBiUlWNps2rCwcNNvrTTwq
qk/2ulj+3E+rkT2H0lPemHz+EOuBk4ZzKg0M3qJqlJUysvk5RpqM//H66IokVKVA
QIfuuP+1abZFmMQJ9Q5TYhhGbmyaOuE99QKo8j78pewwolP8Gn31pZmGI+SthkAw
SCWhg5mMKR4UScLXhIHYnshVNJQh/aeSKg9x++MkLODIJNr/FDbRX5jp8YOiTjNV
TITNQCaG2I9J9iH9IlpqYIJDMwnqUDb4Ej0uW+DdYdt1mQdk0ZdLI3sSxiTqqlUN
1iohw9su5lmwRN77ocsGuO80z3QLh9lDkEezZESTSNjocUXvJogFdfzqAhF9ShZ7
WbCjqZDw+kzs+EMAb2zW/NAVGG5Q0ULubDxBTJoty5Tda+3uu6INd2wI7pLA3J8A
f9sx3y2YzF5zAnuOPvpbSLRJDHWwWVYHexNERuO4sEqRSIwNoib5VIRE7U9TGsQp
zPjWVnfybx4C0XVSAcQ7GXpEoUT4ml6+OJcWmt8zP+cXUy0fetFIuiSim2gIvDzY
CUM3CzNS3YIs0ySILqVOnCknowCz/2Tf9yeTs9vYS/vEb3Qebm+5s/DLxTp6EOjN
R0XlCs9wQ0invfuAWyy+5kE0edx4uqjM7mPzjtUMQdylizFzQ4KHm6JpJIiOD6uD
GLkASoMWaxoxb6n4ZezrP0JFe5ncEeuyRfn/1OgMbgJpmne/oFD58EmSUOlR6OnJ
XoRtt3u/nGEGGVrDA7HgH+9DGkIHQbmgR+2Ed0AyVbZ5FJNlOszt3aTf1EImtFX7
ucVdfSU5cxSbSaYBTxs3pVPVlbjxoP7al1epmykpYYCRb4xQkitiHUTXzzqUQt66
gK9SyrUOwEi9gP4gfLM0paanIy0CWkysnvJaCSa4MLWsU9Mrb9zozaYhujHI6Atc
7YrQk3EgMpf2MRWCnxQgHRg+gCeW5tBpfDw1W1SN8N00KrGzPE8sLLMhuBA4Mq8Z
h1IsIVAyzTJ5zR9916avxiad7peZ3t1+TocNamHQwh8kz8q8mf3U5uW/jR2gqHES
P2r9uqBbaO1tb9qOc4MfSxoW3I6NSbNOhiftQt2JL6ObSpU1DBlQV9r9c0szUPGg
3CXaubCi+j3bjCzLch6Sz6Cln3ZvCzAiSvcKoxQU6X5G8iNhXes1Hf2Br93M1FRs
EGu6o/Tv6PJyoVWD8kyHKWDQMg5eniYXd/NavApSizFLLBKrKOUJl/3FUD247nxu
tWP/IVjdSWdAKN+NSUEUw+fiydnZg1QJhL7rI+sgYwUqaLBPdnkvTD84gWdbSUtv
YGeYUfUMR1YJsAhLSb5AZIfoC98Sni2hMFKJWufo2GiNgjBoM1Z57Zl45fuK1KHG
tO/jiM9benPu3Mj8kQQRGpEzoszDDKws+UBAYMl52ZcFmRqEU/0OOrH76KxS7E3z
SxtABWs9kK64onhSTfjg1LSeyOxXi16vQPqAa79xOsFFvY+F0EEJ07kv9aw0rbhf
yrPVbTmep3Of2+/FAelX8d6m176Lt6v8YRKZp8+jpe1HihP3RteSmPT3EaQWK5o1
ypyLA2NG/C/wGsozSg68D/LJerUvn8+F6uuxfPaG5bxJTJ0jj1zVaHgtKkyQMcpS
zBJofFLL0BMCogAeP9woDouY8csJQl70vsU6k+cEyxNi7az6mUwbGgMcILaRRRyv
dPDMl/hyS+WuIbMufDpA/k16JOdM6Ml+Jy9XGoQ5J1jR4qUZHPtYkZ30QQ7KGf2Q
IcL8gkTIowtXuVq2arGvfdZ1Eemtfhf+sqjwEopUsABVMVVzCUMB1MZY65MFo87Z
/JEd9ObxIsvYxBFNW3hbKsakg0PmHFaTpHvPna+/+E8W7MkBj1xIsLet0b55OiYx
Jg3lOVKrrDywlbwZar06QfQO5bvYyoeOdOBMVw52D2rhOwF+LLvvHh6Jo3p2vvqk
4yPkH0d/8nkOzjdeDf6f6v41BjfIBKPfkrsgpIPjTfyVCDfUKSDV8HbKJWU3i/GE
+8w4l6oelXXUphz5YHe4gMcxkAk4Iz/wAuebD1ovIS7pmaJGs54eihs0ePWWWld3
qrljx1lv+hnb2LAqQiJHMUgS5X8u4VD6JD+jgsu9gN6yWegmRdff1gAYDVRaXvsd
iDhCX7eyFOh2eJnyrfqPhOg57kUWkWa4UefDO1+t8Br3DfcKR1AVh5wKdVZTJymR
9y+Aut7tGNc15+qE6Y9J0yua8eyhP+h5CFIxkxO8Q2G7DQn5pK8RbnnZgyNB8S3V
qvt3o604cfb60EleOPH4OpsTrVXN0bMknPM4ypeSQIeZoaNW4hThUZbme5OHoXDf
QX6MpOp0/30LlyEV2OmewtEgre7TXxM7RklqH/jFrnBrVdXnQabB6YK3+tjDyfuf
hzqh7x3ZU5hA91dgjKbpMXSFFfHLoZcV8DAuzMT2gkm6lrO87/aEVrFFc9/g1xwq
+YPSisF2tfMsPzn4+HNFszCV0r+jhnXZg3HJpI/FqvPHICq5U1dloc5/So2/zO6s
utCL/DN7oWIimiPm2yGJmQByf7FYI6Qf0DsuhAuC3PYz5fAmQ7drHHH/rsqzXs7k
IVBKXHAtbyf0HexgpJUtgOuL31YGwDnChMGTG0cm3c1O5q7WzA0m69wpzbUQ0CxH
ANO2rVvuhfMDiaYkTATVjrcOjUirWaXwGoWxli4mQFt9s7eElhXdqH8+LKANt+KF
c8n2sIqKWRgmvCFLa+uukcrpfjLoeG1mY7CUDD0VixdHDsBf4Zv9L6h5tVLrT5Un
4/4HzR92/TIfqxie0fIoMJ9zWxbRJL3Qh8fMLe6o0J9VliKO8qgBQRUaZnjoFnNt
53Nw3x5e+GmIq02bB/DiV+5fHE1JmpAliIg0mtedbH0wAE2XynxoivN0JrsWimgv
0ZNpxkgJGkALy+ah9ZLHnas+0jvcWMGJ/9/e8mVh97NPUummssTZrJjQLyQl9RtT
ecwWe56fqA4Xh18KehNHDVQ28n2mnnXL5H89OmBi7dmtHV/29SAVtfIv5qktvhwg
/hsXez6ttLtNtvovkpBZquBHdB2itXRnTCnwTETBT8duSfDR0V4r7GV7y0QguUwQ
tqOYB0BFJXodp0tioXsDXraNeTpgriOaxqonAb4P3DIKm7F9UzmUkZl0UdbHS/+9
OTNl1Ogie/ABrMu1+1vB2aona5rEorileR20Tn/JnKOzfJR6Vlx/16wGx/n+kYAA
LQk/Zmglfx9oX+rFt8siztuJpYN4caHLM2+/KlQqt5Y1uHxPP861TGSpjDjfyEqE
XUya7AAZ8u1Dp2GHITufuwY/hxyohW7UhpffozKrLtthKNDF7rBoyCd30+N1OxBz
6VOjkrouzddrfMxHa2J4L5D5tL01jv9TLo1XxHXdQ0/BNisRQIxcctjoyieLCvG9
B8XVLIQ35nI0U/QDJuloIE2bYFGZgHMRkFzveUvJh2txAp8ocnmDlSL0yFd719Kv
CCsz8hXfAIyBkh3PPwOn7J0vC7BTXP/hHLwc/kly8wEmxbX5+C/jd7e4pG5WnqWV
pZkB44lpZ5T3Dv2qgwFK2BarvJHKNez9MDVjWIl5hh0OJfTi5sh8kuuWxP48YRa2
x+PgoqGQ0UpnFmG0fapBNIJibZ/ynKWZzqSKBYFYr7M+dNRL+q3BnlMKYTK50+L9
LyWI41uOpKvpzcQo0E6Bc+B4maUgFV6Px3PHuhZdRwVqqdK1+EsLg4wm9bpO843F
DQ0mmf4+o5iM8JBqeLWaxwtnggRAJ12YEKZ/92l75yG3GIeMJcH2cmp7NVi/IuVK
u11RibBbIZSp+Ww7k1zMetkYXSlnMQ4fMgCz6poYXnJ5+DK9ZCufnTYVLnwevzHD
oVkdJNfZCiWReHNxLLWywkISiiDymOlM44TQL07mSu3LQC3zmwT9FJEMPMCzY4ZY
I9MzUd3P7y9KSf3Gm2fqzNIZ2kyuUYyXS9XAJF4UwKsRg2lURkR22Fs7Iu6LTb4y
/ka9BShddwQhVF3lPyb/X91lxDT5gFdLV5acqjralmdB/FaYV10NJRvBZfxL+zJJ
jDJZyhmUjk6UIZyQeTio1P8IOQzRehtXFQYomaCzba6cgp7qfGKWLuP6EFhO8io6
JU7IAjrlazDUKqTXbZ+NkeBJmubQtlcPC2SI3TepJxckH0SZWdZAVzvXA9B5fO/4
I1rtGYCRApB+FB1v4OdmtGkPWt7F80BsYIXlebIlj9S9Xoyv0zs9HdcAEMDfv6Kc
PEPciVhXPgSXh6Dx6iSP6pB1nWg1nBYKWBU9lOY/tlkYDjOeDLV0V0Ogsz4yiO7y
a0rroOwU6y7mADPeQ8aKBopgVE4lSCsYBEix9wcCBTOSwzrteptR1E9KLL8SpyDc
yS8kJPzfFrmnU+gAzqTuhV77fsUeIm8YBV5CbU+lkWxFMHR4vChtK4Wf5hbza6RW
IqTqcLM1ztOYfK7KWkscC9fBH+tSKQ+wNinI43fggyUHs4KZFenYskLOG4bbt12c
FWJX3UNASkpUpTgDZhCPocu9dKi1yMMYntnwhPtPyumlYYq/D4iXRH71ul4jzv2E
Qvmv0uDF49BP7i5pb9MDcAWqsdoxaAHIXBnnhK7+SwNlZcZ3COC4f3z1mwm7sg+H
z2v3lD+g5Vk764WmdyVNW/Ae9z7GZkB1wUk7speySCo57klPlmrFhmlamqFn2NHA
SNDhJqgz2hn+qplV4iBzaH6Cy+fmeWgKx1dfZ87f7oAq6P4E6YVDoMuoZ6dR0P71
0j+PQr37yv+lamDid+1yj1YnrfzAAwVBKhmJs5NFLyJKrTOiLUgCes6ydT/KOfG6
mdw10+eyWAItmNFivw2xCesD7bTRixMay13QDJeJZHi0wkvJljS8FI4gZTFNV+6g
u+yFrEAL4ESJAoBv8FLTT0otx0YDdthbWiCaOyf0KytaVkdDOxc5UBN5ncsc9JwJ
JeBW7BEjtNbUzZb8BgBw3GOAHqbVDeWqd0jKEMlVUuLuRxfzmyJAYTT0T1ahozrL
ttZCRdNgCCJhrJNlGsQGCDYYDTgCQzalVCwbzwuCASWDmzTWqZZp4j5alURHYalH
xRP2L605i9D+mhTOXMmV/p0+TrjApgonvaZ9w12h3deLu7OgGC3bm+llFLCW2gcX
DyEacTgl6msiH7OFRTFfZ9Dxcas01hdDx0xqAWBsKEol0+g93qIzL9T4BOAvaxEw
TzlJ3QdUSTSbdqgAQeO4bGabbLIi+NfndiP5ar2tNR30vTlVW4wIbP/avmyTIBKc
942blSWmX26rY4H/8TK4dcJ2/gkb/iOJY1GrK8KC+Ax0mEVvss621x9iDNJ5qlMK
OKPxeUdaJuUFEukaMEUKC2LhwiCALh1ySP5HMdw3gijZyJ0wfMh3JDPWMZpfL95D
IDCgauf1yo2zcfA8msm9wcuKvgIr9u0slmlGc3Nl3Jx1vztSPT4/v2zrBKJe15wG
3ObKffFQKGn4fW24QZbH+LgBORKUzM8Q8i+tlOSYUzfcUodV7UWr1OoaOLlek7x8
VRZ62mJiqL4kxkZkCGXaIJh18rziHlNYJ4WjN/IK6xuqoZm0300quTVuJMxSEJJZ
Po9kMLCBOMYMwvIbxfkREWnGWI5/9zyOJkSfoa9jEExAGBBjx4V9ypma+7YlpIuU
Z/nKNZsYXcwJsKGddUM2BjDqdQKzpOW6wRaqmlwXjoU1f6txHjFr/fvQq7M1f2eK
/HUMHiby9wIs3wZnJE+x284bX5vbMPcdFepMTHOV3MHhxcGFJ9cTeNAOhmoJ1ic0
1FnXN8iFRVvqL6zoKPYAGfgsAyci0o7/sWejDBe7AJta/B05eLzpQhG0Xme8KWsS
B8Boipkm7Y2dQEKebXhd/Yj+A9c0uklKRaW46aj40augnIKLpJkvLQNvADWTCtaI
6F5u/3Lp8D4cfsarvni+kGfUILDYnJNM99kxtrEbINJNALaEJCXzEKGAFvKfncz8
YQI2E03FkGVl1MUesmXHY+VVHrlyHmUzuURVsoJ5EkMjYSSCYtFMbcgMPFE4grOu
QBFX+GWyq4Icd7OjGb5jrH+aAMZ8JXBAmxJCBNeBEXJkDpAnONHm2r5Ds+GV0Y/8
Mq664fucI4VMjRlkddFGI0BtVsXBoYOcVMSmwb2mGswylnrOkG19JVrVnm1PSfZu
r+J/Jti0MnhHPezFJOmc7ad5NtIv9O0KrE2lOYNPedHM4m2TlPdpCroLf2hSlaw2
4jCol7HFbToDAz+5i1ITbqCZyBmcZhd9HMlL2B3NWsngJdlMnNOtaUWhsZ/gEv17
2+b5psuHAjxPabkKbx1lXJc0W+61yuyb0dw21o1Epy3ydHVsuQ/2WI1nNPdztXIg
1hz9RXlEX2HSHTAotLr1BJvg/UnuCHvsfWHz0rxarTq5oiQGqc94vVYjvSyj8H4Y
BDPtvNubTOeHfjzncqHv2irEUkbXMaq/yUL2cVtraf8bd80N2eBecGwaM0RzEtKa
MKImYihR10eWpZ1otoe4DURXzIKaJyBnipQpT1IjXFOtA1aKSm/RMqDL0nh8gikP
iShpwm4T+LjPwtDhmP6or3eYaRCXzLsGsdar/9gaJ87wXXvI8Xm8QzSI2MLJ68yt
DNBD0Q9T31gPAgCDuBcgX3hme1Hce/ar+189lUjIP2aXJaelxA5MF7+Jcs6STM7a
iMAnaA17oRI8ClmjtHp4QzieQ8uTzinkRITaAQ30jao49MHbx2HjUAhgebnVex5J
OLUNCf9KFuM7AOzR+H640vQ1lphXHVgnAMchqxZAImjA+SUvrYXGUMuUnrkHO27g
HFhFNmM6nV2RBgW8rvgQPVA3SkZP6136EmCv7h5QhvnjS0/9BymGhCG/ht/6wFrY
NQX/rUtgIVdAu+vIM/LdkBIyL6iQsqAhbca9mBziaNmyzwk5nWttM6wbEL4kyfdd
yQ2W/KQHTmdmua4QW/g59F/61A+9ohw558LNkfhjgX0dbXGgLNhgOcPiw1/BEkQj
j+sYHGv+2KIXZR44ccuqT6qvdz5X5kXB+TlqvBHdmM+R2fR+M0/Xs7i++qPt47OQ
IQ8R+1oU4zAlibicIXLtAzbQ9digkAT3kkOBJaLlPtlhxCtkCLIgiJtV0cgNx5Ny
kRjA4ftunKp8Twv6+LJis3wT7mPJYGUpheIrf/sYD5VMVx5Nvmk+yxqdEiQJdwq5
nQ/nsPqP6hBj7bw5Kqd7Xl2cpNAK1iQ4IgZ3UqQm3WJdkvGMH3NjiinMw5e2CIi/
j6WJ5t5JCBq1LzITUHeF3YMrVCO55CyxjVYqplHw57G9JdK9DuI7s1Mm1zn6gCsW
KJ7SG6s4KgPGfIEp0l6efaVXxMsqJaaa1D4PDQN9ljEm6hGP2ejFuWrm1f0fP0mP
tyFqHj//d1F2+kEZaQjbaYHNcDKTmD1h02mK6jclCG1S53+FvT1WVbbSvgdDbysn
Q8pu9JiIDU8OXGZkZp8qCZLb9Mbu+rCmAT2u/81JpRt5xnSgP0LHEJjOqWTXmiXP
FsN6Vb038Z/VOfI7h9rSCZmFZYxsXk/7Bwey3YZfY0m79cNtCyRcEn0i79GXCCDK
mEUUbPcQIIpqchXUwS+nh1YWEo2fp2Qx8vBFSeaEkAO1P4HsziYfK0CFq+OXdfpf
1HiTj91govK+6OqAXG213ulDZT+7pkqN60dQTrL09NyQfN170+lBoy8WbG5CLfve
V9/uOeJepJ/oyAot1SKckWsbKp+jzUhtGOIfa55fG5Ov/AQVmc9+i18PA260DtBt
GUGjaTbjTWrU6575+XV4VF6ey+PCjMMUK+0tEQj/8Ixa8w2RpmBSyjDXBqScKOuR
OSeCFF03L0/fxHIvSte4So0CNGYyqJEORjCLtY/zgk1hhAzs7QlMhttcsmc74bHL
klYbrstuhPuGtUrd5xWkbtsHHSDvIyBa9EAqf/9qCtucdboo2hR034YhaCyf9Qb2
T2ZwJcMRJTaATkSoKjS6MwrnNXqY0EZphR5Zw+2V0WBPQzCpFFS4J6VvuYLcn0qm
1x3/EDdBvJBf+YzjNnbOjRb0SJoamcoxhQC2QpGCQyX9hw6bDlmMq1fK8ucpKtXx
Cl576jLJs4NGxm8AK7b0eE/NyMdBDrKJliZZ3IgT992NJkObCOK6HdnZlVPIFLro
relZJqOx3jnWjzauh1ve8bAwyZH/a6V58Tm2AqSmp6rhTINSHAh3tBYOVrszciWg
hirsWHiaDOJeFsdcjXCvMGEXdWu6nwn8N1WtDKgcZ3jHrjetw5fWxyIxgZ9gSt6C
s2HOcrzRkkKMZci3vk84G0RU7w7S2mDnzAISbBIIYTTTm4hXN9WwS7Rs+trwoB7F
bPhQBxceKm+u2NGiIlmBOP6jwK+cQ5n9QhsqWJ6l69GqAMFgNv9UrMC6/Ip27fCl
/GqoiX4nuTbXh3oxwz8he/JlPaBNS8kZhjQu35ojtNG5mytxhXpMKZl2pa1+16T2
nLJ9i7iXnHKZEWrVEXWfCBKnP0MjtEWvs+bTFeBEcCxr3RdPYRcZDSAMuZfM73hC
wpPvTvJTIgYVZmA5Uhon2eI1G14c44ChGZQlbZmVU1c2iw1hkuuBTWelfcQmslxa
PXegvkpeNCmsHmyRo8tGzlHzhM/bVUJEX/5rNQcB4wRCIX0AUOFeT7XNTl2jqiSt
yPDz3Q4eaCIdllBYB/b7RYv2xEji2Phk9yifAz/SBQ2AOZ92ukNimPhTWJ5ogxWJ
9tdrh8t1871joh5QT4x7oCz6SIUxSMV+8Kjt3tz6R28VEMB0aDQaUYlF0Wjo+SLV
hdR81X1U/Ul4C+yZUWTYwFdjnysAyubVhtLwFTo61OTc8ZSxMToAh/sYipayZfLD
NcB7t0HDooAnPNqsios+RUACwlyJqHDOWafICIjoYZBDuKhCLADICxAT5O9C0I/0
WNqXSrrbvKgusi39IBtUDGvP1WdWJmXIzLRYM70feJ1mgMEnQbqhQo2YdktBitRR
1ldLo6h652wtTsyUVyARKP9+CJ+ZgrBhVL2CMipva4RCDn3ax8NDfoGflbK5k3QH
I9lhwtITzYZWHXv18lRGnyC/tkGNr3UDhaQq52rKJAwU3uk0S03It1OpWIAchKga
87jzkXZheUrS77fOfYPXpPsDcDG/tXxMi3B97DKSZwhzyV6oKhJcV+4sbKllZmbv
j7FIhvweRS9cK/hskszHQ8d5HlyVFmQQHA7JVGpt90qc08z5ObYSZygkdFbKizEg
YbQtn6i2gFj+86P+3pBzBDEOR8yWpVnGuuGIpf5k5CPH2UiCysXF5U1K75Si3BKN
Yj9oheAX1wKO6lqvyQfqYh32IhLIRNBKRGGsyRJ3u5FHvxfVdCIIQnmKi2Qs7cNR
5WBJhiJskS6/PWs0Id3wSxP/bGIgmevIKGjkeJqpEn1B7ZZrXS3JTsg2eSBeXx9/
VMKQdBO8fe7bT4J+78K7wKkl9UeoeKdCSXHc7PZYHlflxrV692UjfoKk80MdVHzG
fHsVLlR0NCQOj1f1a6T1xgTXzC/Ci3dPaBVzC6fCyZ1/W/DAB2vvk6xTblKa8RoL
/vOnvVO0/YQva7bk1wVfHeLV5kD2DBWNYYp7TCEtgdJhBQAEj1/6PuF919P9O9vc
RZdpv531RW+yKyYHBBF31H37h2n0ONx/2qRvQSE2XyQLy9w+gQL3i/hFS/KydQpg
51nvOAV6eDksKg9GB6rNWeY+wm4+1Tq84ZG+I3ImYSC/xAjq3Q+Nf+Xo/NViM+kj
4G0KjzlWBJ5GloTQQW6MIIg8Dt6KghHLvqnh9PKXPcKTNFmWgFU0BywFXQT8PAop
Yliz05SLjUK/WzPA0+QsMWHqxRZGMKYWbMO5r+jknWafnHSekf1pbYoT1uoOMu99
G6P/e62lIcIfTwvnyZrxbOwVCUGQWNcEq4vv4bysn182Cu5O8VvanqU8fdm0O5up
0MqyQ54acryGYEImTKdw6yU/lwhc9Ls2FzzRs9yVYdaef1h2wW74oQS7GWIlAUdM
rpQRvlaZedDMlezp4pEtUqeftKByejXM70TAOFPHNsYYRGXrsNj2KXEQjzLHvQ25
8tWo66q6s+fxg+LTKuwcXqiqT4KlhKhkk71acwn9gZrJsIis3m5jcIbPA+ikZaN9
etaLADVgO0VnWgiXWkX62OGEiAVb0kwoP1WZLxQHkJHsSw7oRC1yQUyK+7+kh1JT
miB1zglH2rJ/2q4b5vSRgNKJpc/mixY2QL2rCF/QIejImwa/DtfPrpiH1SIMI3u+
4utJfN7Fgr1eD1/xTUChHESZsE5aDTLwcscVgkO1XCpq+Xjv92y5LOgpD0ZnJbpi
NpfMkiw9zCLTUr7psKKxSVu79hjvpt/pZeuX7lLW5VsMUaOPqh1IgYCKE01vYN/y
mEVEf51A/hJmsMGnjOgyPbTmZB+Gg++wDpgewdWgbkn9xG89CN1pk/Yhf19C4OGQ
vVsOsls5ObbCuB1sh1IucgNpd2fsGACBNOnUEldK2XfLNK+dn7M2Nzsc2cYVk5iZ
RDec301YRZ9iplude5wkdTiYiECa82sOZAjoPD/sEzgVlAcijJmcqJNfB8FvS1cG
nl044WeWQYS4N2sXtNvZZOUSIHNldxhW6gz6oTGCJieMzOGlpQhW+8bFev3Ue8WC
7gFvVdGorkSzINbuXPkIpoa5Ntbm2h8FgTZvLpTXcqsEbm9WLU7bWxdWf901ZMli
aSDX0dREoPiTSSKi3QA+otTq1kZ2fJXpEgsn/2I1jU62hXPwwgIlO68/TURSrYvU
SMtmVKXZ0dNJF4++6dXpVi0OBtFfw5RpnL48LVaoq5CpHmykyPGGwlukrk8MRo8x
D3brKqgDCXbe/ji/pv/arVq70XdAm/WJLfWvxuRLq3eglApBGRpirblvEycCJEs2
moFyuFQnF3j3y3NnuzRvyRwGaQjpb0nqdTRzEnRcR77ggwe7UcwE1hvJteDbKpQE
21Exrw5u02W3IN5+MFbYHqcUJK9yIlLLi2mwL/iZilVVBx1LFF/gDWrO+jVlUca1
IDP9aE1Ea6cGQS/vxtNBv7tN9Pn/VG3I9Abi32pBIizrwZiTvo8/DEFwSJgyJ2HA
f8KNztXbRsWDhsogI4hfmk/YQ0aJ/v1AihxAH8sfwK5u/MGPQE/idD60kWQ3tmux
97FU5bAPkfTkyDYQUJ7LlAIfnWBPZp7Bzwb8lnW+v3m03EolQcqxv7B341rf+27K
3LG9V/73Pf7SEOOkKOCD3aklno+/OjmsNDcYf9/j8ec9pSC4ov2nIhSHW10IMGst
ejKZ9Js/k3RFHtAKRryaQYl9hPD2+oW4J3ssHzLzrb+RjSYSbgNdHSzb+TfejKrd
thm9AnpEMYWmMl9XyyflwPE5dR7Vccb49yU/SUBKxXlqwzZuOvEV7A2TxqFRBAhn
JvpLczZqnXKbQHw/52A8bxqREFUKcae6thdp8hNxs2rDM7xJu1D1TSQAiu47U0Z7
p3GmujcNIufDTzGVOez/WQqZwgBBP6K2XLuGI5/8ckdimS6/zeYkXRTDrBOdA0SS
jlVwGIrbT08L5bgMwOPWTIZuZSixJ2KAfFybXK4T68HSRwrrg4aYhuL2WBXpDEg1
so18kKiUGakETa0IFlSPzqUASCna6LOQCMCHI3ltH/+hVQmA4aczceA+Gmcc+Dom
dOi66FAmLsrxRa/FlaJcttQZXFFLMRnZt350BumPwD4J2DCm8hZhYnedBPTG22R+
zuVQRfGfnk1YNbss/XRFGkL9y/PsddgolJ/6W8qrkr1tov3M1owNHQinBZZatFCs
Idi84N3K9clcw2OQI41pfLgjrEko36ibth6r/Sz7q5u7XC5Yycah1K8Q/ISXulaF
NaCNs6lKdp7vdsGTOr1ZBYwDceE84TvA51G6iD8gD7yxC/ZZ3/l47HWnyeiiADS7
pSEz/H94zDVmh36e3pDioWY2u6jfTOAtD2DHgVqRxCrQgMoKpSTNdOOLbK3uzkc7
UxsRl/0xNwE/O3But/s0VuYRNPKClr59t4yS4sllZ0nqV9pBqv9r/FD2rhI1du8s
Idqj5Db29LZIGM2M+7UPKuBA59aRLwlAisoZ1C3E2/0EjxnGsUAPPjgcNoMSpahQ
Ez23mYRUkXz8xfvlNkXGlVOwatoFgViFgZUSySFI+i+/20EMlXf/OSE2JcTI8YJ5
Ht1isqpiW5Y+nv4eBJYWXtgRyFK4tsFgW/qpoYnFvNn0A58DvG39VoNpbCrcJ2T8
/S0zXI+K8hzimm9ARFvM7cUvVSmWmHUZpVdCVDcSDP3bePYmsX6PiWT82GTDsLks
DHdk8rl1ayb+lFloz+vrV4BGNxw5m3DhVOVQ4ZL+fZFOE59GDvuVygHCG1DRw1Fq
O8OeBJxToYTIVQ3HMLETzvE0Kdd2TmYHlr2w/DlBQaVNOUQnJFyQnC1X7G6PcVW9
sfam8uaa/AbEwmVsGXDd1X+/B4aENoJv0OuG1BLXQ7I3X1b2nAzHHxBDeywK6dbZ
nHZ1NvlyOrnBh+wkPUTQv3ElALfUmeBxwfTsoZO+G/ZEUPxX7Wp5Ueev+yXup1vo
wzG3xyqrNuTSkueSvpMprzK4hwHqdkJK1LZ2C9mOYxy8ubGrKZV1S88uUGYrH2EZ
a+XNxNnDfubuq92yDYXIEJZims4pDIG++54FkN+D9Z9rg/PFVU79snrxOPL9AAXc
iOhX+M2vhIjK+CKbHM4M5ED7P60A6n4IROce3QvGrouecjNjbJ1taGtRkCFS/Hvh
qv5a3ynPK/blJT92QwOa0HY/122M1ALgcSzf1CWe54fjy99guFh0juc0LzNC8iBJ
k++QZB7ImeEBvrmI7vBtcSA6ubZH6H84ycVzwS316U4pfMjdJ8XuJTc3DvmJqlVL
S/2uaDMf6GHfyRtPiNEF3EYCTBUpOD5CN2nQin6ntvVE5UtPhykpLUf+d7JFc7Hi
Yk9VVFyGgsLJeDIyqBCfJPz+/bo/9wVKWTg+CJiyNNBSikl8XKWu0xljx1TGKHm1
fdpyngO+fd0w6jf+FtfA4Y9EPPSylYbdJ4TkrCiR2ld8HAGlPntFrK+8gbAjk5YY
COKPeSsasad8KqztfhrIwly/DIjyGaKTW9LHZtxtgAWkj7VZt56iF5+vsG4dDVHa
xY1RFEo5b7OcG8Vcgu3VupcCbLNVbrjF/HEPxIWOOnmj0oR3jqWxYa3z68jKZNLv
5oc5BTAMXzjjtPsJ0PP4YdTtVNtIVpRRQupSckYqvfRBZ8bDkVnEqQyVJ3q6U5fK
zMM700RIpR0lnNNQfh6IsqQVLCo+w2mlSXvPeA2ZcCH6uaBCh3eOx0aKwXU2DsOY
wZ/nEOHuJRX84M5c3+behI8INi/YcnklY/ZYGZA2ZHTo4che6ICSbptGsJIMnbE3
eFmk2C46gmje689T/XQ4hyGb/Rp3cPlossCw85N5yyujFRiHXzn+UYf/24IrzHUu
bUBqk22heIDWDRcUMQdQG4zNhC0SyFbeWBSG7Kuk1vyNvZOuwK9smckGaEGe2QYx
4df1pdEsQjzLAxrEdcJDHTaTW+Hoz8lB6ah+JNkLRCLp7rUfufwErglGg4Nd1cpm
ndqBxFJjt+7JSY0xPYPAs3QKni8w11FMPJTw/EmrFxcxOqoaqfaPmfrk0fKfHrsF
b4SlhY+Ds0JDZyEFIKijunFjUUcv5vfEQYJU0FNB/J4C+HpcwybYpk2hVYrkpLIX
GU06Wc5mQah//8UGNUryF6QoES4VYTumpefmfjNaaCyrXHZ4eQNJJGqIVdHJ9jb+
qHEsfrBcuTjTgCu6p8NkSvee65r5phLGEovn2C9hnMO2KShnFaPL3LxCITu+XicJ
KM184d2UpU838X5yd8euOe/jxrHGH865Yvg63A+5SEWqTrpvrRMJo+QiirRbr9V+
eAK8/lxcsMhUBEgoHoZAqA73TcWu76fQ0kdcuR/Q9Py4yNwjeRAcdoKkbGTMxY3f
r0jGi3FT7ZuBdgnvvcy0oKBq7Khiah9kqj22Du0wE0o62KYt/skTRLJMGhYTjCkc
eNLa+5eBol3KmrG3lgnnYoU/MleTGyv7AiwEBqu+ZwYxQsmhT4efoN7s7GrDkFvq
0qw6yGa4XOEB1g6cMkoYSKdVnQKQziSL2JUbe+Ekn/+eT9260HMyVB/cH+YF/n1M
Xo8EGVo0L1BmrQBZpKlgXf+cAP+FwZAIj4e69Gk6fD5vM53I5fhTlZ/N4Wyf0kNE
mfzOpgY95gtEWGWF5CtgRIdE6DiIahaGquuUecPlq9TLlUKsFmvKaDIeoc3oWa3z
Vu9MI6VwsFz0SStgzNr0+mGDA0qGLCllfGlYOapiZEkOQLkPhNJabOUr9KNMpvia
Mvs+/ISJAAWw+yztmt385ldePkxlRTn1iUkz1MK2nUUeBwyrs6gbSwdvjGNK0L3a
KsB87E4bmIYShI+gXQ6qMMjYH+E0iRfy0LWj4N7s+O6mO8qiKY2VoLfaq92cDNF9
DcTCr30Zo+Wh7LJTevhpUdUYgwDXbmuttZdRKXPudjg/WE/PTL9yB1FQG+jtRSoH
c3AEBJaSG9kjvJfJxlnes8/SQAywlFR/kNmXwqwCLX4gX24M/pvSI05+klE8puP2
21NcWHk3rj14QLQFVQ+fbsNwbxvinPiz+AIQg4bjSvt6DM9YsHHwK1mhIpR0obTU
sST403K3XbQ7s5K+cnxvDKR8lPN+9IunuYCu8amcl5q3tVKua4AopQTpHU4l9VT5
wGx+YDp3vQxW30N93Y+B4lNYqD3vDRlJ1xSEQW/tEnL7ySz8mfsclOMeqdi4Xkdb
5vgQvfCrev5u8w+whSV0lQ/Pc9eal+Dqfca8/F8TfIqQSxY/1sE6dCkwnnKtEU8Y
Ait2dkiunISXYnHv5E4ooEu0RP33zO/R45j7gaatOEEqb+/jh5nZ634/w5BAfay4
XJI375QGD4cgz94Yaz+q3GTeqfij81MDvlN0OC7mbcS7SVhYscSLuxvWgi0OfUAm
//6o4YwwOma2oihJTSYTHsB6RezYMWBRM3e/X2C2JH++CqCKijYBHzAp2X9OepDC
eRDYowfBgio/0um+0ykrBxU1VUPGKgp3I4ebhIT9NOMe6MxKVhzvwtCx+oWr21+y
cq5gZI2dJJDVWJWeKBIXqtUsdBwAzcY+vJpE+hKwvfXxbbPSvGDnSAX73aUxQkzT
Haz1RRt1ML8B/jTGYU/AjgEKJPixPffeKlOh+QRB4xUwgyKH/80pwgst+s+CTu6m
8EufFY1K5drJsuuOVSMFyRK65gXFsMaO5CmsGAxM4lAJS4Zfu3/NeZTx8+cQ0jx6
ddTFn3/bPg+CpF3e+uf2W079KJrQ6BuxoIrw5n95O39Ye0caqVGvgMtJcVBCVOh5
dU3ShvsxsgqL7zEsSVIvmEI58Y71jyoMTJKV39AAeNsAVW6AoFFoW1HV6d2Ptzqm
Wtb9mAOIAT/RXGsVyTxP3+ACRX7HRJlU/1OfxGfKfpf4TBeWbd7PFWLNROaKdPKw
emD+x3obFrtE9Iw5ytarrHEAU3NCk17TASp3dBPZTt6Xp+hFoyvUxPZRuiPiFCZx
w6+dcWbPV1rxXfXjwle2ZuYN7TPlgSIdQCLgiJkq0o6ucqrELTOTkL9LIW9J31Ln
13egFOQLSmlpUFQguemLuwRW10ipSwpFPpNTUXipBNfL77hfUt2crddldoJHwOrA
EzBY3f3epaihnDr3JDpOGTa+qNDyxXecS213ZPdk7nJmfQL/x4Dacnj7jmI0RMQF
roc98k/KKRSr6TqnyJYHjtP54mZsS43lW9953oU8GsxXee7H+jJSaF0thNZGKD56
Fhai4DBLnBvAkWGupZl16qooYr8rn+vfu5AbPlbmQGj/qqfmQ1X/nIlY3ucq4KRb
9ni03NkVx8hSTdDrCn4IUwuBe4sEl+ZcZghqbxSSh44ci8phyUBHUj3tLazFYVo/
eRbWXzMFnSDSixdP/mho+whOCUwj8dNoGPFxzlGDbIlLmRy2o9nhQBc56UKGxTmN
+Yb/7X4DwLbUU+ZXFoKaXFtp+XZdylYXHcxl5Lurr1du9udODrD7IcOgehmWKzyx
QQsgQL61TWXNtOFm22r/JxLut+8xOXLjIjvlIHPOVYuw70UGTKxkULt7P2K8qHnv
4PBnFWwIWqC8fsRfNMLAlpiobRo82j8gFFIlpcJNLUJOfn/uM6V2pj3TuqJYHR1o
cWznlXLWoYkggzn1D+nJ3tMM6758r3WZ6Hez6VQRR248cmGk10/oRYNGPpMm+wc7
QlaL/om26F0zv0mlQjZQfVTpsI04A1DqT5zUv/MHj9Z5EC2jCFHR4WytGAkdo+dq
2lsmjvG3+NFlb/WsKolZZJYrzo1mLpOOHW1vl9ayWYm8Dp4pvt//vhb9TDx/oS3J
egtNMB/I1rBAiHsYLu8wGshkWD9FahpUwJglUIr6UqXCJnjgE38de/7iLRdQ63IH
JF7hgcX6ZUL1wLd1Cb4AiHV1wC7R/JJZEH2ljjJDujZpIQwuwBTM5KpYDbgMg5/W
tGMNI8CSFciyawWjNpHSJCbboSiF9DNgnD0AFp0B4VJC+XXjlMGQKc/Kov7woGbH
bZBs9GY+HgchqVg/FCqIBWxMIiEEk1tCVjWcFfzDM8GcBqpIwQcyQWm/8DvSkDD6
yD8J0dryu3eh1uJTafffGEHxdDS8K3aOhwQ8gEFdiMcl4FM3ESdOghTsXjCrOuif
Z74Qi5hPGr3Br2qXPbWCoh/lCH0g3kyT39mlSwBrHilgOWm6JtU36UsH9QUCvMnl
vj5fU7rG8WGE5Ju2Rjl7OCfh5qq32gR8LOLz9CgVqF7y3shhZmgttUfYkCtwjcva
IE78wp2XdX8S6isVal8RVekKVw+b7DzRbO+022Zqe4O6VDK9WZ1KKVa4TSZSv+3z
2y1d1+r43W8Rs4IJ+hSJVOH2N46B831yLV05YaX9rwAYc4/UFGJZbJuvb0tfhtq0
VPZ9VC198U0hXtZZV2BS1p7Ujs4QTt6Ne/AD6FBm1D21RWMv5gGQcYuHk2NRKzrT
dS0M4dk8LglVahth5Ih5zNna+yaIxTyNOUzsZcXukTNFBj7kKA1vQ6/GJPTc+ahB
OVjd7TPCDrAQeSBgp6B8rp7oLbynVY7Gs6UG6EbxSEy36zL64VgLdwzlPSfnLeFs
i/hppUDYa0W0jTUU49e0cpyA3IKpJr1aeQAbcLU7ZZH19Dw3KH6MHx7wIkMw6HHD
qzbf4GA2oJrHJm5diyqA3sqAMSr0smR1Yr/FAbYtTOTgk9TDwuD+NO/Zw3OAIIcW
MoJgvAa+at2Sm+Ocmxb1rhJoTPkJOGoY2nm6lYfdvHGhAou8pYsxwyfbULi8insO
HrdeeMYlVWQO0aWFHqq0SWlQEQysvN5isl0mT39ex6k7RuQbKcwH43oLty1oPDIa
aYL5FvxP6tHMhIFuj+wRXdhk0T1bB0xDz7keYV4BNUWneBAnBmoMCQNpqjfr/l8Z
J/oSmJe54DmZJM55m6fu0Urxq57eVISRnkvyjjGDntDLx61wfAILbmEslQ4YooCI
lNl5l19GsrnfizokxrsN0gXo5RqAWRoF8z/xmy5fEiGoFZHibuCP/20N6rjTwJaM
L9N5oacI+4azPhbSdpTD6PWoeL64aG2xXWl0lXvCBZ760fHImZFoM2gP173BWT9N
8cLM6YxByrmfQPRUyZkwFvVf5buIXyGgeqFFmwVG6rsmu/PyR55NSrhF/eCv6XQq
gtD9B6G2cLN/uDU8l/41jasUvunUWQZRb4oOyaMiUJKKQ5fAtqmzH5XFWs6jvykw
K8RU5s2435YbCYNtmgxhFFU5umL0dhRXeDr3JRUmAj1NksfRadj48imWmwbSitul
O8gMotmQT9QgsN3RYNEjQp/qEpiSxzEBMzAqjacSsi48n8C44ix4tjrVufu0bFGs
nymLT24sqeohKpLGUle3GBwEPZMv4wiykzFa2D1R1yhxDOxDU6ccMvbaQX7bQ2m4
xLT34RxX8Ccjq2+zWG3++VeEiUpdg/5Fgzaalg4jyaJojixMn54cEN9GTlxM8zMM
YpVD5tQ8u3rww0mg1W4Zgz64iBLhmmqZ4gsS2pyeXjB4JMluYoWkAssH5qbTQ/bE
/8bcV/U495J4ZlsYJeY11yNKi4XN3p9XP4dPVyNJAyQu0TNdlpkv2Dhm9Q2AWXx4
le+ZFwkWRg1WN0P4agPx4MDuFX86LAIqjpUwpRzSBb01G4jV6DQGkCr9gSTwU+V2
RnQjWV/qv/ctJaLKjYx0jdz7wrpKc0epDi5vmAPKAogMYk93iMq++v6mng7Z00fB
dnyNgW4CspQF1vZ1ltEytukMslTJmbe3oOArFht8kiCgbCelDTPxWyb/x+xWiPhQ
Gew53XCj4fGTPDCUag9ezOeFL1PDR5yeXwgn0HvtYwAq9uBQF61iF4px74SQKaAs
WSiTpXgr5Eq/RuaRIMgwIg6TV0x+dThTUWbqU/cTr/CaAZB7x1E3QGpBZm2K8iWt
yJeI8gcrhBTcPELNB62VFz+ccVDecsVOYVwXVYR1lVKJAQuVBGJCsOZvZ61I9/uU
UtrwX/avPdqJwLXL9nThxgtN229X1nfcVBhXh0cm7SO0r8HXrQ4SbMTaFw4VtoVm
/mpedip/hSSeb2BdTH61wv53D8yd2tgtSJzf75yyaJbdKQMA8uK4T2oE5nlp/8YH
SJJ68TmEYK+HSIPXNgt8mo44GvaBQhBitVw04aDoahBDAftbXpG9Qhg4gxJj5ipp
Vh2hdAP3mQYIMD/EDRi2i2eP3UPzfvNFYis0wELlWVtPJ3EHdpRU4K+AoWDDjb8/
6t1mfNNYxSg7PgLRA9Beiz4R7XCD6/qIwQxhrdnDyUX9c8crLM42hANJ29jDjjAn
vi3as/pQ0+F8jmCYLaWyxnJhAyzf9jPSX2UMVChTlW7y3dUTB/TdOyx/Z8cYohdy
g795qsPOUtrbvvdQLM1qpz9ML9fjvThm5w4clSXSRzpGTrHMiUl5UXKf0QxVu8yu
1lLfmJwPkLOZgOPSWJp1NYZ7sHaT2AQedeh2Vb0oi4hAR5y01U53wH57aELu5I3q
/xQNiUUum8qCeHcamAtZBGpyt6MN100oJzFu/HJJds7Xir/nscc8zCNpoZ8HsCU7
FMRuvej9PAXVEthq/EJXHBZmEphWwQRxt/RRLX+bxh8/LHEAmxNiIx02Zmn8XM0S
TQNlmdaGawoqAY0GdMnSjdtlJ41V5PGZlbCknbQ2Qfr+ioudgxLgDebe1yF0FLTX
VM6Pq1BMklAE17r9zixK474bVWUnbYbM+L3YYhU3EJhvv0duVkoz2y/KLNTRZpul
H9NA/QPc1166ze7FndQ//luUQs9pBNtJWXfJXWymcJbifjeMB6O2haqN+wKybIP4
vSFfZ7EbGZY9iu4vKzwak+TdlVPgO1Hk7fixtrwNp4H2Xqy/kM8TSKgUrRBbSo7C
4egl7Uycr7NuDC/jXIn6HeKJ18mJuOAs0Mk1HBnbh0A8QYqghZYBCtrGzfgU9SFl
xyWOVlMFnB+ulSWKjFmqcsDZoKQu6KFJfYlIkL9BDeIEMw+b6uPyU0dYi14KE6HH
GcdNeZ+8v86YqFv+opFVElBMeM465ddKgCGUDSeyRPRJ6xTHcMYwkDn34bZ5irzd
1fSMlED8v2mFxuRsaHtJH7V2PqGqX27RFVTMdOq4JS8yaP2KZfit3KgQTxkA064H
BKw0qEmj8cqhHhba88DTqZpJxcxjby6c1mj7/nE4NgjY/aAL9lp4KyBMlPlTCU4J
iBK8yuw/VYe2BHeVI0To7OzaetHkRL4ptxkAmQc2Bt38A57frrxtqHkq04C7/8o1
5k91GaW3dx49FD8fjfMy4m/CxZhW6GS2YdMjEaQdXF3U8TcdcH0piAd5IK9GcnDx
mJq8ZUFkfBLuUd19B6vDNp3mNa8TIlfYH7+ozeWWk0/YXg64HkH6gP6feoXencII
q7jaLwYH+mpJGuTxQmC8xw0ZjWekzHpXXFEinSy1C0OH9mKygQ5HcAhf8Hp9nRvw
dWNljFMf1ex0B/kc1uPiskvZvySN0umbhf8K5cB6yvv0pCw7SReY3SO0eaWulCsO
6D9Qtur4ooC744YhZXkq+Dtt33VoSlFTffwHpuNDVCA/dcWZUp145d8Qel4tXutg
3tUwvE6dGHorbIQ36crmO2NwcNQwTMFnJIeulCOx9txo21U3q+IwMlClmYmQId4f
P5ggwmGVukEf53FxpD5n4v0n+xm2Ki0L3EGb9tHtAf8lKoSzSTkhjglAWrTcUvzj
quHi5fyFGT4iMt7uHB7cokEmDAkp4xDqTbsHBNU3KemaGwrf4v/HaxIq4O+w0uKA
I8H4iTSnisoo1QXV7h8pkObrs4glJGc0x0jFCQ2eGIUXZlIlLelEcZhOK7enToAy
W3B1U0V5Vhu1Il/bMf8mxWt/EjWMKATyEwo+1vLvl7nbMTilNojvdG7qNvIeBEo0
ktDP0pMn0p/SzN/JHuiJujZXE9MGuiVu43q8U85/BKLDwj3VhcoQxZs1Ba9HDJ2Y
noiaueld1QANXYMyCecDqK+jpK2qFiqofs9EWo1BsxzG/JHSGdGbPU8Z6xpFigLi
XAYFWLyNhlGkKyFRkZ0/Rb9iM2WPM6TuApdP7hdAxm+W8wsxDCYBsHHUMOJbH+tp
ADYYTBqqgRMx3Cb08q819waRv4TrYMpBbNOd2Vgs2gQgdZt1zrUEC47/rNO5og4/
OawhPjBGZ6BowISRFuM/c6VJM01rzKmr0BSSAolACmC9sENbLvnK8dTqKqvWk8U2
DKQi0VbNWMGy3pXUEPCedS/6ydQ3UjeLlrqUhwryv+RzglWmrC3hNhwuEnXr9mzN
gntHTvs/AQEzMT4vZZ7FYs13RM9axFy772eJT1x7qPOUIxYq+QoNpSm9woiSqaql
ubB2CVKpgFEkKu2L1oTW8eYZglgyqiuVBrpZonjEc7e6IkYXCViIXSje858tsjhh
bu3kD6M/W2PIPC60L5NRSNFn7mWY77cRfol5NRceXWEis8ro9M0ggckiOYhBPUsi
mGhULmOpVNLngyK4nPjpgMWDoMAfCg+LuBOm0WAERmHl4SITVyovtMx40RfgVF9D
YhzZZAWgARJfwHgvLVxS0NDs2w42CnC8yipCmI8jRNZs6aYRzIlWPfgt0GOJMORg
3tDtoVxYKqGCUCLmedtbqAiwqoP5DXB3+ORV9L2GoA48DQ5B65aiHvBONRXzjjlN
zab+R6Cd2PwWJn5f/UHN91pvd38DBOMANJJH0zZoXDE/LhzVx6KgU8CMFusDZZYr
iCBaDJJggzAumEuNaWS8ZBsJzsrfJ5k27jGl+YNXcNadeG2gCshdFT6TR89FjHPs
lpZ0naMyRDGvCUrvIiCanROw+0bXBd6qfb1D2U0JtMA5nUX1uEF7MAEnCKo4LT/5
tZEUdIFLpI75Zc0EWUqUhEfgf97UTrXP7ekevi9VYyF1MqiybY3CeJ+RC2uJKuo6
M8XkmgjBaDgm29qtJcm/D/6WBkxZPADzGKNbboExNXXrlMouXQ5jhTYan4yWuf6N
9NXFKzQTwPsKs9FYHhVjqSe/t9nukAf+0QR5e+al7MeH20g+vtzcEvpQ9lVPIBCQ
cMUew9RLxiCnWpG+dqdlpQHSrlqP5BFwbaEJ2E48hjC+pNDpLFN09uH6Ykn+pQ9T
BoOQ8Ey+QOHpq7o8SHLtDnm788Zfnfi2wNabWfCCwUFLGfJKRawNR+dyx2ALR/H8
DsLXPcXObtnSiBZ3Z8gfFMmk8qke8um0tYqOUTaeHHOADK3gKLL3cTxx6fILqH/1
t4+bAuJfbwIi40znYkfwG5GE4aS4jhf8hH9lIu/LbawW8SvNqTlEJNAbmL0HVBB9
i2fGc3TdK8wroCldSkxT1ilX1gsSS05lj9N+MlmnNKGN5H7oBaS97oxqrF5VNZPA
5Y7fIgLbcADnw1Dx64DKYakX9NDHkyIrvcM5cH3qAMYy9O4IaGNVJOGfIJ7cXmr6
GJEnj3Nsv57Xg0HEnTz5qiEQuhl1ss9Tkpi1A6bki2/5HfCvlsMU88U146M8fT3A
Q6vr/U7rIQBOhmNAqFFtXDtuveFewuLc1CRNwN3S0nOd3h7vqegysw9XT3OcUvdg
xGkM6AkfbHST7pgQUVTPyhRy9chiGF1gZJm6lJ+OL/CaXdRm+c85ySoutzH8wmSR
zOlDEBdjRbMv0S+mz+NTnn5ShRZscJ+cHn5K3KeieHATfVwZQfWRBRXvUg+KWTzp
cXdYEZAH05zhfGSZvakVe/HwOHPs2kvRD6a74srXED9bSpg5Pf8fn++4ztbPF518
rKqgTdUA4eFj5qrHpd8S+SEzRt28jKu9AfXHi83o5sUupOeuwCNMCu7s52+Lyx2z
n+qGoEOU3VbygPgxQt9UT9RJrP5yRowF6RE9m4dfi2D71UIqyQs8ZN0Ijp0UIBc4
kKKsHU7tDHvoy09PyTFmzmbetnvFY7FRkgkFMWBaTAoBb0T7ncaX+Ka7kRvj5O0f
9PVjZRFA749l8Oa1ksa5J+UShw19naHYERAx7NZKIyeFJiFZI0wFAamVcDP7vIRc
zQNXgzsKeUPhhQgX3xXmEXSQ3xrEF39Xn48bOrMUyTHkUWP1o7OskTS3Pj6pHuda
ZPO6Tw06dvIPH4EWMF5zLkTAvi7jOJWhj40EPkvTeoZsPa3owTK4MfpExRMGn2u8
/0MAu3xpNUKAIqoLn2TlFc/Tc0zvM/406CxNCrbBv5sKrNK7VWR3jH0QpyGCSIJC
cDw7COQMetvlpFhqu7iLfq9bXkqAaCtUIwwRZ4p7rxyo7StDZFh5qWRo3/ruPtiC
DulfdJd/mOJ7IuwKo39DGhIPBzsdBmoCgyb3RGfSZwpUOUHi1oFFTVy3StSk6fRK
I/T3Rf6sD3fmC6b3WMXq5u33LTVl+0U/M2CIC+1V146q+RgWx2RsBw8ubnABhRio
Bwd9nUt+XrCQt8y1JMwqNXXYo6PGMhaam7MG2M6NfmaezzSA9YJ+AuUDa6e+9Mz9
20x+Xpow/FAQGMSqmulFELusIlcERUkF64Pc6OybYhjE9uW+zHrsEQsDR5LBXUZ+
2NSjVvKrIvXGr4kSL6N7aZv35CYGToCPY/xCDUMzj42K/Z85cBnnGtmgt6TF9jpM
Rk7anj1p7OJM8X4s6juksApQHsvDfG8VViRBVN2LyuKTu+Hb3/Jr1NHEzCKZNoyA
5HvUe1rRlJ6FdqKeGYo29q2Kn2N6GNG8p2qcwU7ffXciFcq1e3Q3zdEDI+T/NVwS
fZtAsTr+Z9mNhIxIEi1tmhjGyEftGRPvBCci/u2reRZ2p3Vy22YFWEkNGTShiQBr
ev1AE04lgZyD8OOatoKpn+3VffHeBTjhL+llrFxZnL1VSHx7gvxLx7z/b2ZcMIM0
5J1y9C2YX+fxbhI10eNOGxd77DOBdKPLAetuL9u5HlE2cwg/fqBtndF/yVWpsB8m
PmE+0VHMKmW+cy+8BRIcgwxGfMflB5dx/MsfGyPXjaZW3S1dfNQ+EDEsgYe6qg03
cw7rD53ku6JFeQtwP0gcMYvvxuDuiji03gSVvYdLS9PtZzMs0kCzpDnoXGeMMLUj
CdM9bEagOwJPgnxbmLRCAj4ki5otA1QOptT1H9YbNR51Hjz6Uv5B7JPXJ0j87cQv
QwutvYTx/vZCpME02BYNeWnNI2D6+tRqorLut2AamW/DYoDHwyPnic2YcCvGtKBN
iqZJSjPKm0BoB74O3WT9BEUsRzCkHC4wROjENC64bSgzO180vpj6Q6aIbOODrdFk
BIC8JbD0CgFXExbqgWGpRuXh4JQFna4vC1t+Gma2ixF+OSkR1HUywb2YNszZRmY4
0PinbFZvi2JnGlsPLmbTo7eFQpp7cdvme37Az6FIdkHTx0ACSvh3dBmfClqREqXo
QJagj8LAV6I8PYUNzU1SztngP6ecdVPnCHOspjrRvMdMTvH1/9hmtALKvBJ8TrEa
8fpdorUAs1/6//YjBH8YWhj3waTkHfdsLsZ0X1N96g1TXdhPUOIr1VRHDMHmk7n5
kE3kimqxc/DXGghejLlmzxA4GMYs7GeuhQrfvTYOL4M3n5pAqnlCqYWgn7OlABSd
xOAXzHqPV9BeIcPTBCtgiyFypaDfrkJRINe2gmktfvvIm79hcRO4/p78gmAkWkT9
O75teTJYsYe3iqrzlAnQqr2qkxm9RCkviopPx4/QIAad7H8D3kX/h0KeonWSyHFT
DzI/RzevGwdV4rcrlSACY63ywqec3F+4ZYeP7+7/ziNquAmpoK4P5VJt2zgdjuO8
I0P9xrJYH6wMKIMLrVHz884oc4YIUqvcQ3sRsozuvN1qvyJrRyYiOXVSEePxKO07
0JqcJD0VY6waA24vaHoQVUBtNKD+udHhIhO+oFw4vCEgjw4T+PFTBe58pRMDbWue
UQtQI1Eu0hg1FPmqF+KGgr2QGGevopTAGMlZnsNiQqJ4cKtO1yOB1tJAt4eptsVG
ANVtUw7c49mgqXLh0CGdxGlhcPAYSLQ5rV8TnUa65MhcTKGE7JiFnkmrzcYGu93h
/8q4hyctVWS8iev8rLN+Qp9Dct3Sy3pnIsgUBVXjFX/E/u7aeBO5Sk9cUNH1uFDJ
RNvp3xShO955VqtUVmFY1cZtUQY/8hYnUT6sldkoeS7AwZwGhAeMOp3cmuSkAcZY
71eYJBIbEiuEezOl5MJfW2N89jpsN/3NDTD7A165oEOvE+MSyJ18RGDyWQNrMMYr
J8JCsnqRM3ankieLY0hscemD7ic4OxAwPQUVFfamNq+64GO70kkgg3I7W2c95Hjx
MFJ4i7Es7ThbLlP9G9TFOw6W3Nypv7q8DkdMQGFe7Fp2yvJuNd+8y54Z01omcqIh
RBf3cbHZd/dH9QX+7u2bZhHhsZHsCV/eVMPeCNKx1VEFPHUTyxa3u3pJ5Ud9XTHS
RKQK6QFCJwZfJ5PWRz8edPRSpOMmZLZRUt9z2SQqIWYz52E1sATl2+68EtdxikGF
m5wg8PeMIx4S5UpfbgvvClmkzeTT5ID+V4gTdiArTaLudOb7iA6NvMbIQqFil24K
L7Xsy9pfVYHvzB9LLd2UO/CNlvfXO1i9As9IfX0FXD5MvKpJdxCmD5go1/9Fq1rB
uDrBbJ4auNNgOghcmi48IFOgiSOYA2weEVhYQ8SE4h4Bqyg2ZQsVJvWq9rPA/txu
RfU11QNakx4XnfCFDrzCatT8Skp1iTRsIP5b06B9zvluut99J6EGX1B0McpbUms4
DXxV4U3HRpPVJwt6A9Lh2AgkkmTt6h+SmKK6+Y7CnlrL3QthgPUPnc54aG40X7hO
TYZPu39toZELm9QI/GToPqippXZFD/BKY9/D6md5h9h/lUwksqXX9U4C2SxbDMov
sA2txWqlZu18leev3V+FvzHV1Eid6amKULDh6aN+cdT+qXaeVWeIniK8I7grcsJS
kri/SIK3jQJB8mMjzymuGUaXToUu2/+WsnJ/ayDNqYksGMB4Wygx52mZRmw12e6g
bC7zzcMr37GhD+/XD+hwHhs6b/A5ZwQ4EFafP17PonAv9GvEzm0ktn9LAtc1urmQ
N16+QvFIw/n96raltVAFxp2dVnylItTD5W3Bm4+Z1htivgMKrEthCVu2W35IT/yr
3VnPqUaKL3O4PnRG8GwnvDZWEJFIM2ctLYjneioiwoSijEv+T0lmEDtNDPFMBw7a
2VfwqM2kvg+2y4XB8OXukRExamBchox9LfOKj33AsxmszU6jH8bAAXavk1Nxqgdj
ryrUbrAE9XdCXhp9PPl+qHAQg1iyKu+4zseOh9p/pKVSLXyY15ZwnlknR71oRSPj
1tpYA9Gzns47jqjS6kwlXv8b2/fAl4RYzxD+s0+ANBBvoQWjd3aXKBS9JcGZUoEX
1unHMeu5O4Le6D8rLFP6dJFsmMh/tZ9FZu+Qui1fBfwn9DVRvum0ML3EKaB+2OLX
B7pPfLgK8pbSt1aoh23GeR+YS3qia4hvpSClyP8E6hW2O8L7QLvgneBrXthPCzHR
e6Aj+57a3vXRw2wvZOM9NvfBPc2w/LPp4Ejd9lgHxodno1mpKZhCdF1LMMYPmEpy
Ndj7GX7c+o9QEgHo8DWiYKkuOA37mgnOgwiD1T5Ckj5EtsDVDN255/UD2lUzncUy
VSHFSe7+tJmAkwjVClLUvrtA/N7JVwWlgIxFTZMbwCjJO6QRd3uvd06uJaFIY2Eg
ouYE+yBxF4aQnZNdp43CVMv2blY/j4j2qm6KxBtri8RxRy8oZRopaxawr38cAmNI
/2nAqKX1RiSPhnuOVtxM1PsQ8auNdDjnPFtSoXrf7kFZ+VhpgUebGf79PKHcObAT
kxSw9uys7rLnI00m0LZ1AJtKejZjPg4C8RncJr+s3pRis+5UBZV6CpdsvjCC1a7F
K2BrT/iOmmaUg1qP2/+dlnM6Dz6blw7aG/sfl3c9wdPZ4jwgFan+Cgps16dzhM/w
sUve8qPpoNA8VH/LNZh5i5BHFTlgjEAKLkmWspO1jVLckTzR1zaHhCpEaELJJF91
z2iuo6t2DfPhfx+9YUhfatPRfvGLcauWSx7BXHHVKBQ/yhZhGQ8Vh5LtnOQC6Bn4
tn4XpbwWe6mJhplJ418c67uM5kQ8mKcZRdCGrzA0Tn1pYYq+BYKRgSPmHSFuGDdQ
0rJu29sURV7aO6bEUXtbZrQ71voz89kprBipwmTjAgTZixzQhNDbxtlRlw1WfbyI
ewi3CTO7AWjUTuez6QUj1a6gXAiG7e9RpyuqUvETlkUrlD0olFHf/np7uTgAjR34
2amvRDXhSB2WWobAfS+qeFoE29v++McYeZAaPTgPYqLc2XA+KJRzibGLQOIpSxac
9Dwa2jS8/xPwKHuYyLOuJdi5e/oQtPjdocUknJRFA8C3ZWOOWFPNCgkbqsuDk97h
NEKaBLZdgWbdO/SSFpmh21i2YCnOQcT6KmsDDvrp8+QTeedhR/CQfbS+PYN42NG6
4M6w06r3jsBWho9GwzP9EIF+D0sJ4Wiz/iaDAmnD5Fk+BngtZD+xWg2GdYPqstgT
s0U/0Iu2T8Omw/cCfaHOR5k3WZ0NkbW6/iat0aFbxKNBU0taHzk8wz5wpUCd/AHd
hOQrlGGVCdZ/pAOQ3ljArSiFEoYxKp6VScSoSfMC9q/YnMlktNPgamWpyH5vDNRo
V2tQbPAtA/7wyfIkrohR/xHsQsuJ4cm1WLFMLEOkCl+MifUk8/RdRlklJrkpCgdr
SINxVcOvd2v7TMJnv5+9EXxTsXsD8foMxOlJ2oZHqsUFOfNLKWBsmUO41FsCMGJe
0QbjxLJC3ZRxYDzqzct6ZRNMdqbdLDTHtEYEJvEVsIb8JT27VN8NELzVBSSC6p4F
QANpmddHWeQlvY+Y/RfExhDEDoKFeHT3Wc0TflmEOqFmwDX55MIATLAd/Jxj3sQ1
DIuSQCuCIj8Nfcy5DHx2mRwhDbgt58EMbvay41zOi0vqu+hm/X3FXDkeKkP3iXlG
S/YOrGqC47wveaSOojwmJ+7IZFguhcO83YkKXSylfJmqTT+C7il+vRK6dAh5CE7E
kuzG7AqkYfwyJs2IlEU77AzRRz55+CzEj3VhJ/fF1X0fu3ZKyXVvNPDnM3JHnX2V
MWZP/GAIP8v/dsQ+1QbzddAa3KD6czhqQC5/fEHCsYYPd5nC2UDxM6CH5K+LNos9
SpGjVcepGT0scxVonw8IIozUQJlnoOwmS/3eYwCix96vDBCWdHvd0AcharKDqxtD
rAGAYngbqGBjEEq8R2TzR+BMJPxmWcJZ1F4RJTpfQWLH9rwS83Wh8kqscbg/RAJY
vFyXAXAjOtlA+rCqYnj51zx/B7ZSV6/bRVyqDqkBon02i+PpP732sX+UIwpGME7H
U05JaI+t5TOJY9YPqga88IbL0jpNSGB79rEsFaktsKPh5UBNLYQskhBnivieV4pn
zdTkAHwUrS7Ms1Zk4Wv5zVZQuZjRbhgAgY9eFHNQAlIPUaJpYjmBPr6+RO6lsJkh
VjXa3tadDyCcfWkkTIBNM0SEm4BKMgt3LchcVIcbbYFahXIiMeIL812TtvYzWz/f
QgBHIkvhTKZRAYpdPlSehEKgW9xc76VJK8IJZE0wmqIMPqS4ZvF8glp7ji3xeYPS
SGsN1mJJPRHBB53vEG1dCEePMkf2phWq9pILWu9TYM+/2cRvz0AlHmo1KWlzBQyt
oobaKm1vkTfD8IPrlAI4E9lMStzYmEyQH9GCF/AtF5Wlmt/gFraDYEiLBy0Famux
6K6SdVLZKBySr0R8tQi0cgqwvfXBI2bnUVIXxCrZI3DfLm1Bc/K+waUGGp4sUO0B
t7WHUfwkPFp1or8xUcl2o1sokhUxKomXU42CKVFSnUln6h9g4Y6lgsNvUFor3zdZ
6uO3zrf6W63dfs5EDxHvjA4l/+KhGKKUwl+NFl1qOToLoAroSuylAEVK4S3+XlZL
Fhg8r6eCR0Mf9cbozKiI55MYxv6efilxyPT3l/xmmPHhDgvd7PmvcxjVzIDHL5uO
vhgohwY/4wSJJ+pMhJZoqhVLNctN4sS4rvxDX/F3Wl1F8RiSzTIkAULgkNaHi7C7
oHWSIhaL1nhcD1QdXusIublYy017+Zc6hFuvqA4mthZlN0cQCu3koEUBhh7IEXjD
QpxYuIVOnbzUA0AyRHm6bb4X5ro6n9NiQPrWp0T9LtM+9cNOvyYOhot2BA67ZZ3r
1i0lR4E9oLvXGOom8ybUSMl2oIYqUPy/JNSNmHpGCgTggU3lEbxVSUvyj3i9fHXY
Wu/Oqm70emuaXCl50hdg+pqG6n9tIPbM7grWXdkLZ5gp240lUJS9ncjtaZRoNrqY
yeL+cHATkswSdX5jQEiIa0uuOFKKnztLTJugvDUi213BtlDiH2VqW+mcxE/bT/Yd
KJE6d4G65VNLTLS3Kv7HDu1zEu0TSuAZQAZRHFCMEQ3HaSnvuMf+7+vc21Ss8+Xm
NhGWiqPteFXbpVub7R32DoNObcRaYIY93zNCk8lRoKicar5DoXW9iuLfBywUquJd
wAnmSJcKFKASn4GrQS4y6Y3hFn+doH4MALxJawg5xhggVbyWi6tCyxSM8nCGoR6a
bCjFlQTjl7UjPHAeBy1z6011CUWCk+S3jf+xDCYC7eJ3suxC1oRmoUaRQ81GP7IF
6BMjFQsSfmxkOSTda8nwjZLe6oE3jUGp55x+fcZxXY+3Sc46fI/RzhdTDo8EvMgE
wJDbLZf5YaACIuGKHE+JqmyFwYoVutano1XQ4plgN0MUaPYPcO8X6iDRLynEltp6
a5g/eKHEV/I7qz79pLUSkGyUhOiYHCfF6ihhvwXoytQQ5QNMvyw765QYaNxtVxJB
BQVzVDps85o/qwbEfCzpkGEhJifGYpD0etcyD4jOQ7kOH0r5s+XqLvGCoja+j1Fc
eANHN9CcU9UuXekoRo27aNXptVT7AcmrZtYBmO8Rka8BGuEQ9jawlKdvVQeTtJ17
wws+K2Rgp20XPTtkF/9Bvv/8WCNcn9B0spsluTGNAVPBLkXKLbEnF1c+psd6koGB
qKu+1UL7L28gXgEJ3yR3uvglmT3fQSovtmajf9rxXGyE4PG8vuv2dS+DZReHBHop
t3e72qd/hmNSyVwJIKj2sWAz+M+T5GJdpT9U4FE5lHx/POjkNaQB5bcCfX9FxR3S
lU8Uy1dAZF3uPNGM6jwuSCB+8+FMI0s4JsCA/7/Lv+M2vakQ1QHR4/ddJvFinhq+
aTU7e/SL4waL7KiTkHGAe5U/t+M650kagg0yXLkQqe7Uz49UjfNDcXXkHXyBgWhd
/0PD3B+AJXcx6jGGoEzodhmRuNDPxZDon+hWlluYf/uYC3Vkx/f13e+W8riBJExi
9PV+tBv83p4WhRJNCzIonY/a/nM5Lp/5qw3kTIe8X39y5f9sNBgtiQlSaodsbHnS
DlPH2MiUKEZfVw7VMa3gx4c8n8LKJ4gKZu1u6kWXAyFwpc+tyZ6PBtI/VAqWYBRH
/VPSmLbtfgoLZSCFuxcdg5UV7dS8O2LVAAfyAXs6oKITMG525sLj3LxIHCdvF+In
QAgptZhHDIJFKKMgdjclRVFM6ZtEZfnGTXF2fZRcicCoQalsodhDC2JBZGmZoqFU
wRTNqzSQeQy899fC2piyJvKxdPlTC/3CgwGS2mdLqBNva6GoEAsv+myYFjtWiYT7
skCsrpmNN6/64rHj8P5OsPOtnR9q827PnaFJSm/91ewGoaqyJuksrm/9mfByQ+sX
1yWs6VCE4h0zZ480B+U7hlqkEj7lY29ZjFf1jrTN69XcdOODJ/7aximifra9P4Ma
2iHfZ2KI+C/z8KAy+owgFwhVyQ1okYkdhfKXZSaVFpEUiF9nWuF42hWKjiT16h6t
uSpI0vz+KyMpUjJkeW0qr9p46zojqVcq0EThqg3NZA100F+HItB6wu3TzTtU43zy
nhZHgkK6bn/+LswoKd+MMz/5Sr22NJGHl/cJ8K3rs3tebxsCuWH/KUROdzRYuQYT
yGt3BsLiJKPaKqNmS2+fO2qmnXzcG5gGRC3cTIofqvg6Ptv889iGngdUNK45yuvI
Q1R8GuEk/Pfg5+ox4lixTybIYTx7U5d+mMMvU9s2+uRdh8sQ8xlPGrMFuU8GQ1e4
Bu4F3kQALaIwz9rqSVil67pzD/CqCNG+Yq2ggOndOsqVoCt/JxEwh679tKrJ1Nqc
DL/vVZwIKzoJbYrYi5LnJLYRlf0l7IhprxhiOVgZi8xmHQcNoxySKLc/yJ4tfBfV
u+6CLVojtXRled9UZXTTkBRN1z+9ZRSZJCFPGqxwQul10cyMoo+W32LH8quPq3X9
YUR/rJRy2FyEXrpl8XoDe1sbmjI5pdfpkpaeTLUDUj6Lrvpms9cfR79ydDeVX+dN
6rTXna9KqHUBMKDSHcfGwdcCLAAhgAuCi9Y23Il2uS+nh2fatCqw+eS2Rz08WGi9
ZealA9OG8LyeFn1da+GfWaa7rhLwhdnr44njyEChs4hmIsX0B5v2sGSbACkWGFEs
f/MYlj/DQFEw/81Xe3U/wVXUnLJkR7vAAHidjyGWcdwXx2fdBlfgl0yTnjJQLwxe
FsbJAvhQrKh4dxKbstt23rZtHfGFZJtqsbKY9P5GxZ6N+cPtd6vergZZZV9DtOpc
Zkw+DnFm3yVsvPFct+eu8kI7Jp3fjSq37t+B/IGX8/XLpx7sLChMEzPdozmM9EmJ
4/3pVP96hdTkhU44ZHV/llb1S3Y/5psTlmC5N+slXBOfVr7vRHg+qCSwMsXxiawQ
DPraKefigJyMUFEF5GDgQeKzKBNpY2FppmsnJvFa20lCHpxBl4WVNWXPH+Xo7S2E
if2a1uu3mIXVpTicAFChcnIRYis9z98i3k8zCLuplzcmVHslI3XrHspEwG/ig2tt
nct3B2hIu150nIPOuuWIcX63Day59F2/KG5gliQ/EmccS1AiFehMEycH6DH1mEBr
9Md261QSYoY4oQS+NpEzFj7YxrPP/WgLyoM5hRSrDBlYC3z+3Rk7NwAsl/HpsAho
MLM6S2GhxZSpLOUFx09S+o3DkRJOavgP/xn+GeShN5Or3J8IOTUrrdeRpsUD/iyR
0O054afkkWtkJnrwoEuwbKZi//xoX8NJ35xdb1x0RGzRuZdR6KWsVaT78Or+6m4D
PL7lD3K/yD45l6kAMouHGPjVLiq9IcIZhl4+HAIlspqCBZI824PPentxGbYvlPMV
mR39rhI/iDeSWVz2f144tf5Uj4ufNx9Zv4QOO9I284xYJedJKehkypPGnhGrbfNK
f3BocjREezs3+bwn3lLmnCH259sk6MDAfl4/bEN+Tbu36c5zsbFLm3KKkBG2oFs/
MQMIimA8pWpBuNFdnK+R4fHir3AsQkob8IV0GrHNcbpC8jHI2gxHE3s9G2vUMXxg
rdFKxsesoerP1KxoVlpd2yKwP/J7SKBtMRwCXffZ1GM0N3yArQUZtQ8CIpp0G40c
IOEYPP0xnLCIU1sDrCaBguvlYm4ZKauRbSN/lsSRiVaYx1i3GTN1hXmIXTZjJLoG
QECzpMDaxwFdkZEiNbBG7wAYxhQtI75WApLqI2407qhitapF+lweQ/3GJlKK0tGQ
3OjfDIAKqcMQ5lPEI/yh/4IvIRGJDdEn4xRp4YwPnj9lLVI+6hbBBWb1TMt6SS+U
WjUX0uA2hMzj/CeRLqakzlI4DVXpMzKjEoHnFs/tp85q7jXNAaeyb693f2DiqvQl
4ND+3Vhhj4fRPl7MhBUZ6ovGTxWuFTZZS5nd21Qx0a61qIsaSwMLOHW5DZqprbux
X2UbHDtFMBeOM0kAucoFHQUMlysd6CC+D5g7+rjUIny7Pk2oQM3l+LzvyinhafL5
PYUwStTA0TevJAIhhaGtU7+KKaKESgkSx3WfKY0X9wv4U05JyfLj8h6oROnfxq57
9P75LpJoKXGECa5gj7amHpxHM6Wfk/rqm8+z4pLhYooypGczv+1/EIWXpS5fMUEG
THKEbonNZ2lLpk+Zs09fmPb7zD8P8eOC6K4O4SYjt51aStW7mkRUQXNsQO07rGk6
N1kkCrc6vG3UOQUsbzoVhjd/ayTJPfIxk/QleWuvQmll824auMGTvQ1ORGu+org6
UYVHrPAPjIxcc+6CUOmsPUWzRFndLrwR7Dz3/EF1ZkIbrszwpxJSwwOjX6eD1eHa
czOgoz7q99dVsF2hzFeJftlSgbJasLDkgt8uYYF6W2ebdvciq4f8rXx3KFijMEyE
k7Fq8C7a0d9chjcwXRb1Pezxu1CfCHqSH3edbYE2zoKnYtiCkgXlzAtAgE2cucJh
/K6OeuLP905bqJyIap6zLqaXK33YXSCG3/ICweYjCIpy03r+iQz4OQ7i7sCncKzQ
qqtUg60m+in8JMrC6cB7om61/LQeOIvgnGaHXichcOSjobKKDDkFFFGCNRz4Gwdj
koIW5bQt+jbfKEkl92MHxAVWL5TLq45HL35vQh4wpB1DJ/gVm9dWgBB4bS1FIvzz
nseBu+iNaR7uXu3QLNFw459e+jm/S3FN8wvAFZN0CHXEtYjhAivRMRy64OCe17HG
pOEEDq1RI/SMJHT4z6ekGrypAdxhQ1PxCq7ly7T2aehUUfjNFCOdmso72YZAIJSY
3ITvm5Fx5a0H9mayBBiPVbX5CkKsJ5FSJodE2cjo7dA5OgmOsDr3w8B6isRdbRky
sFv20KKF/jSVMf4X3I+iNO1r8LLvpPz0204j2xzu9YCctlcQg8H15UgVATggpF1M
XzasUk0sOPq/bXTEr4+xFvUJqyQCmrVuMSUbvroj+g9R6PwYADcAJcpVG3RNeJfn
heeM339nTZoTPjaTG7cdAQ29gJbIiUsiBHOvL6PJC6HzDDTTthwm8cchw3pFtRnE
wzJRWqVhQWiEG6uMmcSJkyTUlrn/eK2r63P27cgLrdmJZw7bk5dew/BOEJPPfp74
r5m33U3VPqFlbPYfQhL4YR1Qd3fgXQmCOxEBOTYf97OYGGASC8SR5vqhb4OzBVSY
WDmZMA0g3gMLT5h6DyZbWvFbUguemQ/gNcuDe5sZNGuymtr2EU42oho6j5VmFUfj
kqn6+rOv33qHEpgwIZr/0GC/uCeJ4grpLWfiQ1bRpDHVX9WSsIxuex7C2khIREbu
nbd0nvydmVMxN9FZXLVzSm8h0jfeVCBR769jfhWPCvDlMUv/v9GSEDVnGTl0o4z1
r53Mben2rIG9FXvDpC71L3oerTXd+xOnM4zizN/W/p3Po2n9KeCP0eBLUR8Zp80x
DiOVq/he9kAGV0UKDUX0Tc1zrQpaJIpnWf0n7WFSgBG/NaymmZp4j7C3lvqS7UDf
EWgq9eD39gnhQyX/kYgAgK0+2sN0u2AVybCluvyfOH9ZLRvhtZ1W5S7dqhVRiDAi
lC3p9Q1Uhy1MzKWl8rj00lx2LOWYyQWEWmuRBU+N0vi4zB17y8NH3IKUiBYNcmZE
ItIHZ0Jg+bt9UpZmh0hpFDjR9v8eEmUnJE9BBcGePd4KGX6oI0twhCYEBkqzyQCb
nQi+Lq7LFOr2UojMSsXcSXnaH5JkW0K7sxPQORlLxfMMv3kgOeWzM9FNigMM2iLl
RVyhsdXxDvS8NXQWYoR9plLrXW+9RvK73JgIVdVyk4ATsOYCDb/xPI+AkqLGb6G2
UhAOeojaejbSTCNW++gvDoQeAuQmYvYGZhHIdoq/JSnsmO/A4n084KywPtTc3Hrx
mHutrN0XbQgrSc8vUrt+rJwXha+yziwIbnIB/SbjIe6JwISHOwXESavd7VTHitOx
Otp3DA/6Q5HUsBhgTj7uFJ46Tf93HRKgBAhiv5cBBP49+eljdAsVv/7VZFetzIzu
zvNtUtmzFv5jgNHxQKKsc2gVvV6ZDuXdEOuF/HEr0U5S/bCclUEC2+8wOrhIIkO7
IhU08NnerqEvieb4obH+/4Y5fjOHCLQPKPn8y201yx+KTKZxv4+AsJmMSKnnA13r
8D9WQlDce8fRSgB3H7jgUzI14bXzBO/bsB1jUjZWOOFJ0w7tHvDL1UmFT/pNU6LI
S8W02XAYsQXn15cokjKKGY5oiHI3wyF+ObNlMEJxEGnNMHG+Nw2rM7C4Bl/rjujq
71PJP4VIZ04dKhfJi2fBq+HoM+dQbHCeu7GDnSTLyv3ATf6RyLSn2nxOUtrNlhbM
FVhIkkjt3SkF3D2wBzp4C+geed/jDTbL5PL04QATHmy/TryjCb8uso9DHX8fjPo9
LulAW+vHhBu5FMFkdom8tPE9lxM/aq6iFnT743gJ5BcDMJ7LLRY8fTF64e5Da/hu
2tx6onVWbtSs+C3AOV9hbtVUbjbJrCT3//y6rIEE+nyJCBciIRIEGbjMuGg5/3b6
nhDDRTGgpWXrfr6MYiPK3Gy7Js+H+CQB8DOE/oMdyvbRMRswmGq+Uik8Zgwhao75
GLOX1FYOTG+J/yXm4sSdPrcSxR7JXw3QbvvFksfKn/vaBhT7LknUSEHPiOU51gU7
pc0CJkXJ1GRCHPch7Ujbllfc+Vn9oq+Z6SuqbGmyLRxRfpou+am29MlDo4siQNOK
lEGVoCPsM9k02qoBidAdhnT1ti/ma+MSbzYs6iNmb/giZveIPSjmqfaTJhITAAfA
AWuFwA0YxPkH/CG97xVsJ2hE8KdPcIhwKhwcPlNzfYjp8P02oe72FcjF9IG/K+wm
1O2nROnIGEdml7F3jxat9d625Ynj425FO+ArmEVo6hJh8SZVY7Sc2m7g3oZ7MCzw
cZSReFs7c+47waM/xTcxlEFpikk09VopN1fYtNkf8JpSyyNAQJVL/cR3zPs/rQxr
15qA+girBtRYoXR46JnTMkzBxTJAq8HHPURvxLDiyRf+pSh+RZ0ZOfsPzz1wv7kx
1uH/NTzAKbe6aK2QHUmKIKDcRsBt30iGRVwGwDokBE5u/48HHVheHal+BjBTpJW3
7axcxBmQ6oGP540dJWsj2hpaecMdbhr98ktNPhEofnwUG+MsX79CJuEVYHOOdJ3e
hBEbu2D+hn9MIJqdm5mGMS4AHHZJD7Y8MnEosPD1MjuJFtOZ/ntu674RgeIBXH3f
3p25hc9R5HizBCzFzzyZUqB5lV/VyGXvwZvuaXcykAqppFs4hWluf3m2V547S0Xl
Ung696IsysL42ZdNN1CC5D0fBe3mbEjiKFrRyCrcSw/Z8YPrkbiiI2SPfC73lstc
JM0DQ/A7WqOEmrfrzJfCGWlFlrqhG8bYQvyRJESi916B0pwktZ6Ivzwl0s5phdVz
00A0N1H9KwVqXnqhEOlvkur2vmW9zR3ioXchWuKzTaGqpaH0NojDzYjyAgNXXm1+
w5YXjzhYtIVLJyu6qhS8gBOOh/1AcdSePXREPXSUsgbRQ/idrcH442FCI6fnz+J7
v1ZwKMaGVic8i7LUxjbdvkLeOmjlvCP+FffzYQsExdXRnmjBF9SuGD39RNL5e8dB
XuOowQL1f+tDq8XoFzHTVHSftv0nIH1KPCNPYC92c45g6d+NI5WJqUvSbgu+DpFX
+toLX6CqhI1JjvV+iUqgNXG/LMiyCUKGm7iZwuP58lWbOM/ukVmuOg4eGC901+dP
0M9UM/8W4Nl75c55GvzfBEbzCPWSeOCkoUpHVKWEwXdKPip2gfbAmj1T1yrExtOJ
T1y+9tUoA0W6rFIIyJs7NkK7HgN5XS7NB7BO9LUrBoEMGeSMeE0WlXof6XoeNdl9
ZqtkM3UGmqEMNWaTXFthYCxS+Wxiqqt03Ee1tieHMOlZCW1/7O3l9kAIKJeDpK+5
wUE/ZZl8TAR//CDEV43XAI/TvyRasU1g2wmaT3LmrJQp2OyRPZffkSvhagRo9LnU
bNAVv05wOmJx66yiMxfdrwvGu1k/u0rJLmteYdfwQaOqR5/DgSlBbesfPFhqz8ES
GAm0UDZ7QBwhr8luNwvTYH69uXN2ddXvXVLI1QXcUrLCtUBilquUg8umS4q/8rXP
zs22IbmTaHbEvos2je0cpQwmA36RRg0A2fayVkuwE/glIWKblhyKPibAvupUEja+
wtOmWa8Y9DZ0skyPNp2kEPC2KLdWKyb3qFyo0dyWSmvVFFqo3xByxz3ZxXOPA+Cv
AMXOvnpD9LQpH7XxpqNPFP5CCMlpOvhUXN57TD8gANVaWAD8ZDBbydVzQ+cFKu4o
MxeiR+AtmRGSAzf8oqmMJN/GUngC0D4MCOuJyOnrDSLcB8NYImJ3L9gGpEdG/Ekg
ykOfJwrlKA1TIYCTSBMu7KiO5Z/r5QUi81jWO+UIHB9Pefok5m+DqZ9iIcGzBLYf
0/Wdl5/5kH4GgPtXr5Mz8KA8WEZU/+i9eh65GTQuhzgEoYvV86H/zQMzeYNaUTDH
ZZ/zNp//gjv4nXUbqlrHdyfXRP81Hb7Gtf9AWeZQlgaRTAq6kf4J0f5sNGcSnXj+
vXi6/3wdu46+sSnZsIogEMa8/Ostf0qkE0ZukPyIC+I2ux4auc1CUNRgW5CwHz1f
nuU5YVTc3ebTbWgTxBzWvaE0lp1XuyxZ2qaC4PulFCCRMtBNfi4Y9GCNWkyFj0yu
ASiwppOiosdWnshzMusiug/W+fg7WKHaPwsx92d3idIlf/nrNl07FzAxEdxVFhIk
3NNafEqDN5c8fglqXmbMaX0oQxlBBSszGIVZ0INrR9PX4gLGV/kArMQo8oaQejci
/rlMFp+t8rjt0rbQJYmuwJ3B6DQ1x6U9fXP5r48RvY1yA2N5yjDDXXCYMYIOGuLN
ZdZKQnnjb8Vuv+rM8u5/bQrP7GmDuwLx//JDmkfRvq+YGsQN3WteKItRJlnwKuK7
3Mw4x3cAD+OW4hgHeTMx9q0X1aEHFo3cw3MNMP4bwtQ00gN0E4PTM61jzL4nywW0
BcAoanOMJGCIcCaqOvczP1bGg3tHuAhjlaKTMuHzANzQML6U7dwyCrVIhFrXn/gI
Bt/ZlWve7weFmSS5p5uX4GKzOBgfRKqJLTFoXhyu7ac50rHien7/jCTyVii0cLHa
YXNNq0B+y1bD90rA7cXqqfHhT59uD6rGpOp0pqbvG/2xVVe981qZQctaG3zEwlRO
I2eZ7czHTTiLfVfeHE27NJtOIZdIetgzTLbbnsjreWJEOKkTarSsEED3UmqN/rur
fQeuwMJjptg/jMxJoL1Y2maFcu8CfGvpGG3AsCMomDMTQVAgl/vp6gWJCrFrZA0t
s9oxRDnLqjmXsTxkzniI1d+z8KVndaaonLefmoQgK+StupMlmalVwnn9jOk1OCKV
dswCxB04RfyKdph6Q0vbsT8bdl4TiWSRZx2NyYA7ftgZ4EG2Ta+yxwgRSH+GWi1S
ynuVQP/cs/ZYumQcMsPEL+fb8Y8ia8IcvmhILRLidKOiLMyGp9p1S9W7zhZQIc2a
V4sR0YtaoiaOdA1J2fW6qZ5PlW8/AsOnZh1XSX+zZgGAEMaY5ZkZSl9n21riuFtB
epgp2kBD1AmIs7TjQNGb8yL4Ic+VV5xpJAwBvoXdEGNqrLM8vT2nrnw2bDtObWPe
pBT3UbxoiCr4DT391XD9B8kRrMcbPsK4gQWJYcYRCcrzDX3r5yM4hCwzmeaMxE8D
u9jLkFvj2JcdjiuMFHQ/nZAy88L6KIcZzQwr7SWR9g/egUsHHCsitR0KLwN+A7yY
ntKYQtFra8Uq5TL3bdl3Ws+8c4uhIjrfARJ/qNQN/dIOy+uDdP5edGBjafigv7Kt
KOp90zlqvI8GjFFuX0HFc7sgetftMZv9Xy9vbRuKRzRr2/Cg9+L3/Cbblm4oyXZ9
nzEfysH3QiyqijqZuB8UixfwXQfgXikj4E180ZGjusbzY6buvUzUvtEfBbw38zrp
SOikkP4e7z4ApFNIlU3ofNC/tBRhmHmLk2W9pGWh1WSPF/zd+7hfj9QmnubO/Ijs
CqGlQvgeyrfo/VifDF3v99sFRhRo+qTXbtNTKXwcYA0FiLyHLP6+Gto2YEzSZ2W/
vXFRxm+NjmAuy5vgvV4twwA9W8N+ML1HKIiT5gyBZ5pjzdIbHCqhnH9gv/0iiIxt
2ftCvAxtWKsS7dQTVO/lcOfa66ec3digt6za3Hh2XDfSr6r0Qx1prla8zPEJo6Rf
x4QFNc831PP70FybQEcehum5XiQqez3/AZ4d/gynzF3Zd7613DzIx4T/S2L8A0/N
MOLmHtG/17hs85jZYZMYhuXBXN8Y7oFSDwHMbw5iyNMrQ42bpuye9k/Chbp+93B0
i++Xao0Jrp9nmp0fo7yZJgy9R1xTBSWHSwj1efDtFtHekAH/sDgRV9L1E3ErgQNX
Tbm7I1zkCTC8ERkcnQFwXOxxpKTpLXgs7YyoaSY1QFIBnna4We3A0qxJ8gjwoRD8
PGNv/jpDHIz+tHfkkX9PV5h5RsWbdVRnDzOg0aTGNrAVpuhAfiL6nkom3YrqfUER
PBo6DiDLUvOPoQcETfmu6uT6F/JA0KPqP/tgF1TGqwF0LFOYSLCXlzGo+NhkBllR
dbMSUE0yRj9iW7FkkYT7/T42z9pIeYF2PngIweDd3iyhMnYAj5gxkJGGbcNHRpps
qKdyFa6XDxDAi95Go9yoEIUNU1hp/G/CCn5AxKe2VJV69RE3KU2S+3hiCI/2QzgN
ONF9RAysEWzL6g/STBavaorzG9HpmND6Uf+TlHlsCqA7/zou1S6F8ilyoi9l8uX2
ZpcjxpASoQQ2LVfYz+RWDEtCgOXwkTwdVLLtWpiKsSwbsMU9ae/RJNG3ePnk17u/
wmXXazUs7Uv4f8o8YfEec7KrNgB8vJ64RHN2E/LAfpC35eq0lynknkQUXGZvk7oA
8AFhQI59D2HFTkLxObPfS7MRqRiwB0Q/FB5FLsgPEPTwszTC3PIX+K2R+SPW1y7X
JAEjLjujT6XfKzPLQDgDcNUZsnr5psXtYU2HTx5Big1PZGJ55aoWko0OqGrzMd/x
mPTVkEzNAIcdAl33IrXo2vFkyVdqneUgju3YPX29isuhf5S1nxI/00jg+TwR5Wco
FYnnpL0p5fPpR3qUPL1p7DGpZNeg3tXZrxhKM4ILxx0VvXfk6tUwJp7e3P+huxhn
woo62z6fRpcgW0Di0tvTRnTOvHeQMAL5CzVpETZpNcu1k8xTqSJp4L036bv7gGSF
fGSGfxiJNNfXxxzB+99NY+7Brp4U9cc7iqCXVuXQeKH0IPG+KjklP/wvcPi0ib7N
2ov+bqoY9bPZV19O1RkruuXNmrktqDWb0E0a/wCFh3blA4BK1e3GXeWJVgoITSJY
GIu41k312Qw1ZOHezdS3lTc9vPtruItRlMtDSl0Pii40AxBwFXaGhWicIoELrdb5
RXYwIXuLFN/pSUhvVIolla944MRR03WjY/T88lSPWRaNkPSyCw5iWh+Y5KMWewhd
m6mFemAahahZN1ssqvhgVBD9U1d1N9av2ozn2cJ6Q1rxrEyIMC8rQfwR7tKHH3e4
jgGu602SBI5aJxyHK58ZP5xSAHQAyMoncX10Cxgbwr5+1F/z0vjq78qtf2FOs9xR
I5n/RxqRDchzQng0Nb7tupcI24JHYCONatnVrjZ1c1uge+HZkSyE9Nq+2ydJi2rB
tGKrmAlzOqiiXbRFpmLPXmiWRHt7Kmy8658mEXbIrifCpCt2NvuMUR6MPyIUS9QS
Et1b9OQmfo97j5jNxalJNXNd0vGG/NGkmFsiqAMiedg7RGOdA89s6wAbT7Z50cTT
ufD0/Si6KrUAjAunUI+tOyPd2LOrWxbTJ1pJhA+9locbI1f+GFP7gbtutW4ye7ds
7vWKTCGsHGvXrIt8ibZo/DYWBVt1f4cemALGB+WDHHkl7RkjsEYRkAO3ay1V4jdw
s7KxfdPIs0AddBP8wuWp0f0lctmKQM+PFELuIHoJAUomjaRthOpl+QiugK1UBHl1
redR4IUCsOMNikASlTjBbW40HA4aEVVm0EA7sDAcmTj40ySpGbJwchC7xasSi8+c
SboqX1Yz7H/VfIDEOu0MlamUw24nW6cuireOU1muvvfrKx2Iey4jnBMgaI4RJaEV
XMNBG0VM7oJS1s29gLqMao2SPfCxtN4q+vnfGJJjPG750Ms+GHtcJVRdNWehsfMy
9ZAfQRWGJeYFUWituDeRgEzrKVNcwBLGT8LtTnCDAwkzn9+oGsC6MjD+9q3aK7x0
sAo9StXU3V/TamW+ayTRUSxwxy+uMHaVqQJeaVITnldzGNf3qE5Nvc+NjMHgdzrR
wE3mLOWaW9pCgIIZ4zJwSNGuVd4b8GRpYbVB3A16lSnYSyqSFbhQd2XLWLdOxLX+
kCGA2MC+vnuUpAYknPbOa6T5tiELn7DOGHiSqaKWxpdd7hoVCZ02bVGvX7do6mMc
bGa29DCSD6XSk/mUbsUanv5RO8OdcMT1OAVlTkcLIPhrVOZxq8h+y602EDzK4u5l
EaAKVt5nZKNmU84Qd0wjkdxpsR/foaBC/PB58t87snDAr0OEWgirtSW8dg4oaWZf
x4JwvFn3F6YZ/oVay7bFLQLXxxCKCnkFvPWpD4jM/IjF2DU3Hsj2Re3VHunVnHfY
vlMcIAvuyMOpb9XFdJDXJI7p+Foe3Q9Ejs31mxgyaId2+82siz2jegh+eEad2BSY
EYrofgAtUktWblkrkFGutaNZqlMDBu7v5IpihYd2+yMn11b19PmcFrqvC37uJk6u
AiNMyGdYg2ewk0K3kTkWur8cmbwDVjvmhCxTlfexVqiSAWiGbYtRx5NNr/dY/GVA
xAkFc8/BtkM0RQkVOmrMY2CXyOc/ocZ9dXiwHqabHi+K6/m46RMlHNau/Zq3yKDO
QE+9HCdBGNSaKGEwvRLm8ZuJezQN8KCi10Z1X7PO2O+79A+eDl2RoGWR5/BDpjI0
u2xjdo4sErbtwIetSA6FnHUbb24/ubWldp0T8ZVd2xbdFhEbOZpQCCJc6CGChY3f
BTfV+Hi7U9+apV3PaYFgrklqXXSvEFrqUe04ynGeNqvdZVmLmpTXIX+PIwGyQSy6
7awow1pAP3R0OW0Z2FKwnmmXJHvR1ZsY9wThnUbcZJk1y+inZWf2+VObY0Hav46x
mvPEiSV9m/+J5PRi/x4jX24fZO3S9HI+awsH+9wfH5A8WRcYBuCC+qZeg61PFSzU
jh7W5m01hRBdRRYljTGxUA4yoz5EXnSw/mkSJ2CL/anzjp73fM90eh0ULEtZfXCu
v0D9d5FAnxYz73wtrYj3ji2WbG/RlfqWpPex8+XtKmrVoJmHgHVnNWMpws22lac/
8xragii0czKq1EU/ZxLQHbwkg829DyqfopQrh9nP3G2fpCdypTBGlH6NxPW+AWRB
u+7WFAix38vDOPW1rg4Gj4Bk2pX8FQ/H68Mo7ApUv99edSRxn4JpuVKMKRS+fRca
GYvyNQatA/Exo9rrL96EdlBBKT8afRTJESEWK0qbGE3sMxEhKSBULj90ScE02kTR
vLwgl6oY72w0V8dHzVhiAKGwH+7Ys5Mruo5zsSj4Wj8qv7oQB74oud0so0lAHEP4
hjeCyK0wW4dJCsY45t7Mx0R5No5IN2TVURAjnT+aGVRp4xF8uA9ctHmAIRdP/bBo
COzfBvhN4ffcIlhm42hw8tsElImJF9PDFOvayIkjeAE7aGC4cLenu9O58rx3jKbs
ToaH1JeHl941WVAVE+l9qxbS3yVSFtmWSeocPMhO0DGyPBUofBI9ZQXohHOLNccz
GPVQUJWf91gA3DHrqTHWSH0l1ui+Hcj/WUEYgOeEwP5t7K6okG9+7VjiBt+BPoiC
cxcBflzh8eyyQOj4E6BTsbscbBSNWQDUjcxkJHI3jSVDBbF+l4CWJnzyvWQPq+hY
xsDfwgEAYuhNzWZoB/HoYL6rmJJXQG5n8i65NUKAX7Av7fgHOzFG76YhZyH4n2qY
R+1QNcH/viJEW71+LZSLA/litVJC+5vXpAk2mR8pR+4EqekXKyb6mKSIZ7m5Nya3
5kC4WQBXjkOi6zcECEtfdxkyP6A1QLqjgavJSnO5A4GHQYDyWj1mVBDMUtGm9EN8
B8oTIc8/B/OvJoJxtX1ig0mOxC+ITs4c3XaiKpzsVHNyEgwZ9iZiIP9NexflDqxz
Kpzy+LK2lRQVMt4qra7MQvbXc61/1FLl3p6dX8LGI9+jZr04YnlcajP4DknLB+0A
s8k/58UtqdoD+dTDNNDYZAL/R9/4AXS2w3CbnUeyLPqmZf4uSxZWF9PR77IcjYM8
iD5RIMyqsMkDPCxTCmxAs5gNRvqYzzokGgwOqwJEWWQW8XdCmQrfWUkdoarnpHlU
TwOgcSS4dOCUaJ+eHzMSjMrNA26hWTb8vpRNpnc/hcB8B9RNy/TAZnXqU6yy8oJx
jeDAg8AB2yRz9OKj9kOrTMsel7nwrlXmR35d41Q2CLZJgfgkfuOFewGXGVM1Of0Z
gO7Ovhiu/hUe+fmcbYzOVZyI238WLaYGS592klBaXKo+My6xWMCFpxhIY9Vajzuy
aXqVYXScgSoe5yQsw1nFUGuxePuXVfwKPXakAHWPxsdpa1F+d5m+jK+SAM7BjOeo
uAnxNamRQHmUAZOJ9n8E/9HwyuGEWBpoNKxU2+tBxNwRM94wgzKVTw7mEpJnLDhl
9yUiooL5FnbsLE/QadgahI9UrRT4pKEol67jt1GuCtp6KOegpLcm9rw7tOmOPPnL
4ZykZAKOFkDy87uDLY/8vqel+VURP9atANX8glgZ4OteivfCxBn1z/XNcVrXA6EK
XfysSuU2Ebw785goz3Al/t9Sclq9frtEZjzXtHP6/Hrnzbyfazp09RCjqOvSx2Ce
pw/xHi9o/RiLmepJhbfLMbdkXxp0UGeba2tbSAsuCgAW7HoHSImf6j/4RLzuZEZp
ZqYZ/VcFfXJdNqshVjJFHGHvkldAsCn/MjpIkLBg2XxGVrJWX/uwcvBXRjLQnSbg
3kHX98ZjUhAW0dFwmsrU29SZIZn2TjJ3KGu/lUmcuar4neVPPJ9eeIhqh6oQVIGu
UYFjqS64Ph6SeEzDG3Ugq5vNdsq1wUCJWFDWhpmEJDSbZia211/IzeVp0I+HxSxy
LlsCIGQJeE1suS64Sp2W79I2DCvH22CnFA5ZwsFzbz7WSk8uVePEkAo4hsCY8xgZ
hc/F90QQOS1nbEQ/I2g+5zCmJYvKdNuC0BquUH8iWS+EGPjYNGQXNgZbHGxfOx5C
JAEpPC4irqp5Eutw69M7X4fxI/lPIB6P8h0XKhHQnMT6Vw7GOMantRmArT5U/xJf
9rRCYbm5ELqBXlq3QW4OddJR/zhkLpsJs8qC+ZKOLVvOlKR1qp9HNK6hCaTp1X9S
ofvpp7ju2MkVdlzYBR+9gsUZ7dQc9I70KwGht4qkJ0oKl9NeBY2vdYiXt85gpcQ9
PPGZhY0cm+l9N4hb70UP+gXA6kPFrhAP0kbJLqHwAcAyPQVremlGLyknG8Z2AYEN
isAuzcS3KptwyLxcMpt3L3Ywoa0kuP6JgdAa5ZSbYSOddUlEODczHircb3wYI7Qn
eSOdmjR3uHVlREQwVck7BwbHaPHV4eTPbegjFTA8e0AN1fSYhJTJIF5rVfpfrTTx
SkvR2xaiRXMYMlFOJJsDLygiNGwsyaFUhV+uxvCErtHcHWgr93f383DI1Dh2sHRH
ENhbiG3ES2Xqe1Ve/luImHa5u4UThnHuIXF98bmga9ES6r6lUxvaISxeQjKAqhEr
bT+1r5yqJTFBpV4SugojSlQ2FGjDLWn9ntl4E+U/cbKNUxgSQxSQOn1L03pqnbef
yE/kvo2h5daMn0UPL3djTWmmkbg9waW5TKrLy9gqop1HZaBuNKxhSXPlduSulOvR
fW15bDFxYAYr+lm5uxuv5LE9pwY/CMJQCMFgkt1bYP26hpUyi+4Kn70v7OsoAT/r
abjWPK7HVM4RWJpeZDX0Bi6cLlWUX91hExqbohFbeEhHGr8nBI10ocIHenGqXR+G
7wjMZ3Jlb8JaeZ0pWAgw06q0sE8eTnUZ6VRo+90cEbGm3z52s3099Cx2Qp0SqgHG
cyn5u2N+Oiz4FWJKZcCR8YR+Gkkl+Ipe7KhAZlVyqLOPxY+nfqfHfDfr+sbcbScc
urOeGXyEkHVTfxVfY8Hkz5TkIJxYaFexses/o9no30tp/APNo2SFLgRuivdi8+Bq
PvJWOEoG1spP+we0/ZQjm2nLNR/X9m6nttQiiAbzojjVgP/g25s+cCeVXQTM9/J3
LMcIHmtK5N9jD+p0gG5hpQ9mHTP/n3HmLaL6Ly89UzI8Y1cZUNfGcJBUJKPPNtrh
Ybx3bBDjetMshGgM5TKrInqgzfJtA6ot969iNU6WgAknfNqBUqlcYOkaiifbygwR
KenHx91rn3CO57FL6HMB0bwPPfyXjeHmqhZPKIq8mxTXlC4hus14R0v2i/7+0Rw4
qkzs5/EHMtwzmvzj8MIAhdCnLuJuFM60tYspovQNPtiRUIiYjL+jSHxTOs0kz6PN
PFIWf+EHPYjSLm1qnCRChDQhXIW4zF0ebnBV4f9OsbxRuXwGg3ps1lC+c65nIVti
juYFyci+2NbeYdJaMO77gdV+VPPgMItpUxuV0sCVKLZC8rh9mwnEKHt4GXlx42K8
0yq27HHruN0tw3z/DLacN53mJXgNtys8dXoiT4W+nfecMqhpRJyoy17ZvqADkJM8
MHhyjeG6COREqPBZsl9RhrteF76eAjy+rUrQ1MS6KNi21dVH5kFi27s60tJWRNL2
FdMAukSCyWvU0H5wx5Z9QomS8wS7KFiEzp7v3wdEFbdp7fg01CnEx5way4BN8RJf
n4ZWTeOqkeAEX0hkhj7S/Yfqoo8TCwbLbkOATN9RcZK8ulzUrpviSONeecIJhq7e
0GRocLPBU3CummEsBtJf0cmqNsPejNoyxuu4/KUalYVsoDXlFJMUTSKPCS5QeZIA
v3Igk5OgZLSbGtfIz8wnOB7VVeUG+EAO3iqx1WLXXOL6+/qMXr7YDnWHSTBP8sZi
KtfPMdrvjDconFRFnEHcVX/rBoRTsy01h3FmiPC+IoqoBmzLUsjpHLLXHSPmmZMH
/uj1VmhSlq1E7hfRpgzM0yfWx0ChZQPQpc+NxEQLI/EpOoVGhyIlNgt8vVtOTs6/
jfqkckrk5Rek7eDMEPZzAl9rpg0YlQtfwgkf8hfKlzF2PhSunD76Ir9skm67HJiS
Eoz4Y8iN/aMxM9ewtAW+2bGzUR+Q81vPLkLY24wdscgacznTv6eQzM8+OOc5iZ4x
V3YW41xwBxEQUKeaXrvdXGegYl3pe58//i5sufDgDRMXhqGCBWqFgY/8l00oQASJ
/GpKrVREUtJ4SAU/xbUpg6ku7uvliG9tPrSFFJXaH05MJGBr3ig65pQwCqXI0bX5
NzwCnQxMPXpqrR2+geqqzxcGtCtC52uN8TMAx5Ch+YRXQHfdAGNv7ig63RJIGhGy
JZD/tsrA1wBFau/zhtwFJNR8veW+/ijnouTuPs5nErd2/UOgxIOodvSVpv4OBycj
4wzVUkA5VvT/eBbKEYr2TEQeG7AxQh1kIDBfbGpJoRxi6bQwCjowA9aCW79NegC2
axx2Qq4/gIHRZSgbHUEcIZgitOx305s1vrX7zINY0tM3/uOau53DvfzDBNvQXtM1
0lzQlMZralYYiQ7YbiZLb06HT06YujsyzJ6hUf4yFG4qwxciU6dsJHxJPmCPLL9o
UjW4HT9XQNJMamZo0uKnJIgZKcyjRz7KGDgKpXvpqO8hRUsUr82DS8+Bx05x9qcF
IdpZMNR9tNJNtay9hDVYkjpKFBdSMmmPpHhCEeKe4G9O2ZubjBgkipPuanZIzuc8
PGGHc2l/d71ZL7tJPHOZzKZ/oQsKz4/fQSAhMZ/4W2SD3HJTgm6Jgm/Wa1adi/lO
6wC1MjRYpsOoOf4/sY8KSBCc1qKnJq9tUgCf7r6LBlv/SMhHK4DUD58DBMXvWO6f
NdAr9fjWrx6hq2jbBAHq39FU3vKRz/LeU8Ny9E9vfWiC3JOYzgKiUmr5+SCquj2q
XIp+9iVJ22UkQ0ZCWUKiDu6jHCTyQpzBhrnqQMCL/XFq0MrSZUkSSw061XbJGxO9
mmwkTtAfsqWYZMNFur0vvOlK8oCW8q9HqcaiSa9gq+a9s6bv68P1GNUFwzc7HwML
JkfXs+bcl7RD2QyWru7YHP+NzQ/DuMo4ZnJvZnfBf6x6cGauL9kbx8yuytvzXN/y
nhXxt30cjkv28gIsKJy2+2QHSu4KYGQe6uRDImj3m6QeuvQSq+97UXjshcM9fWvW
RJiQnxs4rmP2lwl0OsYMo/OAIi+NLIxlSE+3o4wS9TQTQfteeY5XkN/Y67wheVMd
RKnAwN+fnCm/alM+l82g6RwulT1j2wtzibPRzF0e/CnKxofBsKMs47HJVkYHHDr3
sI9GuUQqop/WWdB9hQvAy/+vrNK++v+DJlAldLklGsmc+pdRUdCfcJV4s0LyW2Xx
XGbD5H4T4bw2JLt8Fr/NeOMR0sX/KXvzHgXDz9/+scN7QqeLHIdLwbNhyX0YOmkW
sGfrHaEXx1hPgN2pli3sMs274sBT9d0147FsYbnf2gSkSjoe+00tzi+mi1QTPw+w
mOZ61HUQDKgPEuJ5u7wmCn9nIlhWFf7PiV8qu2nXuQBwAbOxMUDonTB1FH3/4aIG
Q9TsjPfrB+mPy5rz0MnXs1/z8PeD6U1EWnYYo/7YBg3PnNkY6D7RsiR4/P3rDP++
oA79KsEB0ub/YSN6QNsFSX+Hf+qjya6Y06aKvRj/OEz43ay5V9BOhzsw8x3SeZwS
THTHLHeCL0IDZ43y0ngQg8jcPEO77bulHLmwYSHmgG7QUDgLQQrVTuh4k+ANnjul
OkrTToJd4s4dBcga/h0z1TuZsIfh7GFwfpAQQa65EYA/7s5F80gcCv8/TXjHnIiu
hsdgF0aDiwyqWxgnEftW9KfbofjiQth9Mm4nxR4hsJBzCVXwS7eJBbLOxMUlRrvA
LijnxJHU1+IMoacyCJB34/5tGvD/8IupKacGGEOvdfVBIiv6TscvzrgCaDDxwzX6
AwCIr5xY0b0ZRIVwpn0fUi7RpR3SZsMYKZDTfo+CMqdpaEn4v4mYPqZOw6ocTLB1
u4dfPW/vjfKMdXfJw+zxYkZ8DU+kytLz1b/WCoz73ywNt6mgtP94gTtzRT/yQUvo
6Q3kacsgQtqIY1fs0qXWy8FGGu7bK9H8rvv9N7GB9UPeYL6SkMNyhNe0rYxbVEaZ
iwsATqMdLYzqS2w9O1E9QQCx6jqdDgGpgNJ9cEACMluicnNJJEglreV3f6tfdzvi
F9cdi3SyF8dzQicQDM4wR3qyHBBRDHQQsWUyfw48i9LSYtrncOp5p89388OOJ9fT
9oD9gQRnfKgvGcykYykpkWgOYcX87sctMYWUgEk47i1IlmVD2xsb6dusbKpYfI0B
2V+ZM4inF8C67zfLpEY/2Y/RgYQI4LvEPvdBQ8uI/RssUjjaggIpiJIyTrefDAbx
youdmZrIpSq1wcFFd6w52QQZNpnlcKKHhz4xWlv1J5oO6zEhczgDksM3gbzbC1WH
qrog6Z+LLOEfIXWVaS+ALLqMV+9ox1MoB1Y+Ql4Fqsf0QHWEC0bZhDPaCkkw4JeS
OEil8a2BJJMt0lYMAFqImM9qKi/hp7ASHX9Ca6ZOxD7mLV5zMuujuZpz+agYcxL/
gZr8zpy/Xpqe1C5K7JLgzdZS9RCCBFSnWIejg7cwQwPv5P1XIDonR4CoBZwfW/d4
c7MMD3/3V1UsfOdGCf2FW1UM19CfEx1d1HwGOlJpbZbygh/++rlIwDDEGbgJsWVu
tOBJgFU7QZrlONCtsgUdYUiEyAlqoWt0Z+6yjrsFLzqjTdhFB9MJL8xuYzmEhjR5
qwyJZzEf0fxGUMln/YupCMkpyM1J5gZkp/P4yDgA45q9y9kXTMlLWVgZ4CoMGfzs
Vknc/iy+IfuURXl/IGlXe1WlrmWb1srIP4t+JBC6Hs5nozK7sxllCkqogiq2DrGU
6fx85NuVz1mM022dBo4WnQzJet1AE9KipBHuYK0orLBJpoEMN1otJwPqHnAqnL8f
EPWifVJR8LZOuLan3gBztMN2RoM3i0E5rxF0s+rBWIQoSlRw4UGS5Il3Zxf0HaOU
ZikVuDE/da/gP9brMDhhRwwnVs1vsgBvOoXouthNlRtF1Kd5hkAWKOU7o9hAXvnj
/DYRUAgIUrgk9pwMS1ea1hxYULY3kesUMdkOVAVxauHL/blNfLQmw8ElryWEf+gI
3ASKXCGjslblBjLvehSRnVxRi9INFjyeRp4A2iOG+gkyaZt1Z0hDAMVRWsx5jwYr
gWxGkfbQ9Xab9V6QT11hJc5wsgd+2syumA9LRibzck9uEQx0fRr4cJ1I2LTVfOdo
gLpO+YbxWocTS3kzPBG40XtO1RfkZ3loNoaE9FDJPkKxXLpqU5LV7tl9H9Z67I+H
rWKZRrIGsuSjesEhCHRIV0qshhqW3SFWiwSZ+8/Gp4q+GzcNVxf9P0DuNj4G6aDl
c+l+tv46Q7bZx3kOWYBsHG6+Kyrdx9GhVBfFGONAOiNIr1jdLi4eGAX5kWyESk7n
ibR4llCtZ22fbYC2nNgTkneCpTewrG3Z9rjQgRUUXq5xueFxpkKXhyrdZwl/INSd
U+PvIZPZ+k3OlBHT8Xgp7vxvGvHToBNtQhvjcQldRwLXyIE8zufb/by6Vi+NN5qN
+Eb6duchlt6yHaxjjjJdw/eA7+pe0+qhUlJK0mpoBwybf0Oo1Jb80Jfdv9d/pWjg
wschXIByJNY1ypVRvLvYOwyzCvs8HQtClqdEp8V+E13gqgAKEYjMZ3kAqgXQ5wHF
/u3ojclm2BevSn6xyt3Vb87W5Uhi8HoAaqAtkSkWaY2AOvgv64W1K9RDd3Fildoo
6rrx2ZkFD+ePsCQR+nGTvoiFn+xnU1NtoVwdXmIr26spmh+u76JbjfC6307qa4JE
dejGVcxrIqb45BfZU3FJadrP2pN6qzs7+wetoXv01cdiFepC/rzkC0jqkoRFRBXV
C4hAT23SX3S9S0YlELmUnFwyHKTY4/sArt/KF378/KwUMmsCwNMFijZbaU9aLpry
KOpQPDTC7Zyfsc2KJvjneW8xDPbLvEDs9XQGiQ+SI8e+SpGje0RnvllbQdCRa6U4
zGxqJHuJEhnjTw1xmUk1jrhjQ3UEzqGh6IOI+3E4CqOKmiM17DP5ko3zwJ6w4NhT
AeOtqn+0WtcuPfB+BcMAbRZwDaIxd8MDzr2cAwNg3hNgkI5l6/q9eaQorqkcLXWc
5IGxGHNBM2Mi/12QXmD8OgP8IgnCDx/kf8zpWbqu7dVroYVLOHrPKVo38eWlMK7E
qZMI0Q476VbguHFHM9qrEajn8OwIlq010RP+1EfoPFuzbpERrwt8usP3ArnldNvL
f2kzsHQA/Svy5U+VxiOdPfT+xfS4C9smZ4Cvt42APINhKAW6UbU30tOwlP2d5ZTJ
MpdWpOlSOjNhRzBN0Xa1xMw6UBpnFCDVTa8JTnMbWOwQoWSecu//K5A0rw6zPNrj
o3HRfD6sVreP55GMTFFcAtZtztEV9OZS6VkYDmu5tJgTCeJWMBMzv4aSNTQtvlHt
YsVfE9vW1UivzdZnrzaFpDmBpivP/j8WGyJ4Zu+MNl6tIKtSUF8P+pg9nHQ4/aCE
C3raZ4Dp/iXlUCwCmV+UxlZPVjibNvjcoMFHq4Z8SUJ0RC1dRKmu01f5W8REgCMl
qBg0nyrMIJFUpfpSx+znV9ax/RtuWbTQNoEh1gLRSLQYyU8YtFKEuDeUiXbuPk+t
26tD6U6yp2TcD0uQWHZ8Neu0dncfvQGX6mlrrdhjv6V3hCX2OqqNStNKFn4MkN+c
7OoOvjixFXnVFfxOJnMZzGooR45HDHe/o963M2V4dWc8aci+UsrTmIefmVPyE7RB
Lss8n4QVHyd3mqmvXpyONaTI3uIp0ap1kAhYPr4yO5BTVdsvQox1SfEyqADLZXzA
NKcaG9dR9WjTcc6QsEe+k5wDRzK5xRcHF9+5L9UrBCnlf65PVVYqSRuE+hHN/TZT
8gHVxcrZGw0l9boSTuXCqsVXtrMjRn89MU0SFq5l4sHJKOyjBDxzSdclJF5Ge7q/
PdlNzPTsmcRsco7uSIlIl7zYVj8blIFcNGpjBXyYukOJ9fGUdH1UccLBkoRVdY1d
caCjGnZtaLfg9thldqDaSz2VFQVqbRYvIs+A1XppIrZ/7SDa0BcK+lJoOK5GGRnx
DhM7rW7/6zHKywTSriDStD+QxBvlgm1E7oowLzsaFBa9GD6WVj3Grq5D7ORcGtMc
FEpqV157ogxBBIdQuBKAaSJwxGarBm9w07X8dtH91sRTl1p1QYQJYvlVBh/feEjt
VubxXT+rXB92SOl2WYiOqWn3M3SwAm8TW+1+pTwTMfaI7bGABHC03Ez5HFWWChdx
iVeztNfAfmeKSa9wcWuMJtDDZIlGRTr2v/yRO/Izg39giBUzM71JPjDOOs9LdN7J
s6vl6FyoI5PDkQFtg2i5hYaqFePfl9g5M0PtbdVqYgAxlMtPMnv6WP78Zi4BtZnZ
uLT31vGC8pFZ6NQEwRX3sGk7jRglRKCGE61arfjFR25HB5DumNuChELKi1NMXdsu
riNiK2j2MNW47tS7H4EvMm9+bzZoeLOPSYt3qDWuQDVs65qExX4hn1dhKtWkmpaq
BZmS4swhbMP6ofAdqn53u80g9mW14IMCIMqFLL59fhj5vgftAtegB2yxPuao01cS
J/UE9u+LgrcSXBSJZVSyJP4TldCDX2dMhFWXtolPE5WcI32WLJFtTO4GSCHEc0iN
V9yCqrc18Bej+Yj+zCtkoTW5pHeyGrDY7TEmkHt54Q3NVOCOfld6JmwOQ6AWfIC4
YKzdmR0TyuuqxSGUiP7L8RyFXsnE3qTsM+75jGQXrkeQfkaPz9qXrFI30a35Djn1
X8CNDC1JstiUP5WUZIGrDQlnheWolKdo1/xLYamqlGBSFi4rIIM9sDz4ST+VYknW
szlSKQL0/hXqVq0aVnqJyq6MlTp2bneKGGSyKbrM1hhNIdYjHadxH4s16n8FEoXD
SrMh5137ImiaK9atkLXsIScIWBpGn7jmIuyhJVdDrPSjHu2zIO5JlcIsaY86ITOt
GupFZU/BMt0aEsQFpjiZVhtp7kfTQ/GjbzmJXU7M6l3g1340s5F6IeEsupOc8MCT
atiERTuw89h4DVCGOkJwAks6H4Ld8nsKgDOWOt9ybgm4oGWaPtvsWOy0puvFL3tm
LTfrK+GHmKCXYokhNcfsQkq2DpLZGV11Kg8e6otewtMAgKffA/TDwdKhgRKoY2/0
PbkH6VhTgAQXjQVPWY4ZFY2QFus8+ivN5mlVb1kGvBt7Iw6KS4w5JkfUwdn/xrnm
LDZAiGOUjpf3P5lgWGrPgDAHC/Kqj30IAZ6746rLix/jM4crgp7uTks6jee/Kg16
qyp7qrPLWmh+4q2QNKfEJGeCAkWYYtSAI2FSZfw++nCd/6go9ZiveD7oeY3XwosV
F84VaYRWm8Gizd0ruV7Qtt4ZARw3+4Z+6fjxjpLryXdaDQPMVtrnApW3n9sZp4OA
gxjvIRJa49hXZtJHejIPrgautSqv0nSUEl/oM3HOJlmYztw6zCsB9QTyI4Ab24Uy
qYu9jGj/Q5s9lqSk/JXqbgKGnyaqoQFEisum8x7M7O5VSLl8SJzvK3zvC1DQvbaY
B8rktElFPxDakhc4GcnoRNyeoQKGK6eMRV1M13pYALwQX70Vt3fjPyHSAoNyh8NQ
ZiaZF8Fg+A6590mu4HXhrk8B8Al2jL1q+5v8SwfVEmRPeaeyhcN0/k+CRgkS09/l
RZ6o9TPsiITf2rIqxRXOKzjJ7PmTCgyZZt7vC5TwHdPT7B/D+78z3DEUFqiL+7jt
iVoW28ij5HWKYzH5+ZrAtwWv2yH/aMJyRBY/Uz9sa6T9qVx+559UTQTLOYONSsif
kuKk97PzAW0n/TrXyMle44glD3EjYMaW4n8D4Efpp0YAeDCRc4v0w67rPRhjMFHI
XAAS6NIWr80lFRfq+alHkqEb7Y0LYhatL+GdN+d6ZUxwgTL8C0jBYpVML4CwXwFZ
W/HOFVe+jmrOQnLd4V4mRh1XVlsy2ISlqAWpDruD+24WksYfjMjHpKL9GKhmw8bA
wUjmpcPxTjeb4SV0YK1DsQWYWrMOUoqidgIJjO5c7OlWgIozEg1mA7HSCYO8534n
Zv4jcmoHf4KtlO8uantH2PSJRuriXHvNvyNajY6J0LBiYXs3RUmJlLC9dUIoVvh8
6DmVqoPsMy5DgJz4A4Wbrzy6/z901rVLL8FnDHGlnyH2kX/wbv+eBnZRYBvCQ24n
o4+0M5BRDuEoAYkfbnPO9pLah/5yBkqvwj8UlCSk+7E2184An4ZzyLTmfCU+ET0y
+pv/oTjhJbte7FDRgE2/BHzavcMlh/GoQnOUc094/A0pkEqylz3buO8Y/ctdrJgb
E7vGBFZjj51K4vmJ/jIISKpt6fQcS0j6wV122XwZLCVqeDd5+VG0NZ/N5zkLO3cp
KVkj6LzRHLXZ36keey3iSvcFd4O7OesIz+/wSgZm125eoIEhK67F/sAWAS4Ufuic
CChJip4mdgxQ0JvNqfpIL89EyGmhNb1jmo3leqklz265M35xbp80qtHEKg1ohYeN
9+JM/Ponj4suP+/qbrLE914RML1Iy5SLVlnXoa3Q7F/Aqvr97U9wGcBg1bRQcFbs
ch6Q3jJIfwdpkhmT5tRERqupHbfZ8fGQKPAVuEFByLpRmDtxUJoQXEO5YXaqQKg/
tYjsFPxT1FsooMFAiGyMnvF2832xF6e/i736aZTIOYTdOiSR3gkeWbhxqJWbg3C/
2CNw2ALRfOIGdnzwb6bXstYtaaTdVprTGb1c8834zZmT8wFdGInW7ZSSL1eWAM8n
RJWw8TODaRi3V1wfobJvKjoPEjojFvQCEnPuNgWTyd6roh4JZo3pnfsfHA4uAwb6
ggymF5N46ZUR4xvjiWxi9FROeGdp5hSNC4DUZr4UGmVN7dJMYJqbuti8WUFjgXBH
mWmSgFBjc9kjceeUuPb9R64kqLYlAeD0kd7CCn4la752feYw9QHaR4M+hNIj5wnX
gFqXozlCmiaDGagxVlLlxQDkD/0n7MoFdbMqGz6pjCKq/k9mLYd3isGZJTtB5j/o
guEasdz2TE2Q5W5oX0h5ViDWy9yut4pKihVHcBlDxEExBw+Z/OWI1psWYtKTDH8x
sDZIvxpsUhlC8SqfcZDdb+PbqQ7yLfK92UrzULTCf7kBTq9olWif2E0vRzQkRBbw
TdxGhqol8WaUPgjtq7lRdNMt2OQCBMAshAiRMkMeTZnjlkOp30dCFHq0FmyXuyoO
GrFRVPhySMVXaHbfL0x1UbUN8sRqAYkbDVaTM1eqgKfZ4VkN7rQJBh0ZPUzER4C2
aIHezSFb4NEwAdSfNBIEhOmKqOU6YyQUqgQeq9MSPTg7Q0B7ki49T3DWMXR2tArX
pp4bPgV6jKpLBrwYKySnC6zV6EyiShxA6gadv14zeXpeQoVSzpBtxqI45RR2e/gC
eXBvE6VxJ8n8r3BNt8TJ0nvqTdm28/1ROVGXHBPHnr52VlfnESAIqJSzwYnOfykt
WnNc0rSBcL7PZMiWjjzVI58l64ix7f8OGmhgZNpCmLaO/TlCPBb5LaGVUUm0pLFo
ljdEFKfHF53Rqs3/j8R986pht+U6W+081oQjT6YJYvE/fUZWVkjkq//DgxRzeIt6
lIg/7HJVZR/Ya4OqexpwIHlJQIZ3bklLxPwcbmFuMxopsPwDTLSF9UpynsJTCNWC
X2JCtw/Z5j/wgbs21sX2ji72qB6hFp0q/hInogFz3YWyktq3XhEo3pWYDHX0Fgog
7BXWUkZ5toGfHPm7/ehggRo43+AlKV8HKC/+EGOyLnINzb1DVMZOYDujBJbXe8KZ
HThzSoRKWOFYWMqrq8ABgeBlQHvCmvAUnelA6dwY70jl1Pvj/+ePdBGRLXKbVBpt
xvyTq6cU+n/YOZxoGwC2/thwL++9iaE1hjcv9dNGs46OFctoS4tRQoUPs2kQj7Ly
11FV4UkONwIUFp5+xekyMNDFonCEhSjQV7KQgB4U002HfIrC3woTg0iTCfU54g89
D5bnMnH4Xi6ifbq9wA6Kw6GFd2KwEi+i7uW6Hd2MOikm8YNAZj0WMNVuOCTj1UR8
+Ny4E/hT1QG0lXGOayaL6qWjjQMK2n5TnUdgNrGIVqvUT13oy1XeF7K4415w8gyU
m5qLHy6O7NE/eHFn2XX8vjgz+kvt9F1cZ2hj9X60BLxfLXe4IGilAEiWZ3DMu5lw
/pLPp2jwvr6xODdV6ccFKxzxFfj/kmxXQIpbyMrhqEvpjDi0UXnHnNoDOzbEkROw
9/267I41NF63uP1RlyVx7Y1ap+GcfJ3RgPK/9SvACZQ5LXFYzERYes5fnz99Z6xd
UK8hRpivdqTu/Bds8RjFVUBmtWUVZRe04hXTnZZOao0GxhVxEpKDzx07izFrHU/q
b/Mcqy8vrcudJPgZjn0thWJuUUwl2w42UACBhNhslz8Sgb6hVpVFeNl3pzqXw0yr
ElrcIL7Hlq0uq6X/1h/rwcdc52fNoUNcS9D2ysjA/+U0vYgQdsbINpRzQYJrzAKe
0KKuxl/GsGXybZ491OfWQzE8qAHbxVcgMbCUD0JPNQt9GE8o2gpMC81h0gxQQnpl
cE70vO/68vuEXlRGXO2DKfN/DRhHcZdmG8deNoAvdR7UDhR5jGkAPPMi39gu4arH
2hFtg7W2bAVI+PUOKOb9ODAtR6N9TI8clRz/RqVDEBIsJOZIchVwuRrsKw5Ttvjv
TBwEynKLd5cXBLOMP8WZBMMt3fE38PHh2HXjjXO2blxcTQ0QpYi5T7HvO0MZpOV7
dhTEBm5KXvJXszH1j8aTuL1d3SvziC6mj6K4Wy0+8fNqiWwV4aTDWiP5uLX//pzP
azIUTEbFQpIqT33IZJdKdelrtre/jmeOSRxotpN4fyxbIunjyJYjEsXZtHqaspzA
MhpjO2iQdQsFSz0E4KBypECpT/9QSo+MMWim9UGKkOosQWHkbgOj37yHt6PseYwy
vilvM5MPewRYSwIbF4DCvLJVI71pMc/WIEwqXj4fOsn6U+skxsH65bvbwGAhdKjk
cmd21LVo9ewjaxe7+32sbfCRGmC1r8+Xk23jwIBHS8/+2eOQLk+jVBE7zXrH16VE
E+kjPj0WCdoYz6ThoGXB7CQhbLNqvW1YMCy0QCqrqddpe6+9eHInN2motNWL0Cli
mbV3vlfyfP9R62sd6wVTRZjiZsYbo9vyDCvgWmfsQHBdkojFElIxG3per84ZsCrj
RkUA4/IxKZu6fcglO7MRfdTbTU10in2w8LOXiCRZ5vInRCM64pd/6cyQjjjF6b4E
h/UnLZB7bqILU7D5jgN7qc8lxgTbQmw4BZwF5ckOrbKa3lL8OtNJvh9SwE2AvfA+
X8pURnPFkksYhX2/B5R7z7/1cS+mEqyKU/yRgqboI5wNlLsTGSv7NgggwYk2O4oP
owqmocBWSmb5Z+ue1dKYcbMj6HdxiSul4DI51y6oTTufVgAqDbABJtJV/GmYAC8H
nlSc2hkk0Gh8u8wws+EXLFGfkB2gji12/tJgLxU8inkTwaTO5xv07Ze0PlA/M4YO
a4rKyg+SXS91hD6WUnl0SRa9eXKY06lHn9TwiczC7Dwf7uurZ4bz4BuhLPLOWX4J
BAf21cYGeSUy2kjLG9wd/YI7wxOadavy1qeq4A4cs1GAwXwfpYA80z0dmgAcvw+7
1v/MyY5YSspmUVec1GuGGMwzXeK7HYtHxjAL2srGH40sJlwDG81ieP1euuBxQoel
tfyUYdTECWDiR/JT1sAm1j6OJIkosEjgVtYvC9AEMKTaoqXDO+b7T5yS+NqbI/x4
IvijRypQHANNgfYjiI7OIe8oGH0nrw/mdqC7yGzEutULiBgeBgddi7WKsSxkgKwa
V3hOpChEgvvUdtrqqlt0paqLaSw/YwK9Bf6Nv0V2ZjcuJEqPOh6eL9yNmPWY2T0g
OgAu5GhMSn5L83itWsGvr6Zcsp1UXgiF9/pzdx1VhBKe0arjD6c9jjiZu0an/laX
MfhLEhjbC+ZQWjQKSXeOwDsJpSh8ZHbfyCPTHgnZGzbpddmwJjH4NmNfZI5aX4BL
DXrftEi7uNN2G9S/lomnZKX2VkEwqmSmWkVnwXm19XBd08AmIDGKuZ0d0Bi133AE
rTxcY9NEIGHAwT8L+BfiQ3e8zDh3Rw22YUrLVknIu6fqvNE48lojtm0Yc95XgHWd
Fx3VL7LrTF0vXeIFfx0/BjQ6b5eEbYo1Zby6+4HdNayihyOQz/wR76GXAtrZVg8f
PLibX61G32uFvkpKkicHvx1QsR5LE+/J+iv+MKIQg1e6aEujWLH7kHVK4Y4rYw1e
fYjiPvBHgYJmdIItu+rt7CuZOUJApknbQjZQXccE6xxLZ77w08optjDWOm25iiLh
KQ7NG18/I0EdLsnvEtXhZXTdurVU9WfK9oJuf0PP7mq/yLSsgLoTi/xWxu28E0XP
3+V76BTddV434j9gLaJTMogHrJfB/ZgPkUGVm3qWzIs92vqn/ERK5KSx8rJUOJWq
rPBFHZylZ++kCzs0SX1eKEaGLGpu3i/tMotCm8waAmiD9uLdeNpDJyi9SLBlDIQn
sxrQPtRo9cwFV5upgMLuZD+SPWfUe0cmMqLLSeIjBb+xsgr5YGWhRRZZtVfAz4vC
AFG5nAdCR3074bHI0OdD3/G5YnTFpZBBYQsDzHFsiFEbHXBTfusPozqBcfqbVbM8
6suj1BolIDf6vYoJnOv0mitdpZ+BQv0sewVYynM/RAfn5KoKyi2LIfqh087PnRZd
gca+e8IeUHVt1TJsK3cuio97+F5zhmUKkCczlsiRr7ldOnQUBGnjp1L1hh/rzV+Z
YfyDcO1NzVydiedLS+i6JKzY1CWaVHE6bTK04uT6mXD4Vahs2ezVxxdOt6T9Gg7L
liMlVxc7dZ8PuK4x6eAajnp4EnoHsZ6xwJVSO3oEgsjsc+TC9IiHBkEEroYRmKIt
/u+piWV4AznmGA2TtaB0c2bpm7biiKFLat2eOv3b1t12zuIxkmccKIGPVUV94Icg
W5YdC+JCpDWJNumxCPb/9taaSYZvgX6wcZPpPQp0RnwqG95eW1tR7kGgwoYF4yWJ
Njj/+7ewsyKFJxptlKw7gudOiBjISGEfgkT7DajEgykqPR4aq0WYidXcvyFjU7u7
OG3fLPv56PyTgt9h+D6oUPaqfQCjR1C4eN9x2uFJZqUmnRCI2OHVkg3Pyk8JtSI+
gwh1ZNTRJzOjZljKINzHFZ6XDFGuQJy2BmDZrmTyeNknwMU20+9bsbrNlllKC2iE
+kyAfYyFeJpGKRdhKz7m7zHph/7t5TiHybntDp/eLrVJIyGIdAb7AGgur+YfIt6K
0WLNjaWz0wRNsCAnOjf1bl4ZIBcBfun+AeZywKoD4whqeBA4X6Jwl8Ii4cP26H5B
JqXaSVN0cXO9hNmPMwWDSBS+M0LsJM4TTyiRnCYYt2uk7SI3HgipLZ9KSqrcoo3H
OYUOvsatQERCtVIy/M+TR75Vs59Z3uMS8ZB7vEEgFg8SrhOD3wXZ+D7ClBFrizro
lJMEJEK4GKY9M9wpVi1G9X9R5FBVPgC6wGeFtNCZyRSYyUzyFJdf8eVyV6zBXeKO
pOFqGSUHkiOJZfe4EjxylKtUT/JvfQDZoKi5d9ilojNWykDdmN38/KH+7BP4Pz9W
rRp8zLhAZQNNJbDTb+o0Gqn/+/AzcdMpVdOB2AR86Bq5fIFmu9d993ZnVc5aMtIP
dz5hCpjy/Z2EJeCqEWsDkn4xEAPiKS2ci4B2azgMCbyKIxKeN6I7/gaSPkz2C/sN
F319kLby03p5+fCYRW2tTpsYWKlQLRAOCqLT024+xH7Mrb/F5p0anVIidG1kkc/d
E7ndHbO0C5vtpinSGwow+gffUUfCQ7krSEzcBYNmS9lBBzVcLpCM+naBttPafnWM
kgqUuadjXLE9GCBpORqolSOl4+q2MVJQCnvwmirQGIxJ7MeXLFu73W+cnKorLjJ4
JdSKSRPyQ7p8mf1FXpYyaO3lro6+qipVE18UzozeewRL7nz6YOv1heSai4WiECqg
7hugNEaEbT9/RIhXIAFmc524ZY5KXfuvY3bO1HIfCVjSDJidfMlTc7+CLLEVPdPa
Kl9uEQbjwOeTC0JHqy/r8GAgmkWhtXLPeocPsri1zzzAthceHCKdK1ZLuwGhyor6
2uRs7MpGgGx+in6HUu+ASrn1B9lLFoXwA1pbTFE/DvssRANtU5v8AY9Emgw3IfW4
AGsl0EFqMpCt+iaGibLpfo5Ts3btULMtbMcv1RZfH12PuaL2kNkiXDGyV9FrdkOW
qrAn/koZuk9BYHf6ABFJeLoA9A6zEJGLWywB9WW5Q9+7m6bUm+dnWv3SOhwk3L42
cv3dP5H59B8TfMRCTi2+aphfxF8JlxwHqoT2zJ0qBw3QU7/rAGKywH14DJwkYnt/
96duAJHBbiugoEev71jt1wmlH8vanYev1BhhcbrRgg45eo7WNuzyuoK8AXAWXBvS
eE1zGdz3242dQdnK2jWQmg3w9WRId6dNYpYts3FKLRHTB6hOISZ/8LLql5iFMJf8
/5PYzYGFwu2FD0oEDeB7A1ygyUM2cs4NLE7JsQ/VDVPS8DacgorwNy6qwJ8QTvjY
gfaQSdkiZsLVF4h665c4gpbTK4Ef5zOg9uNs0SN/sIVuJA1FUtSdq08ghASLm/8c
SXeH2SGjhScVGX25n67Ceq0UN4TdOXAItlH1g0SQ+baqstoTWFWLfoHDB0SN8298
Nkgi8zqIvbijrJslxbF6tLFUW4VeGI5Phwq3JEvONlko+kojQ2TJQneUyc5Bt0Dn
LR4TZkG1oEljFMcvDaEG4rVP43tRwX4Tr5aXhOt7zHtDQ3CJeV2ZQ6kXP8SZ1sx0
X0qgV8eZyzp3/Ca58jZ6OTiUsGMFHCIceqeHK8sPwOtRqPC8lgoV2TnGwGhEgPXl
+2FpHTgjr/AJenSTS7RTrAugbNpvqymyylxsdUHVoRCNYfb0fV5CTx58sJWJr0fN
IoiBw0ao/tttsURNFPTq58TSx69szRr1WVi053PDoXt6hLyI4smrI3/boUswAzu8
LYf5UmRlsp/VOvwbIC4qELonS8nqHSCWRzVP5SEH4h3rY5OvWx9LxH0quqCDnfK/
r1+SHrJ/ChahjuX268HElYrbe9eT+/2bU/wELCRHP4tyiPTqtgICHq9Ypm3QXuVV
3qaDOGosmdvQr0gCENK/eS/MjgZHORXcrnpW3/XAuixtIlL4WiGQIOMoQbuGzmk/
LtA/gwEA1ppBU1/isNdq/+FEtEdxqy/5u0aSJGlRZ2/OwVxH7iu80GNcjmDGS5kJ
YjvOkTiY5wR1DQYscfwkBbWV6keVbNgAWaPhKfHEQWUZDcTovUMAjnbDsS1yDceU
s/7NhSgqaTShBJLm4Fc9NIpUiPiAVoEXkxZ529xDgw02OHdRhmUym+gFik1qA3rO
J13uL8P0RpSYEWD7ZGvNoUWt/PdIgfYWkcwsIKozb7uxEywXFtyYZcIwUl011DFN
tQu5nFvIbyF0HkFIx8PlxZ1QpSWBH8/Mj69msUBKSMgZhxb2aC0s1hShr0MAJW5/
9zBU/l1e2dZP9ol/mMYeE3dNmDXfkXUCNepcAEbsQwF9vmYffnkjKqMYlaCAH8DY
Hgpe42iJV/MGDN3cf4lt9RC1Krpjf0e8hLYuZFAJtgrwfHQMq6SJsKIgn12QRjpc
qI1UdUiyJScu208I/wVbIJTYle6gXEvMEYMu1Ef8F5AYkQAifwoXJHjpSgrPKD2b
fGZOMxbJqlfe2RrL0Qbc4B0MC9jutpuukZ5QzTXDBDClZb6SW1bSXK3j+ociG/Cy
xzepBNkQw2k2oNaDd359cxLQhUcgSiSVivkxhuuETnGa0WW9XlC8+EzeJ1RYE4nq
H0o8lfOf5HEuRcDncvOsx9pbJ0GrBYgDv+Ac6/NKzD0AlfxEDNjQVS0ZlYS8xTlB
SnClubNVC+vLqp+d2BVa+AUtrORoXarHBt6gma1L56Z+1/dFAQtoC1T/aJUcjr1o
BRVAsjoE1RQttNp6cFUmJuRL+amdK13RE2jscjYLzo3D56GZmeeOJlBSDNodZxgV
hrH/Tb+IjJuVj8oWjW81GaE3wYqs8sj6xHOJfwKiJ5k5PlURMkGo6/b8wQTalSar
1ESd1bOUhuIEMHgfuXtFmzciHxBHpB5p36KKHdpZcVrCiVB4g+yf8A8keUzgy1li
qm9dw8WO7iRnedURlCtPK4KqWqCYD8L+It9MXlWfCwoCIn3ZEdhPo6LveW7TK2po
cLtXdWnUtnkj0puYMsjR0dBek6QWfD9IHPmOCEBrtJG6XH583L0wm7lAPUy9kL7M
+SCiFAnoL+S3pxKvVS7R5d4OEFLnctAbC/zLQ5eMxzEnsyr/leuDTTCGrPIQMCTr
GiquBb120RxsRciK9ru7J6ZCE+kls5OqOzyfmMtQ9+urCuhKObbAda6doAl4N2DY
gbNhJlWzwXvpRZad62LBG7KvAR5dLeS2GAmy+XHbu4AP5wIGRcFMyhkNy8Zcri81
U9LA1Oj8h8BwgOWSTw84BexAVJlYXFts8efujaxOG9lR7uifvgewbsyZe2Mj0tQf
SKCV81USILjYwaUH8S6+ykckmKRJ+8qWjOsnmcWHQT+KlxJ+XyD6ExO06nxuO9Aa
ixuVds0DIEfZBdBkWMYOLtC/afB9+SfptMFNX/Z5whulPILejUYF/xkv9CueFxcl
FjPZQgAIMlrEiJKOLFNRaKobJZShFYeKn2UPMQrm7m/ZP9CfSn29Nwrm/PlWvm0g
YVLfKzS2+m5AlWWzfjClQlGrtYrLH/ECLEtMDnnQe41biJIfKuc0QdppqLK4gWM1
5snkEVAkwgOCuwziUt3e7Fd6X+Fauio0/wz3Z03vBfN3KLfsLbZtItHHLov6yVdq
qq6xlrp869zaMP1DN+KvNCWjJja2/y1rdYNuEuMApxLrNRsNOLxzzMjGnGzmaPhq
Vu+E8DQXfIsvRVFKq5sXqff9aQY7CIVsy1AofT98vUBpznFgeIQxNJYwAU96ReEX
+dfByhiU6vn1IQxLLZK7EOz6VZ/5skrBH4XD56FuwqFA9o4al2t+LZC0XNtNd0xg
QrxFArXvWgh0N9jgErG0A2tQpCumdFXbc4V9ZFrZH0/kPqErjo6KCk9THc7HvREC
NVktkthQIV4aHcrx0Nb1aq+R+fqZYJ6K9sgxsCzdUNJR8xo+dMVLd3viMGZbuxsX
0reuTVhwe3LBscMnTf3AxRH5Tm+DGxVmYETt17ZQLV1G2bVxIvTH5ookREXl4jdv
xIw4KKNuJ9zuLbTBQUiVm60lFo8d28kK0lI4GBxaTJsgGB+2TvU5ilvbH5o3OzE/
NuMC2qzFlsPT1yq/uQWC/kCSgz04u/YR7iZs5nkBQOx3dYXMDoBnJzvxBrTU8Xzf
5Fb4HZvRRJd2LkqX4Le+Wi/pHy3C5VUCETGH5zND6CXQGaTdTLeKms3zl+OGigit
PWIRPLiXZ7Uzjr9NckOTR8YoMWye1vdV0OEJf6znkIdok5WxgXBStBFE8nbLO45i
jEQnraNsAAttTTZtRMXmIlCGVYEt8jZCFQbnPINh/jrHNYjDikgy+LTw6tUAXQRA
LCzOh56zmPj1GYcYPujcIRD9Eyl+Dn52z3FWKTyMe+/E/ixvrb28lUwPIZc5uULe
eGqoCMMJ6QcaPeDMD8Ca/Ti3U/R30xx3Jnzv5hu6Sb6jzztX4nvFqDAR3EhF9eJe
dR3xiDOxMBenr1AP8iZ9+gnSYdz3yi4KLT1b1KXndEQE6omtVyRB9DBnOdSofJ9U
jLdHkF58JzZyqgVY8l2TNVcBVdoOt8naqVnMGrbl46vZAqhk+wHHqmMkuyPGFxKk
g6fLlXBjmsY/8ckqT2PihHLbxgDFB2fGMMPMdDUrJdkmQqAZmVqhAZh60bJ+2zf/
gLrVcodz94argO7pvcqcbypwoTPKYBDBeqiA63K2FCCo6UitSl/9IhzHWcf/Gs8h
Xu8zefBIbLnlM8C9gxIK2QuOomZ+VU8kJiBc0E1164SASaR6/umw9jHcsKjoQesC
Rj0bN1UyBf4J6iiQXKFGTqSe9pSB5Wqb47OksYGILLsHgvNV75bKyBB6gKjfG5bB
F0IymGKcdPfa47AWRCRwySxibtp0/nMe8j38Y9Ql7BTXHeiFHRhkFx3my5aaU+6o
jVkB0USFl2r7lKGzcCZ8VaPXjLjB8ZgUdL8iWntIfbgNKiFiZPTm2f89j+7UeQDL
cnQv1u+dtE2ph9W/aQh5HrKgKtPznfYYSAydqXEOpZm4pM7+MO+EEPsUcqjJz7di
RLJVEkVPUjjlQln1ChfSGapYYy+P8Dfy7ET9BFp8nmQ/943teox2uCF54XKBAyEW
PCNv7l9Dd7HhaApwk4za5FQNQriuPrWd4YIv96UMS6LqR3Se9LXn9abDRJOIKmhZ
8K85DlzWLQrVnoEBi/WynLHDSBVkyM+WIdiJHtWJVHJSammCwGZ3Q9rLXNVmI3ks
1G6Xv5N3R84iDkyNALHxIirCK8HSDgDoVaHQ3p9NK8FhGDww2rx2r3yQf7msFTDD
4hxt9kdnwKCfay3X5fRx0qgcvFJqeFJrBZr6hocPS/VCnxcbDAwfol2fVYEigd/4
1Bh+xWAVUS8xei2MiIrASv1zBHqEPOtFtBB5uCqxb6ATPnjvtJNgrn+tVduwOaV6
AngO4bviAzQdqo5vZyIZ9KVDNic/8BdqzbAHInbRx2botoq3hIF6mgBXYk2bdSMf
/cl82k3zfzIHiDNWsL7mhRWERbT//iFPhvvzu/QG99PdKBf0xdNWiq6hsZiRD11R
jieLcbaFjX9TbcrpPTN2WYdX/gTWxNsvNJo1TKGjzTKmIoRospeYpmOp2wdC7Eqa
TZ80/KT0QW/FMVqmSj0RoyLUuQY5+6NO9VBUK8+tzoa6IFQloREqAUK33u+pPASK
uxXCf8FbJViF61C9/lhnLWa5KTTGJyOukTVZ98Xt93xOn8m8kxd9/nn7ocd4l7fi
WwLDnW1seTrFoh9nEcgYWCvKVT7HQY5A2G4FQzmlUyUHBXltGnZlThQJBioBhLxv
6vvl3S6+2P1HUxohX/MudIsCjoFLG84JR0xM2AeIejMKDcFEU1P4HAUl1sRGBgW3
24FrcWdQ5Q8TYFVURNwWBhONYyqQUstAj0Vmx1T6xPX7EBh3KwoHarY4F+4ovy5m
qUkNsnqLXtdxvl2IOphmDJynAwnN/izfnQZTygyGmjehyz7JtwMqOE/PnF/7q+sP
O2+wZ9BHGPJPOot5dgdng2hNnLjTETLCn8C8qm5FCmtW5aUpUmpcwjPV4pBQhWO8
XTzdVaGSFfBTeSkkWuDozxyGuoljUmughMCYLp8se5icAsEhM5qDDSnURFvgWBby
cow6nNaW6GyUBuDH4DJcGvCRpJPu2/H9foScjkGaChv28Uucs+qM+QFSbOqdv0D4
e7R0vo1LEvh/mEr5i1PGP1/+D6HOVbSR3c/2Oqp1KhSlL7Esba0DrzPiqQbsQO7D
CIJ98+yxRPOPanRWVZ1R1RlibbZdOd5S2ekjZgVQ7UaWEmjz8vQDm7cCtR2ZMH0X
RJK371LsR3oeJOhz9po0Kweg4t6mPZ8ldBFk/6IkXFIsLqt5zwDcL4yS1AHbJJ2f
TcM5qTvLNEHiz1shmTI6SRGMM/+tYHBR8DNffyZJYLy9zaWPUcbCYdWp+M3yngzv
Hxv9Odz9iEkHx1Mm4cXWvaBJCzI+WIzAKi8PNfd9Q7mt6WdzSu8I59ZMCiaNyQul
dqH78ervt968yhuzTtHqOS8c9EXOPYPBurLtPd0X5DFY9Tbv4kroqgnE+RdSEUrC
6pWS/DsjSRR7cSnBuc6DPpZrLJ3N0m/s0K0GdjN8cVkjrfKX7Pb6kTGvHJzVmUbS
/Wppg3D2eoMHYPCvI0Y0E+w29ttvpQ+CcMVoHCh2OGOrjzweEPXzouYdbpD6zRZw
INNqshFgMbT1GfrAB6lJouvFG2D6aObaiIDy7uzRZ6OVsIUP3hT+1B9j7LRKDPqu
CMrS3eEeQ/9Oe9T4CGKOAhT40LzKZOtNopxOnN8xFyz2JJVeCjFcuk0aSiJ48eil
wP4cOkG1OhMonh87KVQXyoPfa/NIyKhWdYC98YBqZJpNMcA3i9/U8BmSECV55yBK
ZWpZaryABcltsN4RLaRKORftrUI/AR3uKX2jOIOTYW0qsts7J+ZhMsAas0c3akjU
+P4MSBKV+WxboAbZqJbsg+46cIdPAydD2rZTt+Kl7v5Ixf5hkvwk8MXTdTTrPt4i
p7Ay0cTqsuoaM+2d1iHMCWo51u1u5KW8qDTrDcr8Eh7nihrlAW5ewSD0h8NEAbo3
mZicKzSbxBCQjpErvKk0rpCNjMy7AXIuAps9xIeCgAhzxszF0+Z2Lc3GYC1+EmuN
soBM2eRATa8+lslqxY3VzR9JVMjgi4fNuNHjz9LXe9yDU49tqNcTM4m4eseLDvMU
rUbmOdlXsUrzat8NAJYerq+6JaUFnVBq920OsULvWoUiFzRORJwZC2RID3OaWKmM
cwVk/SWsszYONwppo8cD3YFq7q4W5q23WhkEwd2bfAayXJMoDg9tQs94cGQFQmwJ
kGAvX870TIm6wYLi6toBag71EHF/hQ0wUHmFAzOFHH8N+mb95n8RUIPrcRKSF6CS
jIUeWvzNf04ATf0Am/VKey11ho92VMeZdccBDQjpQ7ghqv0E133n6KoIRHEtU18z
Ki+yGU3MTiFCUmSN/1kF6O3xIRSTU+z/BCb879IlNIbs0svhai8Em3QXFd0dwJwr
2GhUocWTIulaub2l+SoCr+LjUSRdNz0k5S5OB3ZTZmvR5bnudBRKx8OqTLl4SAK/
fPGkskQ7yFVLniwJFLHKUfroTIT71l7L9rIznk2V8jcSDShpdj3tvV8Lb0J8wLS9
7AUjIEzYYhXXIblOFiiBOaAjDN/sKwCYLx90zbDONZfohJ+u08dUkm/jCpJkdgcA
T9J6t/GO4MIhTkn7JrfM/OwU0763TdUGwGVYaczXIcn994Bu2WGyAN2gpQls2n3L
GZW8pMsLnzMsoqLYc0eh0agH1vsuDE2n9PQ7e7lCXksZqgz3/39Ax6pGAU5cPhks
XDXQILh3lt7bvoOK/X9Rh+DDlbIb1GQsqln9Zacn167g5tOL4d3IZQQo3A4uUCGU
uqKw49Ywa8+ZGkLL1zmIr1v4VVsWRXjyVFZ5E7ypbC4isXedSZcWyQe3Z85mV0iN
jlKdctQ0jn4zVUPugAJbm9yh5psCy88buLGDrS+7ynPh/FrjUh6HrCYFWdh/VFor
dJziQ1xt+DL43NZ7UEMN+oCUsC72bHzurPjXIJ6afQ58GQdEVAKbgRwThHvHClXB
KiGIEZOqB1gvzKeYhJ6PTa0hrFdZNZ2cvEs7odvToYb6PHKeQDMAxQeqEsFtb3ty
A7ALn9pDuPZoROVv7lysfQhCjs4+tMQedjJjZu9TQfu3dsNrzZ9MhUF31iYJXJa7
5LxJDIS9PJcKhYh11XUC7Y6QiXhMCCOVLL5ObkZSvksm+UnQoRU3zYxeE4evcGHJ
Wmq41dIunt4gpv3UpWlSD11ASV8fJ9Q0P0u+5ky6TBVSRJUs+rVhrRnHLY6INghy
oM7RTxTq/IeX4dc0VUqllkRSGmtjSjVwBsKPxy61aES5kSYAvApOfdbLnOtKAu9v
oTJZK1I5vH1i6Iy3vyqHjI/StEx8zMxdz3ZKw6WlNJtCkEnNzXW+5WbW+DbgNWXt
QGtlHSriStf5RgKWdz0RIGraE5rG31Qo/sKZjH3k8T53fw856p5FaYIXmTpVzFSF
PiA22xeU7Kb4bd1cZ1T8hcRiJAuSp+1RRTLLybSK6RUsaz9PbNOhA6tPmdzlJ5uI
7TL5grQtvdbuAuEZeYnIgEoaMg5MIWIbm7Ceadjiax0wdflnbxD7Nk2GckNKtk40
e/Flk1CYmwlAAyOWcKIwPhnqKQi5ZyVf69G75QMPR8zVhASr8+PHFM7uyCt/Egey
qd4jjfpE9o6DBsdrUmp4jdJMMU3gGnZk8rsL3SyEuKAzkszVSq6N2M5FHT0xRULs
CvMIeIcZykXxlAqKDUmci39xSBxxrs2kk2er/SklCmTrJmSp2AZAhz8d33MUFyME
Ik6zb0BTUY3yasFh6wobGuJW9DCUpHkq/8HPqL4VJJGOSuCwwIFw5ainleDpsPkS
DW3tFeggPKzE4FCKBH+ny4B+5H5EyYuT0/R3qdFJEwOQlZEbEuBaSx/uxtO40JmD
7NCvytH+QzVHAEGP8ugRuHMYEZ9M7hbKpujOM+6VgBh5a+8m0UHOVecRh0uvTl3x
sPHxtwPK+bh9gdMmVSewu3lFXKbFn1q4S/6hM0Yqk2huxKkbR3Dh0MKhmjCmaWcJ
+ZSch30gKaidlri6f2JVpUTvpeT5bsbYqHBdICB7GSPJ2RaQGurCkO241ceEyq0T
ogm6MjovN3j+HMbJ4ox2dC9R0MMRWAGcATfPqVbfDzjt9T/3aPMowqjewh1gc9kQ
p0V9TebPHRopk2G1ghxUdy5wzmLQHlycrv7GGUhz2o1K8LnJR9Dv9bzWFKVIZWm5
KaeMbFhDFqa46KuaZ2e9q5j+acC/wsGjV1rVGe+pcrxrDGdBuWXIY86THWw/22eY
EDOR0xk9tcLf91xDc2jT/cC9eywYuOZi0B31EKob74j/FAVCUTpZikNzd6JP7v+L
vd3Wl/VeLgBx0LzSn6hii1CHQd/P9s3kb6NTpmqLpe13PGeO3DHZU5sgfAauYc5m
wYkh26waIlDNHwvnXQ5wpPfa4ee9TVbS2k6FgHtY3lydJ+vEQ6tnIjzdNmoQ8Ws/
f9QCZNHe0hbSG3qt1tFgx9QGID1EFN4cJCivyX4MnKL+Hc9TvKLHCMwo4/grg0ti
yCnni7ALqbMk3zsXwjrn3/i/hd/RdrQfQP5bTWidVv8OtJa2C5rvVuh6umoXn9B3
EsOKnlyEIUGoWDYqXfcqOXuPMvano+huf7DrMDmFBuFyVwec7XPOQAein7AIs4Bd
TDkUL/JcpwipS/mWmHup41zskt8haIlpVTWJO7mau22IouUYzCVIYxODE32tV4de
75bIIxd7DC7D5cJZNb+xn2TzwEaj/JQmV06eER+SuKrGYQy5TUoRYDha9KprAqDM
oQPkqnK06+Xo48e0Lrud2FjsW5yBUUD5Z23K+Xhf5XdLRnmPBZcpmxfLkQ3dxg/x
olHYi9momxiCNq7rkLHt1EuCrK67yPM+cCKMR/JrItKt7A6ORYYIb2um0npCtCLK
l0OEaQp8HrdA9VxYtCehKyQ0y8T4TWZf5jvLNmRxQHsBaIR+5nSrYml37bheLI45
njgR1lww1axgzw/xahAbNwoViw3sjfi7FbIcqYm09t57V4X7dS6NAnbsYOBgY+Jq
xpb7dqmb45j18RMqj7dZ3DX7rUlzSZjT66aPKHKFW/yzrLx1wHV+nLvhQyYS6Yud
qHHUfALWspnW72PQBX0v9QpjE02V71UtsQs+0lrsS1jCfS6B7viL1xB+NvuM/WAC
Os7HJIGcriXL77dbSj8z4dkeuiPH/WJthHyV+lZU/gqikn9Kh3WY0H2rX4QWASpn
XWpCruh67HdQOlzKgn682/VR8bmjocEp4AqeE16UFCkInorxHgWy7BBzqu4knBCa
wDh/liIC55zuCf1W5regRo3lgIm0KpVOLXWMT2JMqgLThjn99kgNHy7CQ/8GtIY2
20VMIdGH3Ga1d/14OyMzlyEXz6Tf/LQQL/gS+gJ4icy6VRnARe2Jtf4dkoZwjm00
vLj+qCmqkGJglzUdcLnBwc4DoqEXCnB3IrbnHs3nJ2L1341B3jjZYKEnqKHQLmqz
7uuyxjN7Qttbw2kauYnSKc0NkxNHznP9OWCh4GX85lhQXrfZbcRq1Ld0aObIrS66
BfGgXfMwNLbcRVmTqOcxavYW+oqyDUSbCSgHBpEqj1suwE+RG/LUQIsB5AjCqo+k
1zF16S2CpirbEQKgrurAufQFBfz1E8VWPVSolvuugG4oJtA88rkPIEALujZyEDWu
r6BHWUgwzyuCANROCcloP1wBnqaShJlMI9zqaEX1IH2pcCzjsBw2VrXY324P/OFB
zqrA/kdZwWSUO9r5ISRMlXKmAdl7SKFK81I5fWmnQH3V7V7dSADQcMrvT/dLA9nb
sLqw6Ez1p8C1+pdN22iamQzwDtRrnGxjVIbl47+3JdeeFy3KK501lCiZ3WlvkMtY
xzoiDA4+R9IvGwEpSr4iSS+Fz6k7jtN7qHHTnmfS6jlYpqUR3KN2PZ73HYfxhdIt
qKwlkS2oQjhcSsluEqIZRPJaaTCF/GVIWQYBOKGdTiUfolBIDh5v5DoFm4PULrz2
MKOA+l0t9uGp+1EfShV6f42BBu1AnlFcwWBkDdLtnrpUZ0Txgu1jw2B4sGhg7uU0
bapctdDmeJXhYsjTdn64EGc5ZpnQwQtECnUQct/zmSKeNJZxpeyq06VP5jlQCcJf
h1lqGzcEJZSVJ3rKG++22LDHGkM149yxSufDGH+q02CCsPp0NT1kgbXts7huDbMl
ayrAq0pjh3Q6dc73Jou+Jf8azjxZzQBJuqPEB8nLakevJfEKWwtD1nhv3iW+DQ3e
17Bx981fadOtVu1gcrszG6K05Nlk+YEglSY/IofyKj4owzxlWG44EdH0Nj9qDsTd
uy4P3OK7kTznkk/B/koMHCsRk7ejYRbus4lysRPiwRmEMpP+suUZCicv6G+3nliI
Bd4XqLy/tD0ScQ3jvJXuR3xcOsXTDmibqsVyacrUymlOJd+DyM4zIYlYA0cXMWRE
UVWdPWdiZ7fd2sbQt/t5r6veIIJESlty54MwHrq2xFP5hRgcMq7PQP6N9ErhN+xf
xU5Zv9ghU5tKkybs8LgKggE3JFJ2gdYXq+mj2BDmzQDYvpR9FzmPvMtRRp7Q+wUy
NtkZoQqmJq+w8gXOFeRbF3c4KNOElHIMVTAhyBomyVymDQOcUfMvxK6YnaS0d487
EMUl/++I90bguw6bxmEgMX6buVoq2OKynpdvJHeLHYtVzAVmuScUmm6AEm7V3IgN
PSi2mylBiGv3SUXFpHDX7hhLztUvDXfjQvZZ4xoioCP24Kg+DoI7KHyg5WG94CHo
M91nH08zhCzwUVGKFkA1TyryvcWRZVplE/u1Zc37j5LKgjsvFGrpRHdUEYM6ECep
4OgNOhmRwMl+FQARemDDnXhg70r80dhXgGl4k9CuK77lsjvJJ03Kcra5ZXnRhmJK
8IwUd85x1LqVPznnY3SLkZ28I07R+C2I6iICSUbZtUsCXd0gurJ6X5mfAxOlBMzC
S6uotu+0yZdGusA5ajeDubC0wsriklP/Wf+ZTMP327GeFavFZCRRI7hp2o5Y8zuf
fOm0LUlhi5fjY3hk7qmDQyjTL37gYTNQ/nmfti/XZc7I8Sbd9/QbL428+mohRMn7
kzpEXuDsRd8n0Nccc7Sv5gWLYQbYiSmO99D5McxiFKr/tmZOTDM57REH8zHKQXyx
EBSkb4EaGiE3m52GPDrV6zGdMFh8OS/EJSRPmPMNQ16eXl9Lvz5a4AXPzQpHy1H3
mMqdbqEUDZrEETVSVdheP6WEd5q/hgQE0OzmVIyVQRRhvj91xhp86gFEtcODbkmU
hdMVDQgqGoqxME9wkoUZ5VqT94IGMstaa75dUSEFbfrFzQ/T+b41zw/ZbHL+IezZ
AD2DWYULJqPH1RIBEHUfsMksp/yeLDzEBtI9czDiZKrfIf/D69Dl0wjT7ZVru0v/
mPcuv4/fZOL1U056oJAiyZ/6Pr/rWL7B/sIQ4f7np+ZLIHE/XD5tRk0dewc9wpGo
wLMRuFqCBkpMMR28xGYRQPQy58pnXlkHWWSJltZ1x/7KfNa/rkblRkpxz22LPSux
jJ4wtfIyJESHB4PkB+GcZlv56wP2ThmyRgxx5Rx9acT1nBEZD8yHDRYQ9axYwysz
BqmwBvZfOsCmRLWhoixP5aidI1CZKY8IgFjTrBS7lf/T0YnqcGE3RoN4ryTpXPDc
dxJR9I+DPOjf5J6GO/TWLZuB7pQqTxAAT2Mx9rO5poYB2e3ECjypNlR5WZdxCJz/
6mtzAy+enXo3s8JhR55UsTGBsTQXi2fw+U16UvLUBPAFplpwlIx3YsmicO04hMGC
aLlp5x1POi3pe6K4iJRHGMYP/zKD8XeHa7a0qDF0TJeccBM93EAx6XiJOgZUKTAB
tXCmJnSm0kg9oqUMJfe1mhXZuVLVSDbrYrvSXCt+fLNt+PHewmJMPmJHiktoBWsG
L0WFdcPcFv4PVbbXuXFgU0NBcro2dlNiz5qGVAEmcesN9Pgm/rk5K9KaIztARDEy
6/Yd5he/E/QyNE3g71ZAX7qjMZvxx/R1ugVQtrSNVR6K9ExnaEFYpHZhKEmy7qoh
am4NSjWp905HdsptWxNx6J9qSwFu2py174cuhFDuDk0L12mOcNhH9gxuD4mWzNmH
Vb+KQmzO6M/zoVUED0k/drRDBT8Widdtvq5252mpk9mSIxfDqsaZ9VoPKngM8+pl
OG83aMNRnZ2nn0QCtHCAfYFHVXgvYJaH/woDBceuma0ryMJtburwkMsDPpcu9oqo
ipLktBW00J+Tw8yLIPoTf1FEeJKuPLu5NvnXTcZDXnlUhwSDUrDj7cmnOxdEZCuH
JvrxrKTOfygKDgcnuI9VmVdWxrlq5hcgckTaEFXbnypmkL3qQqzYHC5vGAn2HT/l
oJQ2RPdWz8Bui+zeJ1av7eBMDDO18WNMnhGoEHAoMlmWpHh3zGypmD+IpObm3/oR
FxKB5eJwASVbggDsr/6y3bf+4lZEHKNA6f730ymemniES003i7hA4r3QWVRogji2
YokAcpkt38ipWOMeqeJmG3fPgUqzvKeT+P2FDnGDzi63pGYItlnKWwocZP1tj7Gp
aSg1by4E8EFL/ysEqPAb0v/meSC0RuabKClzPlvCTtaZdG57a/bDTp47gOlDuZOU
y4jPvaLc88GcL+vl7JCtx5fCjHiRuMBbdyk+uri9tpouYsTWR2gIaYfUFqnJV9aj
eekv2OnWsIjcpJlkxQvQ0fXhJRdeg7ZqL8rAGfRkh65M9/l76HHvE+fqDMHuUyrM
/2JSDgCnvx2qS8JEnZVcLpmc1OLzY2e76fN9/GR8fFL1AETj1kxJvu+I6m/rI/2F
hsBdSejY5RbQxC3DVK1LoKS4IRDJBgBmuRZLtiMMCM7fHfv1oSK2lseoh6YD/yj4
cmvrz1wQ5ojpNzHyHs8KH2qqYuBCqlg71obpl1jqkQg1gzbTAF72gE13e4agRvAP
B6L/bGa2Aq/NyMXJjv8wOcMn8rFwrfzAW96CzfZTE6UQoN4cmjjmylZs8nwvRuh2
pbYsdwNLkeWH5EL0JL3AkDcz8U1BLPGRFdjdE5gZ5xH/RhHfcLSsuq2GmRYL3mfL
tk9dcMOVLrrOt5Tfae5BrwOfA3KhCwQzoMbZZi8l6Q6Usw03mfrpFtmzcl9Ok12c
baax8Xjab3xFVWqRPU+gFjI04YM8yRWk+BbqL2c3VpnYCQe5BZOdGvtOPW6Z8r6W
C1+5f3dTayXTRGYhb7DSkVDV8WU1crnd6FmgY78uzED6rNLsPm15JZVkOdRaKsSn
ifS5aYLiQCHD1X+4YUC+Gf396zXonapnrmI17QHAV/OaeBY3eB0YZtH2ilbeYDZT
2ni0R2chwh//nuaVNLzUrkk4T6k1xd2g7ha9iWay4uojV9unI7+uB21nbinSjxCH
tIN+Wm2qy0uHhDaPMldbIPtA3JtC8EwfwsfFeUypuBLINdRy0/he1uJp9dhHUF/2
4FIIslvz0Fsn01dVky4whO/TPiErnGHS6UC+RB2a0ttDJB8c1e4UTA5jSPuSgax5
S15+pKy0t3k+uvc0S2rVdUCqEhZLiukODrN/dbYWk4Dxe+GocZA4GC8pCa7eNnzE
Ax1cSRqopXAaDIxd82Hts4obWFY5Hp/+H0gyhfH2bGq3vrVS/ZZKH12ticWKfvml
p2A+mI+REvxIRXc33D5pT0JL1p5LtmhJwuGAD/q1Zy/gd0LDbpSaxsnGHb38E5HC
A+FK6fOlE3EWWl7kWaSOB+EbiBZX6VDbMhkUgN7p8/XP4jXkQO0fKLo4SDVXyrsZ
43TR6Tc28GcihbseKs9nfTpMyMXEdTTXjDJNvWrqrD+XBDUbTuRFMiNg8sBMdcP3
AI72Z8QQON5hufQ2lUFOnp229m4S3imvotxHqOmZWt8DdvjxVV+4NJz7bt7333v0
SKRUg1icr6K419fJZILE8BuH9tV8nsOsU5peKI4oy8CGdcWs31QBpGWgl4elsC95
lDjxdj8CPCfvHRHG006yWHSQOn/4XrPcPGMdfJR/h5vAYP2HYkSyXL1yieJ0bRT0
rXf9gXS7odOv1wKXe0eEZLIWkqiDuB3U0+708olSQR4E/P3ijLxDKDBgSTaEa4/M
R5XQsix3UzNuJNwGtHs/m4203220pVcW1KisT8h7jGwv/oLe2TQjjz00yjGYkZui
/BTfZJIC9wLnqLkB9WTXg5O+D1WlKWYEJeizZeFZCzoe2q65lYPIOVBnH5M91WJX
Y/ui9bTwZVg9IXfczvho/9Ajmq7oVzxLb9NeGUyrOTYDyFd2p1OCaWFtqymlvQd4
rv9rPm37J/LsPy/MjVCg+wF241tp9bj9kL7iLqZ5ygRryJLc+q+jjGXVlTLyd+HU
LLk1fXoepZOZg1yv5VOYaezWRj/T7S8/axauCyTsEbDD54j3ExwUpm4gvUtguagV
tAGGzFHoFxiTDd8lcrzKIYtma6xSbmBuZ+rybviYVdHXaSZXIIWLLu9D45QvOOvd
yCKD0TFSUgivosuAotvnbi5bzxPhLprw6S6kE9T7Rl7shOCe6Zw0MdxRhli9hEbw
OHxDVIdZ04EMwYKrmW8I5LaqU0sFkmg8Ks0CUknJSwwxIqYK30P8jlEJ6SdmbflB
Fcnqx9hI8HP1idcCFu91/uIWOTKtkZ4xRttm9jNAaZc9qSxb16Xo3lcFI39DdAB3
ozPf+Tvy52Jvt3Gyb0vvnM66BggwzfQ56bv0pG9SeThrrzHqBieXnGBUJASyLPx9
jydJS4F4MUbK4yNMdhNC+uGJAgH1RWNaCjwJ6dtALXFlvQxhte/9Hahwa9b6Mq7+
Q0lHj5gP+BxGUHnLYm2MXgcqfofZT02fGqF8339GXBmax37amYlZ0gh+DqfzU5Oa
9nSIOwpMs/cudqp5PkKbU6ZUoVjkp/LH4/oIdo28OAN25G5emVeKLdJ2O0uCxdMO
eddXSBG1FSaBUmefgP/Fy4qT1WWiDhci6O5OyUIosuEDDPWkJyciKDkLusTGFSM0
Z0Tlyh5J3FynNfVeY91JZpmr+VNALnOcmpE9LADU7cOieyOQpRrFZPpxUZEhI5XN
WkV7B3UO6NdWUr3YFNAYyAHZ4yAdqqqGdT2FPoTFm0LYBGvqA/itMPDcosVXODxG
s5TYA0BIyjgdvunKRhnZczahXKWPc6U7J0T1+sQ6jm5kvyGZ+ZsqyRHsDn2ItdJX
sw2L7DEnD1gsWPKss7JgtWKmh/aCmc9mI1rNUQfRmRKkQ8EGuNp/3d7OGRswycba
rr+XKf1OuXZlt9ix6bojHEAvdeDEHX5eChBTfG558uo7opIyqFp6u6PBSgtnehcq
Drg16zLfIHnJG+KaFg2bDf4wtHhQ4DPwYD/HX6JVLJKZ8sBPw+fLGKF9xvm4+rNC
9zDK9YiQAJ2Z3MtLkjAyfyX2ex5XPzbqKa8qCuUIuWQQ/tjzQXxQvXrYFzx5pEUO
lO5ecGK1LtMwbtqViDGkOGJG1HYljOFy65T6mlFIpQLuiGnZMTODDEuElGBdFTwt
8b+4hcCd4IpGCuCOLrU3kBXT0Gnm0JiZEvXDN056q1YqDra6+pz3gY7sG4CJpU3T
Xnei04Q1hkggx6kKza4lXKxHjU5Z7n9mBpsZRCewdavBAkEdomk3Yz5HhHET8Aj+
OHQ4s1QTOP4ppqxUN67FR4a+epPpcKt1V9cOeyjue+kZyuoTPlkyV5xKb7fH1VAt
L4u9SiAlZRUe/aCEKzrUIE5xoNhTilP2KL6JvBxRyPYPzyvy2nyEN8eGYlIwwptd
4jBqjfygAag/4q7sXJ4PRrjYeQNoGuLDAlhKgod392pzE6dNxhOOhZ/Vw1ThVGOT
SqVIK7iRse/TMWtxll6k597O98vuX1LiJXIbv0LsaXanOh80cyk9cyn85yuBE800
gBpIpqTe5rToedezHdzBaw/V7sBgoAaxb5x3F/rz1i74cWZFq953pNVWcYh0iXz0
O2qcSYjQX+BGz1TuuhrfhFwP75FYgTmS9PsSUak1/2p+x2F9K/94sEUK3y9v37L1
dpJHqmT3qVTcEjCBSAXgvUVyM/qq9H+ZX0ORRt4qktNy15y0NkB60d8JSZ7td3XC
aIXqsmiR7JZV7xjonhzHhq6x8VgRduIYb/jBiilkRH8a182KDYzZpO0ZxZdljXJ7
2MbEtGwjRi1zONZOTqDIUa4KI1TQrzjLcKo8Puenh+8lk/iDz+aX347M3YGSQmSc
9SP/PvfAHLKXycekY0dfQO/R9eT+9ULbUmbvm3c3lUluaqvukKrdo8nHcW8Oo3fW
1QZXHLfqrU2x4ks6T++Gh0cXQBnJluGHRhyzvA7lyI7lRsrsueATcK2tTkSjNvpC
1Uoav7djbLG7sYmt73YGMq2vJqN24VZMLqVo0e/ISJeBFdiwOT16v7Ah5UB6IY/J
MdMdXpV5vJ+ZlX2aN4cOXS4tBI6yC0SUQ6YDvcbk8wH/fW/pjtk6v0o1t3RINHEa
sdXk0fTwjwl58Nsy/64Jc1PyYvGi/B0yaXF7kXzyubc85qX2/pNMXGi1iKbVROV0
i0amqcc/M1dTxYK4IBJcq57k8UIJh1LIpsRo8x42lbK/n0MOrGV050hxASbVzZNL
jAdSxQzsigrWumdab0rf+jMYb2wIjzTBtQ9o1oXrJyzMCuKpd4tJlZHOXn0E0lDH
TffJVlpR/ZHjWDBZStbskHikSwGK/lO22OtW82q+9/qWtZ10qygfCKNwzjAWVj3n
3l2zdobmAYSSDYSoCPDzSwpWIKZZhDc0gvYuW0Y2J1iyvugqCEu4tS2wmcc1fOA1
GgymJVTFdA3uh3uo+jEdtAmljTmepFNJGUWGvNIVhSROdgFYNv2kmFi96mvBPOF/
3nuy7D/3IoZtp8o1PJB6SqstS1qLChVCgfyNLZ9kaok+SacgaZz3DLbHWoVHjBF7
d2ABSHgwTQ3EEumISAOaX9CT1qybO6ezHcS2NDSnf4H4YOfrM6mL2RIFc/M2kwaQ
jKxj7UQ56pFCxsCZiA4TLRRykSQLIuFYw+bXnkv4yDwtwFoOAXPtY6+qIPnNZcGU
W4BeGz11e6xAjDq3mGnb76uPugvvo9mAS1dFJhOpF/H7QsROnsN1rl+OZoyJuo/f
Y3b+g8fQnFQypaBXrnVfM7++IRIiQbR26G2lwHgWNC+lT3ElU2F4Iel+Lk5eqaq4
4uE/lel9VS30D+auK0CcjTz6D8xqbxXGjTY52v8tlyzD6VUWL9Jw0JpRLD64QqqD
rPRv1yfJw683buVbK5JC8kQeUcdo5Pc3BeX0dy9ttWfBF2k72ImSIlaMFD6mhLmv
WkU8dzSHJpMtU3E/dq7qmryw8xbkYFWQd5LnGBN9cECFec6BQNb4Hzvu3xqdJjYJ
Sz2tVbk9JbAnR1fnVf6eB3cnlfm47kXaQ2w7YlPdgol5g1C9v/R2pda3r+sFJFio
YWawLFiIv6PUHYFO4eY2f16yvestcjlTvVrTOWOT8H3yl077PLtP541lMOVrkqCs
fTjIf29I+MnlgTmqCwZdJor23/FqQIZVVFdj35RrFy+111CHIOM3A7qLlgSX9lsB
vjiu0pZS3NjcalIVonSnmhaKS3pl2TJYF61sJJtn+eaEa6tMdLb96r/KXVCyb3R2
d5dSb8nVwwYvZaPn2kZxXHuvx/fvf9Jf5QNqeHnzb+9h6oFUIccghpVsDxoRjhK8
QC32SJpbYecyAqFpgUPsgT66r/75SnKi95f878n6wHi+NXb46FFC6RX+j+t3E8hb
G3wCDCbicM1s7ZQdQSwJNWB+AcJMBMGiIKLNGqP0Sr/zFA1FmhDhBSYc+Xap5rRd
chcfn8pjOu5EBb89x4nbZtRVJsAoNA2XWfSM+GT4ywOe7oyqKjfrJD3SQlIJV3tf
Rfv8irNnh/bqkVK9raBVA+qmu6bUOvTJaycxNwIbvgvyYAiWYZaWn5YsN2VPB8NB
LcyUuftJ3ANiL7LEacyZaayAWZ31p1Kn/XQQLqJqBalLaXHZnhHXBKE51gwCTFyS
Yd0ExUItRNF2xHz6kh+UHBcXK8sG/e/XtFSyntt0f/bnXxcubtzsXhJu+kqBD8SC
jdhWxzbwfEHGsJhvIGDQwCfOPbJxPRpjrykmr1fNWC8EkrfukhRCWP15caUZV2jU
QMFOxz1eWW6FAsdRBW/tIExaedUqVtAXdMoweXFm2XQYlWEt46BOBEJUdy1wlzpv
+7XpA7y5MKT/W4cRA/CvlGnJwrPrOqTWNWd/kjwEW8QvyoD/VYwjcUrsoRNFbk7c
srg+xfPO+719RH3oNnIlSGi5Nzxb+Hw7WeB9nlFEXnMviQNNZlMkyig8KzKoP2N4
z1XeE2P9SgoC/basCvdNoF6Gcw7ireLSyir6nddadNcPWaY6k5kN7ct+0kkNMqyh
PKQf9sO8BRHhcgsHOjbU/vn9nrKBSmGQuAgN+mkneCU3IvCayWHadQEWELpeCn2h
XRFlgFWikDfAadA++pzkfyyWLgiCieK/MF3UPa3Evk3G76wu633WVfQkzo14s6Cd
diA0ZFg46c8KISb1NcX9NszRfBB82vlrCU2Cwi14Z6KhEyqWxw3UcVQbY2UFVNfP
Q17B7n1p/GdwyRSq0nAyRaxJDqoLrvQaFFgaeL+2Gt4oZcr0O3f7C2nIYe1NTXlt
Siz4pliyDhUQE/Jt8WvJxlWqnUl6FXpdCtnDul1/AOGfEPe+J4Sgrcguz6+AJ/ro
JgzY1bZw9OCqL3Qw2GbhDX1MdA/fpIvHiZgQU5CMfREvwbmjFKYJJYozuFs2oa7l
VX/l7NgAiEr4QCaNUXn5f8CR4DEqqsm5koNiFb9ow5Zu7bQGfmVBq3Qh+zkZDuqo
NKP9TnPmU+CM/buI/HaeQKWetjU7rHGuSw3tlO6SmMhYmCoVz2I+pTWOEe/oJeni
CJurVIMwvoPBCEn3Gc7BAJCYzrwrrPlCMjKfPHX/ZfU2pujSoGnl/Uzf7imBsp1V
DWh1UKjSREFug5LfqG4SpngjQAHrb+dduy/tb7z4rDFTWtlLE09CIYBEFyQxLgl5
o+cyFBO9m6VWkWyHD21btCi4AIpltmjtGTudCaK8wZi59NN+LzdGMtjFhYIGgc+b
hlnjNcgjNM4nSHrrvjUiRy5LjuJNc+Rh2g/GKOyJxTl0XdBcgUYWPrFIyJfvIMFs
BclWIxHqJXViewGTsrVSIRlJj2GDyffB4e/R+MA8/3mZtPNtSpTUmtPGaKFiW+/n
6CtPN+kbUmR9eZTEcjaeuUA6V2yUgtvitViPVG3n/Xh0tYpel+BzujjZlG8YOkHM
YD3xtZYr1597GJypGAiCg+WQdxeAnyfsMRP0e5SXzoLZt8amgCYvxQcQbwaqa2UQ
XfkTcMaesYCxxWVp5iZFvotVuopNfdIMuBBXGl2ahrLLdRtYDkhyI2ABusuKg9DM
OfkEzxPpvXlDjirWG5KHsugpbw7yXeZnh5+aF1WHowBn7Y5h1AfReachSTy8RC7g
yKESBbEsuV4Y8kh5KUS8fAnUKqrLFtaWud0/9bpKHb34eFdjIQQZBdS8BnNnVFtT
SyFZ5iYt3V/RjXWWJpxwKMFyBTQFRSYDTfNe7CKmudDMML0QFlrpax8nRiBa19f2
nhjRiif7k89TFMUOjLcMla6F8mU2/euTFnFdXyU3LO2HTHvudEHL0jO2GJAdW7Df
+Bhq7mIx6VOn0oNwvdjWAHOcm4+8kskLw5lazkXmAy4EDtmz5/lYyHVMXMWEDFFt
+zXHjwfG5TIVa54zJAtYprEhxjE85Rcx/lA6huGA/5G/rGXHy6AhM6AMJ+8RRzrb
MzNnbTwbno6asQlnX0V+x0qlCGZaQ7HN9lP58NsoALefeQynksflSCGYwGkI2ztJ
LWyQsbFqWAYguZlFl+zZALIoV1RmzJhE5ZmXLYe1SL/TVhoX7W/AyJHNh3S2IHi5
7W6jTvAUleGUviGJSTDQ1/X37hnuSkpUlhTagoAS34wIiEanGmuDFepL4/R6VzY0
LzRFk0S748TnMO9TGaM09B3fQr9uRLKfOFvhIrABHcE5hh5mL6v69a6CM1CJS462
U8myIt0utf53HKfj+yReL9PmhHZrSDlWgyXip8CAE4427CdBAOuaY1/1ILzHHl87
3KpXM93BHCw0FmRuWnAKN/2ko1cHHBGDs/5ZMimKZRX+T3l5MAgaTGQpnFiZD5y/
NyS9rwu6+nmKWL2Cq0y7K1uRrcxVGqGDh4YwWX7bdQSoAtsTi7pKf+6MA0F3kjjM
KQOZSSzgJlsN5BoWxpqnNR3r5WQMKbNBMKQS5DPk92PWPjetbGsenHg8cRz1wA8U
INyI6rOwJUfaEcmUucSa6oXRz6EYlZQMMQP05Gc8SJZxLevI6h1jED0beTZbrJvz
PxsKYy/vrsX2A9T0TcMbY0/HuHJ5D2ZlPAk1JDZX+Ix8GP0Vr2KEHoqXU/iFbT5P
Y3lQajenztvHZFzRO1lpxWLF7a8RU4wY++eydraEmhEToKr7xuTfhOX/eR7Ihj7C
pML57t+HiJQ/dH+B5O2r8wBchAJOzJ53jE8bs9pL5c1MvqO7kKM62Ovu7Vd47AVt
CnBP/wawj9Q/gn8cIvO8BAPmDsI2e3lTCZqZm75BXvp2geiIRqaAYmd+aeJXghuk
+Um7RbDdnU9pxayKc4/nVBDMjPfRAu3MJwxrvNS9UrZetHYElzeDjtaqmnCsnIBU
qzmJRxmB/vrInX6Ddm0s/QEph1DFcHWtMEd1Y7SUe3CQD/YYfRyuRj/JwyeTmnvb
jSySKZJIgqZE8mybuJXv8KvdJMbqVjVutoGWEHKSZjPEJYJJJ83TNyHNq5wySo8W
wnGUXy7ze6m7Ctag1WT7EUy3/6bO24MaGsavSxct+rcyeH30JdX+B52WKNRPhq+E
jnQ33AUBeTW2RRyw90hxzzyExTNblTwFXhA/48xG/bK7pGT9rcvEBFGAtK/RKRVX
0/M53k+gHFMqqQYh8o7r4GtWO/+79aJoNVNOvY1CVg3e1eKpmCQ3TMMpGuUDCIgt
kVeLdBIvt7wJeAuTlCmIpJHcP37uQtnkeHSQq2s2wbYA9Tk1u4P3y1+V8AVaLg/j
7aw0H778kyTW08tGO1/T7i6TiL55A/CP0cj//BVIKjNouiXOiHYo7a/3nQtmC/iO
wF45kzMiH4UTYkMgM0iS0KIDT7PtKqpgpBx2b4cAQdI0uwQWEeU8/RgS8ZFupxGf
wXn7y8IG+/7V1yE19Fu4/skM/nO0kqVlZvmHnQ0wE4ciPsEmpSxVglacXiDltU86
n4aAiH/rtMYM0GR/DYyVciOU6f/XYtbHcT4ktK1HYtW3+VwgD6WaG98EsMXfQ2P3
qGNVrurdDQ2Mgzxi1j1O1z8pMtYTY1RbfUTK7j1i90w4OLWn1qkENXq8r5dd1szR
ULBi23O81X4u/xQg0kOU/UULbkNGR9zpW0KNbuOL65cJa9eYKTph5ZCXmwabhP0O
/VL8cyKJdN+db+2XY31Hj7ZWaRf7DQlj9ed8qDVAw0pW/Y1ncp8aNui7AuBEK9zc
YXMA5c18IKHgZzkeloRZNQX1ursJ0YGQS4NhPU4KOS8SmzaUyFAarweqP+FtnKEb
uToZRIGY8NI5r8uYOCNjFcv1krZ7y+OM1dIp8y1zBIgMfY2jKAa6sSzTcSQdZyQb
rLkTJ4ZxCjkSWmNhqADtBas2GNkt+0Nm12CKZFnvSMAL40bmgx/tjbGFp4Qe425c
iVOeR4fJ98ND0rlX0L2FUo5RS3iqoo5qglE+BW3IilbXdkOzYdZ5WAqGY4H0Et2G
7A629VPWB6qB+AX7ijkLhInD5mJDPbiIp9RpLgcoNwLXKMNDyFtN30V2DJUGDKtd
2JMU/bnrzCv9jO5j6FNpZLjCKOwqbyBBV3FVzlbFAHUwAtCIf6nx5Joyk9nzQtlY
kZS0GIkPiqt7AiCglPhU/pXv8s4wETp7oLrfujOEZdutL9PbUC07fEhDDDzIMFkI
8ysfWtYWCpji0TOzfrrAcJ3l58SpOyFgNO4db6AKVVdeXjbMPT4vo20d1lup4eKI
A8EkF+TaP+1xyido6n4gn5xizb+cNDZomCdxiTD8s5MLEalk3oHe5L8JJBLsU7pj
1vscAM/gifFu5bGmpuGTboKC3W/iRn3mccAJlUn/nL3ymgzcMD3Bg2n8YBASO7CE
LVlBca26VBe3/+PS8dKByNazqNYXPEhGHsdLUNH9mUmHwimkXDGCJKP2af8dyXcV
jzFHzttEtxxq6741dXbu2mOD4XHm82rzg/Qwb3qyHHBFOItRPntze79wAqSDunhp
/mb6TvREthy0aftiTyo1kvruDIdG2JHivdhHMki49UkLOpJIQeQFXZR1P7R7An+L
Dw4VgMoRw/MPDz4UTEwGSWOpe4h3IElrKJCOCMNcDbPdCIYOlhusSzm8zb1P6BrE
ozQjW/9FioBrPJLie3yGgJsCBz0UXevCEEDEyYuc9Vd3UkopHIUBV/kmKH17FXvF
sO81N65JITf4OPXKD42goiFGqE+MrNxKseM4FVh7XxRM64g+vyGkyOZgo8xH3Qer
Yp5u1rcjVhvTVP9HRBN+88cQu4tOwcySwo+/jKRUNBdZagBp1g8E7V1W4R57qwWU
uoR4GndeZf5+b5MftPrTt13SRKkLPGEzJs2CjOxj4JPt5Cb9PM4yZAB2vu4BD28O
LOb30dsUEu7ahebLGbQUd052SVOHrKo09sc5DX5wx6pUhRP0wiUdTSndpg9p5xcm
9yeUcllPnFtJtA5TP0jWf6f4EiOx0Cyt7yBKKso6Uu8Jb6n7krBtiGxAi7wdUcv8
J+5lcS6QBWDj+eITZp0zYMnvHGa7E3jM/GusPmfaZ5LDwnqFK1+mrg67SdsWnF4f
3jpDNIUO5ts0Miyn3e84daggRnDYxJOpIKz8nB/DUjmjCNI/wC+ZSu1rDWQeyU5y
b3DoMgiUnldzTPfgofEXwGybCBy0O9vmmamcUqj6fCPMHeMv+Zz8/z+TWPaR+3DO
LINKWc4iykrg0h32YrR+JRp9GQy7HwQXfrnDD79T0zGekt+dk8PvXyDLv+EDF033
TWREQrOSm6sUTVhXmUqfzi3BCmW9bsFCcks5COLK4UjV/XNHSLCfwZff50LN+eOi
KKWaygWSYWJfaRXDAPKDbKFhU6NYCPzNopm4TUpUyFpX4bEmORq44lZwnhDUXC3x
P2JTFMl5Sy2PRMTHByUITMzu+HyybQCfFKDHsp5YtRx2jAIZaPLynHQCZHYAf4zR
aelG413L8O8OxJxdXVdsiGlbgjrdx7fN9iY67wAsrTJOnwMnhPRMMjsjbLI1bXGx
hnhfwjs7FQPFox/fEKMeM2KI4M7MEYdQC/AGpfVa9wEwDAGoiZRKOEF7jbIwS8Mm
cGct6D18PqJzkpMGzyFHOr4QsNyw1hFUwCzUwggcYU2Z26xes7qssUeJqa0MrsP1
/qdZMSdbnO/0P4egCyloZzTnwVB/7hNdJ+iA1Ao+KB23g6xJO1l/EdqI9dXmLYm8
MN3CxvupnnOZV/SAA1uBQTHfkAWNFjflFsbFg7yKG0Uw93HCyUtaOFZOvxnScNBz
RSfM6KiBO4cxSq9bWQNJv/P8JuL/XpQxsLzh8/BgvEFGQNoLxD3kWiuUWSYFXmmr
WtAFmpRmbwqBgfoJjE45U1XsYficHluOxKShAR/VRa0ou9haGCcOCedYHM+EYfdQ
1eP5aPehaDSvqPLgh7QiLb00tGVYa/hhZaVrmoUOXk/7y2euFtKu72vozX5+eE3t
sVWAA2+BTbyQ9lFyf8fMoZIXXGCauBaAVHsG/Cl+Dpz6EMjrrAnWtZrYMTEV4KIe
uSOR4U4xVrMrzbx99hDbT+nPTAkFR/0osFZ1HdqwlmPTiEDj8d8df3PcrVtZj0+M
jDW2JM1aNRwOiCJQO1sTqMQ3RTcLNEwiIHVWlMErhiELrlvxYS0DrtoPFMYTul+p
iWY7DBEG66TEVAv/oxyijrgBODCVR4Nudao43pqPaQcAQjNRGVE1p2JGsPox/eex
Watt+TyFfijdjOKd0ZJ98cJ87Gup4d/Y6+PbCuewbhDUYsFGxsAkQsLZfgNMNs2R
5CWBU/xGsqs0k8k85riFhsSDjQVzNrUnKYMx98DVQXof2IK9rwTIqBbJYmC33C+b
EpFLOVi578gnVuoymYMPBbpDjjTrNaTSCfw6A4eSl/+UW0Yl51qrkEoZyBKV01D/
fjfnw1LBVFgGZum5EMZYqcYKu7te+LDjcndDRR0vJqv6pMTvmXJbQodiXt8uE6ZU
9HV+r9+vyT97f1xVQtmNST6PhuIFnbb1mhtO8RmmNYJEqZaX34hk/qLNvmXUr1j/
19SUCDxgT0835zEvBcWpMXNTV/jA6Sf9LIffnxceK6mgKEDx9R/XeukWCZUo9lHI
8PF0T8o+Gy4LK6Om2yQYOjLjgiYrKqW0qG6s/uts0LE4TTW/LIq/CYi8qkRe7oPb
9OFjnhgA12cLRrDRLAGjAL/aLRdEYLkRhPVd0RvtcX1hkBbaPzTPnQK6FzwsJiX0
IpyyzBqiyL03Ck3pas8WZDARbMjaAgkjrlk67lo594BarlWoqnCJjmWw4xqmtI0T
YpamKgehXddWjf78XSrvJ+qyMKdbbtyQDCGGMLU+vCekO0wAWgUaI4RGAqdfv3My
ui+3G43uWYeTAkxxJDWv2jg77ZOHXMLRRiagX9vtj72kqg1nDjnHLocusgacRgOE
Aj2JHg8Rv5TmMYVvke6Q5lfaCNJQgGH48DJQNaePO7msvbMWDDpJWT+5mxcCqcW2
VX/y43J2tT2NREcrpeB3Ug3I3pPU+1qZ4nGvvkKdSKIKeJYst3g9KSsWtwuwtiva
dkRdFo2OKZD8Ggy3bVzRhqxbkADD7+v2VZP4F33SOO6oTSF6/NWZIrwexqgSRxY7
ZBFM2Ghe9mId8CQm1LlKnEFRaTDSFeWRDoO8JSTmhd6BXtXG5RYzSJYiH1y575Uj
z7Bavhj+wiMs8ZaJNwp0CzwY9ZfnhMxHH0yALe0W2mWQ2MzcRQCMv14IExgQ4PEL
K+E2Gy2HDl0W5UuqXvRj8f1IDGDFcxznslgZ5ZdvSIA3GRqcxTY/w5u9kZaVz4Wp
/HQTGR9S/Kh5Q9dY19OlyE8SA7KhyiHyPdXBeLqQITWtqjVGbOr7yuguKJIgEFxW
o4pwoD3Nx4NOrRKl8X2JVg4j26gBu/Ui6c97hxoe+UhmdM3PyJdQStTGTs0nUURm
pzyn8PQsBweGGFxkhegmBAAaWXQ2KdhZX5DLMsJCyU5aKYW+4T5pfrECwuwSXwvm
r9+vJPwBlPpAZCr8Ys6FxITF9g14DYrduvQCbWLbDCPHo+WgcUIsBLZn4HWa70af
LYtD9CEprWcbSMF/DECpt9DVL+oMnO54IWFqyg4TWp17/wZX49FBkDJYErReAlb7
q6lNsq1mAf48FQnKQMR/k6fJCedR2DVY2vNAEty3aD0AzlBoSJVqp/1vwxq0QcWr
lsJHMvzk9Kau7qWLdl2pS15HxX1bjswJ2+1sJbJjXGn1r5t1lTM3N97Ho3uxxlf/
5jEKCu9X+A8vzG7mu2VqPkGfTJMTJck+1lJSXrCdOFtzvW/xjwPbUrPTp0zD8kRv
/uoSi/UeuY1TtPTv81tomDKiaO13vOG3cZMaGHLm5dvArApG9up0siWMEAGeloDF
fO1CqhtjLld9ZdbEayA6Rb9dddByZBeS/OS63dY9dIzxIrzhbJvdQGEnii+qYKiU
JQpJlyYC/SI8dFmwrPd1ZSLQ8ljA+1HaPUYqlg6l2n9I3r82A89F4vUReJpKKqxe
sj0uWAFExScAvraxxd2wRkifv4XmqKjy4LCpHLDs8Ipkkox6EvsVZwh/L6D8S175
mmQKvHNVvhCA74qoqeFUeFy2WpZBtS6Y1X/jU/DmRxiR2HAlJaWWh7IzkEUOitVX
LzzIxiCWgIBpMjjnDNgqlabdD4GriAt13cj4poJWBr5tc7wjoEWXrYvpqKK/bkK7
tLuTCDPJVXYbF6hfAsc6pLzgPWXSAvyvy3uSKnciIcolY0+UncqZdCPtdQKtTFk9
V6dng/Qpq/Mwluu7hqTgujyv/wM5W3/Ue+zIyO0qiOgmUNwTi6hVCADcpmhv0oHa
T8LqSCUjjc1PAoigyPOAGVo3Q+3nZlnlHYbvfIe1H6EG+7yPeHhUpWO3kqCyUuom
+OeWRM15OI67hmtL+K3rviSzjc4AzVdadV/psPATbAuBKYOziNuKEy/3zL771b8u
+AhKq0xMI/Cm3yTTyUH1bijy6F9a7fQGJjXrLoIvsddE1ZQukLuXTcA/nnmpxZfv
JB7aNAk0iJ9AyMBwSlzGJfsakL5KVl8ZmvmwXkS2sJp5UXTkn61wAjZMAr3DNLGI
hczFZT7ZFq5bWBX/Sx4L+T9Qb/pKV2rMLYgkdMu3aNV6ROfmbha52QlPFvepjviI
F5pNdUVFzmWnOOSbEYkhgQd/QO23jqx84cTN0/LdDjJ4b1UCJhqsvny20airtx/0
+6cmQvmhEQ0BrCNc8eRFKueoUb7GkpZa8dyWJcAgas6feaYJs0fYsIs29Re9WRbY
+TQcld2OR/mjhDz1DAYUP1A/qvVkHFCwZy+X8sODwDYQYK9rbrAJUAiD2C08lFz3
80inD4q1bNEaNLd1AEmrbaRogkUdKx9Y7iPALwRYjPVYFDWD0GT6AW5lkO1arl6s
vEHTQTRgRryYFkCbeWVTMSAbV1CkrXPeXOgbYvarMABrEhWLUcDtU4oy7wdgm3x7
3A42tmNfbjTqdtMrRjQXHuUHAX+EVwspeO74+BXY6irS7ezLO3EmbOrDxmXI/44r
O6WKc+gmkrGyo//iPT7NPM4x8FKR30c+MVatihrlCs3lrLgtbGKV34vDnMWYdQ6g
CM0NVAaM6VySoO4vA2rlhzhETGTD3fj2sCq0/YthmqHSFrjaDzzdE7eqfUOHBxTr
cnMIw2pvkdiCqU7maEOgR+AFuzL+ONaohnV7XwE+GFbS3NgdOXnIRrI124H0GVzn
9mv4q/ojtKaqnqUhFpdIelhT66ljPOQP6/QoVbQQs6r6jHNypZBkyuhEONlRnD/C
KlwCF9MAytNfkGFGSy19PeIsVqNcYh+sDQ4c0Z4PuQCYK/vyJAanZkV/+SrZi1b5
AMvncILcNSAiFt7/wNpF7yHsp0O7BWED3MOcYByFl1ra6EhFjXVHgB89OSs1N2v+
Gmg+dDTJ76anRQRzO3M3sYU7ThIcJyaq55YddpYaDGade1A6etq/r0LsQz2Dc1/n
oCC6HEuO01zY7+MhyM+cJv0m737EDTiPNmgwzpBj8Dfy1BRsOCYfev5Ernoj1End
8MEF1JcLpXhAJWj6fYo9UU952xN4vB9ewrnaZovH+vw0MNiDmjIbd37xmszzlhax
mOu/OYtAVDVLY+HtBW9v92SZqITCA3t/SOM/TrnyVX/S7e/E2gZuqZyL6SMOkiSh
MWXxzdpF70lCeV7NV2Ih+MuKQu4JqLmSRBvjshm1b154P3oYeq9hIzrm2ewZKTu2
PFipmJuWS8vsQWc9va9XYuUFbbB9RrV0AYMtmnQC88110WlgTPisz0pWgZSAvOKj
uKk2BUA2xZbzgONedL5k+hWlZiPwFszu7iPa5b9uVBtQbBZxm57KQaAIl6Xs/Ldq
7DAtQyhsgF1w+5cpZdl5/9FFk9mlG9Or+BcoHVLlQHdJ05IWiDykIZZhJVrqlrKU
CUNUv8YD8zolLmnmYsRucS4CT+v4R4JXMDqBoRziAqA=
`pragma protect end_protected
