// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jK9VYKPLrYcxsrok16Cil24UO9oDyEoV8sMxFtmIM7arPD0174jS2xmrpFdE6W8u
S9trmpiJM96Dr3S6zRNvBY5suERwpQKS60cmmYLUbu1htrxX/8cB66AbJz9ZbBc7
oHa0DJm0BIbqVTCKzQ0QHS6QQC52lbPYljZMQDCq1rQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
0kzpCVtDgxPTLrW2DUp8CNOpMAmi/KSaV0nFfN+M2E3xTv7QGnPa17yLEfnaqcDY
A4EsdhO0UhjQNNPYnfgeCKVPOZoSXyiaa19wB9yRSmFs2WeLyT9R5wtdUFugNwmM
Zv4ma1yEx2B81LHCeJisxEefSeuuVJlcaznL1slnnCp8Vx98Ixi1s8g4LvFbywAt
vxnIB8Gf9iwaELgpskZ7TOfe83372VNGvuzO+UZVLhjnh7aBMU/WXX2FtlXODR4o
JKmaxLq6zz0ptfN5tclT2D2SNjBAMN7hr61e+a0wb9FrmQ2oF3c5Yceie6LbRM7Q
YAU2XzgXp6kjNA1gvfpZWl0H5kttIYC0x5WC+jjXyXCamgIe8GsEunrMzbiq1U6N
/2KwhGlHD3FB5zdHiReqf5e6xgwSjEcBU3Eglowj1Yvx/SvA8BMjGY1/X/gLJfGg
jqJRG460le94+HIdM5SMRZq+KXuiPwqCrxJB94haF1AgqqvGWyvlHN1FEtrIrRGC
gnXIV2LnrRtpHpmDxn4d8UJmlCvz6WeGgTbaLEXVV63IwBtf7npbpGMezAHGHY+m
eW+9aHdrLGuZOKcyJNnEQa+4OW1zrth4l1hWnRYZDm7gqQGeDgp4dD9hfQ+fSb4T
GVBE0wHORkhRddO4TMstrnaLIZ31s/htFg6QDrpTBzH06M9eKWSp0QQQ049hEqwX
3xl3Gzc9RCqaIu6LHMQWi4FlI0QtYi/OVKZAMs/psdsryTdjd78vScqdg9zrxQcd
6yjYRAU48wqir7SAmWRwlH6hJi8tRU497UOJlqDjIjS3mxt4r0wODQbZWFXBmk2u
drSkL9CIWhwFgFYqEx4dlP+AMc3I2iRqs4JKauBAlONXygALgW+eeK92QuGxT2p5
hn5Rax9JiCi8DmWpiqjfVQeYryD/vJ5AZ1Q80HiRfsbCc42pOlh9GSCkS8dbo8NR
f9REdW/VMddWagxw4x5b1FGnjVG3GHZLzIf4Q8iVftZ6xrVpEO83CNA49ki1Eogd
LggRmTqoaQZVG51aQtnJda7jISnq6d/sTSNc+t1LhdylLQrcwSRbUB4zEK0dLYU3
IcWQAl+6xBebgL2tKEj1IIXFY0+BtGUDPkNRiB/MnGIQqucn8U/fukrWT+qDf6VN
N+Kku04YSvu9RwX7GIt7Cq7jyvzqdwaE85GrJBwI5HBhOrYnNkHgQgkkCT82qF91
khijrm9yU75wJINW/zsjB3hht3Ohg1elO6e+JF404eCbDBHyHT5SOvAcVrpQfjRa
R8YryD/gIxETMFoQ4kXUioTNbaE9P82dEHsNU4W3p0dWqgbfWCLk/xWVn0JZXQS5
UrQFq58BSTSXz9HOHWCW/ISRqnf0DdERIuve23kQ1GonVCpeRAlNAoS85niSzP+o
DvRUx65+OthTO58wi+XS/FHgBgHrFwNenPd4gUfF3dGMWhsqbfXLuwnhz3jpLhIe
ZoKQmRXC8qZdnyaZ3Wv70KwXuguodpeFJDJ3nrJqJ8+oMXlQ+Q4xp4jdE8NnKiKq
Q7q0LHVgkdzdBW9wbQRw73bQkSQv18Ke83IsY2n2f/4xQw9KnTEX+rtW625qdy7P
vKlusdkiiikbsou9utPTky4yjrlLV7QXpu5/Xc1WYHAsa1AWoddrzjH8rLMgPcTz
LmA0XLbEgVt2NXUUXOxT8Kxe4PWqtqGuPA9YmfR+lR4gTEVrhFG5W8e8lkWkuNcN
6bfVKq5FnL6YETIYG5l8RGofA45SWNdMRXsyCwlZ3K50D4AyK0hwBYxWc2z7e8di
v/mqqeF91mnKMF9arpt0ol7wv848GAd/N9BTFSVr7P7otbtpkOI5Vkxhuy8Gg6+E
lxu6RzmGGSm2uoo602F4041BAobZZrPJiEY7pmliTkiin0ie4aDaQwKahoYJtxn4
fW0Gpf8tK5e4cuoDAAdOn+qmR6ndHxTIO7gzY/RkX/3cLwZIIteqSUXFWXEd2s1l
SJLIFsZzoF3qauV7WLHquuhHI3Knx91Tkbc1t2iMvnkqMzpZ7KVFnxUFS0Gn6hN8
7ugrF7aLxG/ltpPAEEySVMFI0lFqrqVbvt0ggjRJ8yyzYKw1pP0i4y6K8D2fwQ1n
OX6HhuIrOCVGHtBADXNA2804kQqWaddSFcIreFUPTovsXm/FgfJ2BU7hsHtniutG
D/ixq1znhzdne/Y81F2Fki1qIQxWb03Kko5bZA5S3WLtpClXjIuDKUqFycozhzKo
vMjJWc64s1ua+tVA9dl3LoaQkJq93dK51BNb8L+7qu5Sh/4e85tYaUbcVYZPTNky
ooQO8WEqCevlWT3ug2Vuf9kJVLNCMtUL9ifFAAPK8bVbJUfqi+Rqlc8yhrAb4/ch
kM81HZbf9AwUeXyq8PcQfKBg22tWLIIPLY9oN33eMIQ/dWR+j3XulYYO/fA8ALs7
0vIiDSnc+UXMIaRXg0jXnzfCavHntFrwn4dPLH68N/vJ3HAjP/5Honyr1DJD5tYW
7QJ8/VennHlFld7uWl5iPaMtEayM2M/tnfV6sEYFiXOQyhS9xaUDaYZkMw7/Poex
IDhrdiBD31Bv6n+x7E/2KFvCucHqigA/EtJbVBGBZD40ozk8YLuXgoZh6Gd7R/l+
TO9c7B124O4m6WZYIKvkM8nk3Hf009MYoKbvw+2Fne9ZmBRzeO7PnwwPDbPVP1JN
Gt5WF1WqTTsgp236W9UG8kd4M1xA0k+tk96pST2MqjwsAuWOAne3RjQuXiIQxNpZ
GaF8tXmV5mFtG25M9xyAWmJOAhiF/dsTn3Spf8/MvUFb/wBe4umYVvY4s2wuj+Ru
U6qQbTwIxsV37iMi7LxU61QIxtNYWvzj6R3ij5ApExN7JYppGjvvSILLBB2D11Iv
PE9QKum1cCoXYKhxY9mqJsWGWA2rzcgz++9pgzu+RJwSWj5rl7IaRgtn58gr4Hes
LxBpWHyBZEC9WbgfTO+IAYf9kYj0kSoJU7yhNdkjIG6CLctM0lyjykohipOzhqmr
9AOFmmaUaHsVF/+N++x2AjDzupyMpITaKCAG7s0QC+Djz7BM85s3LXwVpyL6qWk2
2BYvJF5b3rKOdkByIdPXLINFwEAdJd68KUrlkcmRAcLOQysDOKMuOYerbq92B3Ek
557sI+WmGvAGgADF0aTU3v6QWLK6gKm42Yvaucmy2VCvC+BdU9AIOgvc4p1FkgwO
9zOSmjWLEy238I9a7TyfwiXS4XZH7aHv/ZyIPhXcGaahuFMscV8sIMYWEzTX3TP1
PCBxlyLCt8oHidkFmwnw1WgJ5mW9a+QGlro47uagT9yA6DBgfAph2s2m+6BekFiB
VT2LLQovrm8P9KSL21vv2+Z/4mfeQMSIocljLr56QwtpS+8UbhRgKE8yOmM50I/A
2UQeEasq8OKZTPEqZ4RwSL/dcLinFLTC+58OArdQnLeCUWUFkmEtUG2rt8g3h7ew
8+MAC7ehw2305I/tn/kXkteZFahKGkYYe5Fl5mawhS/jCuag97UVukgmYsFLdRqt
jU8HEhAtd3MMUjz3RhO0HKFsFryHBs04BcRbqp8iYH06U/UoYd90E8BKD8VTeFgH
CZ7Pa1WIfC1YcNhQb+bFLPN3tgUW85M6gugayLkUZc7isY7jVx5F6GqCDygGilQO
hn2xvFisaQumiSllK+hwqF/MF7IJp1bC2/aZyLojfngVl+SvmtndYLmjSpAEZFWk
/M8jcJX1e+vyG26nGKettmBWONUNQ29BCm4N94C7UZHVfC20wG1s1/HoCZGBG87F
EseWwW0wtFeVeYfTIvXGCANvJ/bObG7DeV9d1LFj3vDYMbdj69ljIMglqOdTkGgN
Fxt+ON0jD3S4gBy5VmZ3up0syaMUWUubVAsCnVBNMpxpcfyYel86Gx4O5TrfraSb
RHYYb5Qd6h7Q1PcjqWMkEjbHNALQqQSgEe39smCDS8tu/AzdkpN0dUafwRSm2TJn
KRX9vGpwzdMQASdj7lb1Qoyae35PewEMBG2N+1c7WWU7WoUijHfV7DpEnzmaN8zX
a8ilfSTT30wtWEYRbw8BAFBdwzh/q7LR45FSU7tB+t46jVeLyA54RXDtkHEPowzN
VLPmQ/IpBwYm4u8FDaSDS+taZyXLGlj09Og4LU+D3fXCTaEoKGjvd1ripzdYrUzB
7462dVSrwb7cSxCiz/rPqKgkMqh3sG55sg1cGgvdR9hSy4w/XMA8+Nbixdh5Rlez
3v56rHsxZNSjbygPg6q9ROBwDRw5eCpIbTnIwqg2F+Yqo36p4f0DaqVazTe5ISZw
/mkXp1X9TY3KnipGD+UOtHt1M/ldgFWXSLGvVx2Bq/LJcx28Kc2SdaoXQqLih0So
9STyTXKVMfmITbqNWdDx56A0aXUxNJ4yHLKSpi9jHBdaSvx1cSBHQQdSDSJct+Pp
KQ9XAHB2NYhFxsB88rIOIO3I6s1moRF++LYRlGEi2Ve50nSvQPq5L550FKljYpAU
JO3XnAo2S9EctSkxkol1a2n0L2EGkhzubU+7yLgMP7oqa3hZqNdmKQU+IZ1sGct8
rqjgoTJ9HQJWwb1qMKy3FYM3M9X4QANQx6JPNqylZ9/5DCZ8TtGQSN1+XGBjwAwc
rS4WVPXeUpVn8wVsSDEOoiLjCa+DhqmSSRvwossg+xYUxDXi3JQPb4xmN6wwwu3U
pgeyqAAlgDzeFrQqwwdQBYc6fM+d1GYfjt/ZVldAJb9cyM1Yier/NYHHWdE9idEY
DbkU/gEku1IOaew9/Lki2m+DJndLfHepnFXh8v13oicW5TyXxdDIAJDIbvI+9Ewz
Mp9p2v9fxejCHqTjccp0Wqwk9doWrtO/WqG6zOJqWJ/s+HEZV9po2n0KLPMeqyrA
A8wCx8TesYRgZON6qeOG7DVDmzmoFJhy0OPlqZYiYI3VHMSP9CnEbNMqA4+uMf/j
QFlzJrGZtb2Tk3fAOym/CvPw2JZu2xfANgueTHYrIaL66UZCRnUj/JBPxz/JRd2A
liyeM69YnXJy9RlRjtojJOZnPvB/BfpD4LcxY/nHV8GSiYciXNEgsMn8eQ3Ryb/G
Nfpix5H5qy0HKoKJfW0GHVgmuVMy9KO3dPvmxOB55hx7yc8RbuZbO4e/Id2FSojo
a2qcbJi5TXsTZwMFxbHpPFs+nFCDFhwu+IM7Xg2z3xz6ICHRrtDvRvb01+ooPmuQ
dUX/iVTir5I1Qw10PUe5ExXpNEQLSc/A3PrsZb/1qFUTS5Xtp73XJuKEROuvq1+I
NODysoe+DqiQ3ZOhTDSQsf1f3dMv/M2cTGuRtOf06b+3Oyl2ryp1Z3IHP4HR1WEK
FCno7LzaKSekDFa09hOwfb7ncRgDlLIcosM7XB8bc8niG4P1eAQyg/3LCt0RSGux
HtOCkqLvVJpMTCxGmDeQYBbfFrH34BM2L3WlrIqp5FW12JTEiE8aiu6znLorsIYG
LlUQHgpVse0KeJvQjvfrXFFBWRQko+h5/lEKiVZ19l7TENqrRn6MZyynzuTB2oOb
g9kNllFXenQZRZdKh/jzwb/zYcArNpUQsI/HN5pgZHwBMN79o3NvBBh2lH0JG3dL
o3ogSDcLVX2zSkkrJ3N/SahfTePW4vEFQqZR1YGeKquBCoWGwVeVUfL8WBKo2vGy
ZBwQTTsRYUhIJGc56K4usz6yhvv/Q21I/if2FO6clTxgm0m15lWFpXV1YPC761XS
yEY/n7udDAL56M82Frz5HpvTXVYWre1N/gY/zxQjR5V0qpvNin/0Q8JaD51WEBCa
Mtcf/kz7A8OS9H/9b4sOCGorfvJD0flTWOYgds3dyJiHTAjV3vCiyFLbolc2iwoB
nXMG9o5kFNeXFEm1TTiWaiBQiEgTaH+VfMtCbSPfF/1vWYmUpmJgcCTPluWOAmYg
YcGlQja6ovMZOuGvIpKghDWl/WjrVcgmwGnqTlDPIYJ5Gb+izVy23keMJB2/Ama8
toxOkI1X28p7rFR9i8KlS8CsmZY0IXH+VU8S6+9fwU2crZ195lwnoIZNbnMnpE3T
KdUq8BtmqfNxaslv0dG+DuUuSfvUfxxL5ILrCmgkoe7I0VsxmBrTlk+4Rvrkx+h4
D1p9XKKqdDuqHgMndthXeizopv15amsQKXiPQJhYJGlHqXS9BBUBVzj4N42X4GCk
QEwiHyVfwG5iACC9Ce97r/7RbByO1y+IQFWsvPbJJTeQtNPddSdLGBJthk4sJepp
nySohUEESF69aGBVx6U0hWMGwo84INU2YQlVwhfTik0yViiI9H5kUwtq5Yfqq0PQ
xrNfxysyI/AK3qkhZBA0lou8//LS2V5C+zadCTDW+/5mAha9jTF8jCQm+OWy8xxA
HzD7HQKjmb1CHbIdWVa0uUSMclTDHOoXeRCkskGK85++Ad+nzXJ0WgqCrG9bFgB5
HKGK7OfBFS/NGQ1mZXFiHutSJRKSsFt0AiFiCOqAGao8Z/uVDOS2MZVPsJDgwNXO
84EGCy1CudNdyyFbH/Z/urQhr5SZ0bUiUkuG6hwdXWowPFblepcp/UdPsETV6AH3
xYVJMevYbOFHJC+iVHZYsa6X5js4HJQhJwJ8cII88xd+y1FwLmam+BL304SEY/+D
V3/MK9C8b30sZTjBZD7sI04pNA706zDICcXhqp+gzMoiDyPtaS5uhWQN98dkHxYF
sj6h4yXeBA5LbZAJK1w0hRU0jGcYJru95MMEOb6Z3gZh+RQKbbJwrRZBExMSLapP
q1hZ24wktEocWXNcpaq2L4QVEgSiBGCX4PeB3+oUy2s697KOMaGh9F/9YInVhfTJ
sFdfC7uj3LFtJc0MZpS5SIOoUBbF22t0GeY2/N2GyFKBLDj+IamYIMcXxFJqwlEp
ZkYowNLoxE4hbUw+lf0nlwxP42vWnh+1eGvrA4EXXu/oGjLC+Fy0HYXTqsFsltt7
yLgetvziYT3kTCnl/KvxTiAZXHHb4Mr28NwyptSA7YynPkwglVMskNGrDx3N7fbA
ClrjaFxsZvbeBhaCIak1fzaF0fptOlQWV23wFdUTafa3SmOL6HniwjiBMeQANQqw
ojM0wmTDD0DbxduZ4jQPlb3A/FFwkLuea5dS0BHxdCA85L1v0Yk2V4BIF1g7e5cw
W/JcHex+NRNkUSNP25KKoCEx+89/Pw5s/3TLcVWxgJP2YOkvGFCDW3wLtJu0yATg
kGyR4vzGCdySO7eWJZaw09V6FUezp8Y95B4LQkfkBcAfBGKHsqq38P2VKkYMBdFo
Ep8Q2ul07os1MY/oQje9S5BX0uXH11LbwE3NzfUbz4R+3BT4odCTpEOlqFL7waLZ
M49qthP34JHFDt4ViaCYM13FnQhModpjzKgl/UIsnsRoJhCvgt2cegYHFhtoXSsI
F5S6CLN94ZtHwm4qVlKTYz9DxTV6yG8KBlwC5ePPEDUiNSuAeaqgM76unycvnBDt
b2zJLM3dSinWra6THKjX5F0H9yym5geZCCvWulobKimHznexEYZwTbOyUfWCtKMN
ik88A7jhQ2wwvnxNNLS2Fw==
`pragma protect end_protected
