// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QxYbF7NbrOWMvo74O8XlDzkSFZ63uUSnq+LHv8Ca1tFHWA7WoO2vNaTkbOwmdR33
Ta5Qve8yb7t8U3aCLagbAioJVbWwVaPa+xy4aBtUj9tRXvKRUnX2bBSRWPl9aRnO
6Mv1uc065oyk6JRrknqbsy2mkhv8YX/7WzjJCCQwKkA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9648)
8fqFgsI2Ct8cUng2SGp1NnfuSbNJnVyZvLUg4GvRWM4XjAn6fBhKdeXSQky/fhkX
xu0HFLGoJVhDbOIRLSfXM89XUrB10lk2xD6uJxGFAmf1HKbCywOc+JNH6zDUa7c+
/84f3RfF7pK99DR6/xDz0K2aVZRhG09PVFoZ76H4bPN9pYQ9J56+kgrxGLy0+f+G
r+YIghnlLll1NCNHXsvMRnaHEsky/PCOMIdsRJcZJVAyMO5GS6OjExLv9UunOVJa
o8BKsl5ZP3yCmQJI1+hiJKtpRIRBsEyBNmY7FFZ9tmV1f/JG+Zs1V9iR3QrH9aKL
PGI4fYVcIal4P5zD+kFeg3kJJCd/6/dU6nDtYmNeNpHqzzOxJPMtz7jHqskWB8Wr
bigPz/7UcXY0Sag4r9GYEj5FVoTfGVEOZFOYTy+c9by9RGrsqZzGupV4UAWtyhMp
+aT3i0uehMMC69TRIcWBSx2gFiLmewuvltxjHL1GYbRfCSAVgZ93iV2WNGKOobMy
MdfOc1L9wEvdTwkd+91F5MlYHn03l80Lnm29plbarWLoAu2Q80RK0J7xcti6G2aU
XrOuJXJBSmIn88F0MjK9sNu/BOrAzW+5t3uYOvtmavJH8xi44gHS0x92QUG92i4K
8pbCBmP5FtJfS1cpczoD1LqKeMuN2EuPYdyZHY+vuYBVLQBTWCrgSB5eMPWSkS77
+/P7l+MdDzuhm2XorPRXIBWt8djMXuPhZUmLU6qLPotg9fk0oDmCYfF0iZt5GOp1
LClDpBJcU8CKCTKGxw/uaVfLeAFRhJeov5gAplXKC9s2ogdaHVHpJB7pCzFLJSeZ
UWmEKntLc29FW8mTeJp0y8idjKOL9jhN8r0RqbQYny+7PWMszo/7XPWpyFoAQNiT
Jinuv1q5fYKqZ7NNmIkHoj3r1TZBmxRTxM/buKMvTFKldIBaf1chJy/v5dSqkcvM
rLZktczMT+Anyb9yzUL7J8dVhdrzd7HUHowEMCbHuv1LagowkBW0pKyn7ZhoeB60
UvtFaogu0pqWDioKIzE509wNUWijpWjI8inhED1YNDV/Lx12RLT4VogK0+/JL6Ni
qozlLRMxUFSMuRcmFg7BhP7HVXFyhKOU1TJyZPhiuQHuvR7QAmyaxy4OUPGplyqo
SgnMbOTfJzcLk09njUn3vxyGrmVKbNq2XEnTdr+ARAuGRsjwcWpGTQwBXdWcLM7G
knUUSXh5+M/A685i9CqWA/GRAMk0SX7GqvAcCdP/Qq2rggibvmJN9e0dq+khJMdJ
MGU0o3vswJZpEQaQADNyMoxgx8+HGIUPX0NEzAW11spcYjfpHSXKvsU0hwkNgTox
QtmhLAo6DU5WLVH9p+6AyMRpEbhl6MfgphxlKbDTlua/RIaCvEgTgzK0fyLG2/nY
IIk+gtOuBG63NS1dKkedZYtLSou/dszFCN5xj8XIo0lvp5GS7tTlHrIQRSUwkJxL
lnk3j4Z1TKvxR7Y3bKBT7utTP1V0K3OzPR2FU1YKqNtrHmc83+QxuRCSJsL2LZNe
0F4vSPDzD7kntyq/mKRS7crpObIi6xxVjCfTjaaYcCvrlOVZF9NRdiikYtpic0E6
bPyds1iNWhl/1N2aSOLdx9gVKXQq258l7eRvWLmbCK7An993AUIktRYIs4tMp+FB
v+bD6fpe07iMqd5PkbRg59wp8CDra4BV82ZtjsWlnBQzh9zM/VYVZGqckrlWr1rT
pn/6xfRDgkqJ8n44oJX/MoH7WLRNGMq51OsCtCX6eWKQI3wX5orbnQctyzvPW9Tj
q/DSyR9JPOsOSC7va03G0NjwIHBchxewa5YKMGE/XYptk+yoAGBYrwoqPi7dcR01
Fzlk3dhYKQ7ojA8x+sMXugFwYrWJkaySLnByLCo0wZRmDswlcZmHYQZpqXnCMFEJ
TNVuxv5vtUlDTpBoNkDNk+SxVZfDZwncd36Nihbhe0bF7aA+KEghg5KMcDYV1HWp
8+ZsJrtRRKEgNRV0zOw+t9ZkpJjFP6Vd9nBfqtI4KNlu2dAVGIOVMozmgnb3bv4w
lLY6BOTwf0mqEYGkxhFZ9H0dTpctAHqRuuCE/srXbt764SsDoFf+Q2CAJmaNWwKt
mGygSVhxwGE9BTchllWBxjMREHBbIUvl3Xu57gxlLeQIi5LavuIRBtc6FYri9wcc
k0HX6QcQuUENGLGLp8MkGNk8GJprCtZde1E18rXDGriTu4w3ujsJ1iv6W1KNVFTm
LIvnmRAEZrTNcPu9zX7EVCCxNtvBhXx2eCNKyf6FlSyhSW8m1u99THEcOwhNJKXP
suM8MD74Is9NQOoeda8WCLlje9VHVwmKTANk5I4iT0ywyaO0I6KzPfmPPy7hwUtP
+WEIzeG7jo7C6Bipnxvn4Kh/HQLqkrtcR2rG+rLOSJKZMN7sNPKEbVS8o9/6SASS
BmWjP9zN4GlQxs/m9neSwMS8Nu95pWb6kjWHux+YIVYvz6YA1g3GDwsu3/c+xaWc
pwxF48BGiWUBV3meLhMKNM1fGxsBVykt/geYYhtsW+YHUGuHJgaChq3R8VNcX1qT
UGhSRWA5xfK+bAG3+5f8vjZ417goyWidDyQ34OOHa7bLWiFZ5QwJnDxWXEjW25UM
FEpLm1cHkQEsTT6tlT6DBmE8N6ljCLpc+NHknHqOydGihGL2BR5Hw8k2B3LKOgsm
KT4s1/R9j0zY/9P3V3/fBoD3eDBrtW8sSkz4XopMZE70RS/WxXtSCyP6PbRtbOuc
fohJ5Pl4zJ8hvRuIIYD/qtMnbo9tvSD0Gis8I6KCQ4HODhWltKRilyq9RefSlH/h
HUd/vDpdyj+633maCPXL0VGjafzhrnp6UqiH8TfmlbSU5nrHg4pXOKZohn1UHA2Z
3cRTLfDYoJLlIHTYfyaeeahqAWzWGi0JT7UeAIXAIxN+/i+t38mV85I/sHNXHAn+
wHB97IXpiJW87BZKPUi8cMLFSFdgFrJpXkrD6/f48b9MTg3yVTfIJyC53LYSFB3K
jEDYXyPOg4Wbf8CySdUEFeCFtxg+NHJ4Q48qVm1DTNx5qha1C1Aks60RFX8Qk/IR
r7hbA2b5VH3Ev8C9ntC0eMOqJE4eqaUsrgiEELI3D+j6vrL9k7HT7pCqkiDUa3Xx
C7bzLJ7wtp67PwFq+WogOyNEpQujtc+7l6AqbQs6QyRAk84IaP48HRGW+pcopMPu
10q+/kVuCU7yy03HlKmhOFy3jfxUCMMuaVOJb62ON2VCFQ1R30CrGozd0bvduQsL
IKFcslzK+9r6qLroYNyxbTCu2pP1TF3ScILJ5KmlKbcgdQRz+VZuwJmFOJO2r3EO
xRNFa/RPbis/JEi5F7DKCf9iU8+E3kAbdFN3r7xak50sOGMmwnG4ki8tQd7Fus9W
3ObJf7PXIJVTuIFyuwCRp+CqLCAOb+/x61FL+wCuvqU2phH+dx1VJlogXt9hddBO
99qWCiRzxZKFpj3vAFdzK37LGTi5Vx1N9ke68VXdm2nYhpo6UXMh1ZNiG5xnaEmA
Tqcz3B4Dhvc9fBqj6FjlP8tS3jXy2pvZ7MYihRhDzQDaBIGrfoIBtnKcLT0871Mv
FwbLy4HE6esvFG5ZLJ6sF4/wDL8hfLDRtDzk8iGtB2H9bZdU7qvvGxv4BMUcdYUF
vmTo5EUcUaGZqThGBt9uhDnR8pkx6HbbJMQds3qoXcalEJeTfu7xGlKb34kNIn3t
2cDEqY1Z+3JgW5hH3rLjFql+UMa3TODUulymjKQOD7HcGEO7mAPnMvOPC42doh1q
vNHNr0o3ZzytnvyISZpAJLuHKUA8I5A5RLC0iufboQU5GM54O1LDxE+Njp3tpPRB
yoYD78GWnZndusZ8V8OvAL2PtHI4UapAs6LuFy81ze2OmF/80lQS4fI7CsSOty1c
nQCHURUHcZ+Su8SZAfHarONMlD6gGFPz/lejet+J7MGWp9YnAxhM14mymF8hpgZX
XTmxPKCkM+FVhvrZ1knaaZeAXZTZ2Ay2EtCJV+QsYMQ3yu1Ui+SfYvMtOsgZTezd
rNCrClTx2zV4klk/oCYOhX2eWmBw2tvddnR2SDX3XtEFxJVRVe1yQGeEN9ybyfi4
2R369p+UH7Kdm44I/MESjwFw5ocVMEBhMo6zmcCwF5DImK+qzzMVHFpLLtLBqtfh
lmgZR1uF7Ps4Wyeyaorc8k91GZHIY7fbVUpWdoSM8d5ldMemJmlrvmWUdXhASXTy
kD661yLMiBbK5J2BTF/h1kw/1xszqsxQQyVFxSWgxdhdGVxnb9UC8fvpivLOqLJv
vGzXpNQr1WqjFfgbFDgKsGgJ+1M5vSSJRfxeECWUTYLaSE6oBPakC+VTaWaenR4U
fFGwjwzOgffyIEJryvbJQQvyWeVx7SszrgxZMUThBx7yFJN3DgpjkVtYmRaIZ+05
5UwdFW3VfmWXPR8E1ZcWr7cUJs1dMoWwTnouZmsMWYWW/mgvx+HaPhJAn/2EEca9
9yXgErJUg8klkoUAKHqqoqvJG1KsAqKh2p2DEU/He4R1bO0Y10fYdQvbwXXdJSfZ
gGHmOGj3NiJW+XInIVhf07C/yguK2tlJ7sibimgTSKGAiVpxvkpxEjtezHWcJjkF
NIXsSQl25fZeoqhFWPX+BHbtAZuZ+I1X05FfRFUGfHNOnr6BapgRU4O6Lv91OV6n
rT23sZCp7H2HlYkJSK9NtHY0xx4AmFiq6+EGmnbEobDk0Ttrip07kaCC6Ibl4KiI
Ta1KmyIhGd5GDO52+UGmJ/q6QdCVCQ82rgRz908Wzr6ozIebwanCnECsrBesCP9d
NHk4Sv+87XoKKUAZTRSi8/A6OP674VFj+HY5UenrcyDi3Pz+XjsLcpAvKRHplc3V
IQ0iXi2cwwslsxQoeW5xpZmJyMTYmXkmTiFHrXZ5iP70CqpPefrDo2CK67kxbf3A
mxBlYgRjGtaNuX8QniV7ffu8c+R/Rnpq3D3atufc9CJ5cYhKleIxAsaM4paWWUa9
+b9MQb5ZBK+biRJs9WZnPMpviX+1906vdUa/dyIJcCAsqJGBnGGqe9gtyYSedP4t
9WS1vs1DkE72axJNLG19uY0frmb5phaMGR1qIs4yKflV3v96Ba9xuoGFUd6W78ua
ermXUAwLbGJavBWw4BWkU3mvFySblvM957e6PjKUs1YQhmJSj3mt00pqVWj9JFNk
zX9Aj+Fo/FCpLrGGOdNPMZlSmp8eO9+4eV3j8EVX8omHdp34XDm5V1P5dd4lAL/7
/P85ej8FRRUK6ZEq79kEQZfNn3dSVRMBjS+5oygRNZW+b5YlT94dfh/bTY5LWROD
J5iGRuBeVWRpksvf6GvYQ6YUr/fBZACfWSINbjCGP3GMKNLfZwJ8qN5zsG3VWe/N
wjWjz066XGEfWEXUplE78GNZzCUBZrxFDxFvrumWrDSepLRj+feeJnKD6Gadp3cu
1xzX3p6pt11yqif7QMoVFlg0+BQAjiy0mHCrJ3cxPlUXn9YmUfn1L/TZdPNwRWwd
YDJ7p+NVALhPpWCM2XV5z/s3/r2ThYCWhmyYxILrMRbP5E32W+/JcXDCQmb+khAT
TIhhUN5eK1CCeIGI0S8FCL3J0fNEJpJaSlmZdbImBSoNTNHZO5Blhiw3QNiJKM+z
1v2JrFuoNeiAUpHK/3ej7jc9mXEAcCqmMEPefEL2r4Y+9aKphPRGZMarpGaGeeOY
+/5phIE4vz7qPSTCOEc+vR7Zfqv1vJ5Y9zmhN7A2QdNr+FWR59OdAYXROTScPqZt
EKUnqBXMVaLBzc8QfsHj8Dr6NgWnzRFCYLMfo2/XKzrht8bkzVKOiBm0Vlp+Ra9N
u+L1sKfShLE9fwAz+T0LYS/sx54ui7nf087zZm55b8XuKpZRzlGc1hDTxilvF/KD
0/sCEqxT23SvLRhJ3HusUSFHr07Dz55cyd5pWBleh/pn6mOYMPwPRO76hT5lCq+s
KPxk+Xx2txjwT8iOeTGQN9ryeXOawOxoXbJEu4t4D6VwVMV2uyWCdYWlQGnQZnN1
ODI5sN65KGwBadBja4HLm6yVMYjkbKNNT0tuiA0AX6ybL5N1iBKmPczzPQw7ZQQ9
i+xeyKaDKs4UB4XD3Qkd24thEXO7pwq5bcz5VM92mX/oAKO//xGx/IUvaL9gTVTe
HGXIuK11qNiN88Rg5Ypq2SpstwpM+M4KQpp3rAMNti509fZVhxo0yw8rL22+13FK
VoKliuBA2K2ygN9Vg87pS5novSbGJTQPt21heNXVaF/EytiecXJT1mqgU3qG74UP
MiCkArZIoRXC2u60i9Y/DFdzwvg+DBmANXc8HpxJFZ8ZDsZMyV7z2UoWCur/AAYP
5HrOZnZt0x3BTuYWlzWsfYHQYmOiPOgLp8TBcPDMaXJcuVcLvSx7M6eZxPCjtVZd
utbrFJx/ik1FXYYjAI/yl42VMbn44bkPjq4KnVk+EdsB3tRxwa1niQ+7ltnmzYo9
audYSx+b1pHF5hkRd9pRoyQ5IMAjsH3jYY0KiMH/WpHSwLb0Qb5lgn0uf0x686hD
gh79RjRWPKpCeMuOUXAzYpAihrhFxeZajjaJouM1q5g8nrnrSfjhXsrOOQ/FmU9q
I9mwqeoOE996QJ5LImvkyw4zfvrlGJXPwmk+/Cy+YDg89Om+h4a9Msd7pfUwjdLE
zG9QEdHWtMKudBwGH7eQR4BfI0mVGzrx+FW3SVlki3TvpYIUogTQUcPqp1kFn0Vr
eUCcPcLn9KXr+dPr/Sn8RiAH383ZaG+T22m15h7AJ+AeCom+Y4XsGO+GawAwkSL8
9CUvyZ2sN/3cJPjP/OhLdrl8oF0QeEggy/DEeUG10MHnPbsnhcSFBJnXwkC1eJWt
Q36ZQbhAps0sSWjGk9seMfzGDTR5UeCL8Ae518ihys3oABP1QGBAh2J/hLdQD3A6
iQ16STTPoCPpPeTfLcvPqGnuh+jF+YMugfKgbsrplwZhp1g8qQjbJa2A2/LdPmgV
YM32iwXpg0y/l8aw3CQDixzYyqokzwpoo8cBlBCMK5Q/TXv6s+c4E//ApDDJ/fHA
Mekg9SED8K49N6a+GU2N8rs8y0WdqcSjl8SAvPz4NJiv90I7uwc54eJQWguCwXJZ
YeLrYcMTB6vs6i9HR+lZnawE55+UUapzxcLW7Rxjwq4Yd6FCyNEJeom/EGpg3Zm+
rnKnacRmHxnwmzgKQbhJ6B34RX0GMXRKDdYSc/Mk9i2CHC+Wnwg46kSE1WUDWRvS
HkYJ6T+dw66atU/GJcBxZswJAT55NV6OcTVJzpb4F75bRifqatjWc47ygeZQIppr
i45oe+Wv3VDrhqfJLhExurOlqZ1kxK6WyVj3t7FNf+UzfMCviUiMBShSafThSTvC
CQPQR7JH7OfObSCgL6W4C0XFlcdDSeBHmsWpFqUY7lT4iPLx4KhL8SaLeIiOR0Mm
03IAOMk8SXL6yjmieF9Oq0aO2ZBge1pM6LiqQ+0Ni2qlQIBskyDzAOVsBDDalCrt
jnirJptN8Qk4v5LxK4PJt8Q/x6uPC6QT4YcKQLqa+8d4c9xd4PTW+ic9Ay0ZlhKx
RVBTInpybhpI2WYIhy1GQ2Mx9fBH7hNz02NW8uaTJ8uH8pWO5btzvmIhfM+1u9jB
iQIGB3s2pFwirSmjouy9mi6KwT0tut1LMQm0NbqvNAuFyeEvyaeRyAZ4rkI+yfR1
t9m44/cfQ3JfVvdcOoAxYUsNHJhBXial8HBD+XduVUq+uVpbmeUFpJCgJJO3MdXj
BRq/1fYc7qiJAfFm4hQUb70hYEvk6f4HYzGY3F8osfZT3BH9Umxr0/SnDPK/zmYA
RV75yMgiAQ7tm/L4w3m6G8EZNiYpVcrwt9lkCUf4B+M5ZnxPuOZmz+neyBv8LCdu
sh/OUqMoyr7vWBmSo1V4JDV4M85rFpp+1gbzfT3m9I+fCYxeIY5XX5mFaQdMCNpc
phzyV5SkAl2j+FzqqSamWANQbjM2T8R6g2QmwdSJI9zU96+brBDc812PJcDtk3Tm
zj11oo8kidutXr/rl7CzlTRB+V3EMTiPTPMTXS7hK7f/Hsi4d0bP9RgUj76V+/da
RLGWsZfmHiiJnjS7S9IhOSAPsJ0jv1YypzGesLZ6tDOF+X0g0yo7W0a3+eazveKR
x5oOAnUweaM9KSSlG3XlrLSHTy9qRGYyKRT5jWhrPY+C2kzXkDqpvVPZwFSdxtL9
UA6brEa9SIE7fWOxEzTjJHkp4UFJ+qrGy+gNexCzJXs2sHteS2b427hvUSRiF4Lk
ol0AWLv2YoVyVEBMj0yGoiW+8Yx/90r3tJlfLgHIVj8+BkR4+wB/HtHYwtYiVZY7
YXYA+jdDy0UrZk9y972pGiuyEHEp9moZmGHS4Y5dAc2yyP9uwOKY8GSSk2oD7oWR
urN4I9PEtMlkiBYC3vKUy643PxegAVYV45CtwDM58seIj3sn3cYHaU5f9910bv22
XkCqeiPD70DLAev24is9suuXUWi7IdIOc5XCG6elKB19liHDGVDY+gZrZJ4SC1SZ
Q4WZ6AkqRrZazXcgHeF2UPnMMhyR7gw8/xKwkF2QZZw87cd4qpCSA92O+lpfCnUJ
jbiqWEZmXt/2IEBYug0eELJBpfT2UnTuKPDW7UWyFkzA2ZjDDi0aUx+yzNcB+iMW
47B9a82FLq6jt4xsQm6jm+jsTjj6myMMJl2/urE56cK7pHyREpG7qIGLvizkUHaP
Hnz4zV7nS4YUTnh5m7Sc0DIn+uNwe4+Dh+FkVuxzPip73D1MZYEoeVZZWjq2N+4g
fcbMyaYLxOyx1/LSi6XyX9zv4DpH4+Ve0UA8Uv9C8kfe4vYDTN5/1r7OWrg7nLX5
2uGxXhOBQYcSdC9eCB6F0uETvbBTNb0BRKvCXxQL2lGNwFYWquKk29mVWTGLuxNg
TYWSaS4k3aQbDyPyjOgogoc4hQU96G5lK6pLn1guqG1kcwnj26rCi/nPQUp1Nvxx
NHR44Q2s+28OtPguPRygcqwTFKry0dm9eVx16vcH4RT7iEvZVv/K8UNJSpkKxPHJ
9XMSK5gjKOxX4xyaJ7X9zJu4MCH6v3VL1OB7F3cv/9P2NmlqxqyA2rT0XFJwgGey
9EsrLA5Iqbs04pG0YCa2bgOqRklyb/IYT0QLarFymx5//f/Do8b/Bnm+N4B/Ii6T
G7ChXuCOihXustfwtyhs47Ae+88rX3FixIIKOZyT8RXWTN6gIMctNPRGrAF7qgkf
QZotuEwilBay1q0zRlCPoBykSPn7i/+6QmDNQI1JFjAhS9TSD5Nkp3Nzydzi/UWp
iyYejZcUOdyJYVBaP3b70T1IPR74ogVj401vg2iq8S7slhS3EFtLJA04nNSgWGGW
pWZJbVU9ZbZIav+RbbWR3y3qN/tGBCWdh9QNyqNGRbFv0gr8Fww9hP0XjaRx800U
/4koZTfEul+3+MnUxed1MEw2qXZZ2OPXIMdybf60W1npcjtqoH8WNN5s3tNNHSx9
3cqRF9nAHrD7JX1PGxbLnuW2Xl47CN/CK1JdVsOvTS//TWmJwI7a4lAiGqJqmel7
5LD7bSC9qXHpQ5Ca8UT73IdEaZlJE5YkTCLSwEtZW8K8YJQ/j/QHDUZ0omtw1+7c
BVu9czRk2D/1ztPOJIvhfnV0Sz9H/FfwtZCxS/fpcCU9xE4rOMXMs5byQowggoTn
OspnRgE7CNEIuS+byuZg9is5XdcMQ8YA2axqcGan+SLtK/0b1xFDoP7iMhh+pfGX
FkIL/AIgjOen4Btr5YE1qXipUujEaVK1pbw7cToiLpDZeRRVTU/tLl7pOSYoK9p4
ckJt4oDG+zTdagTquKE0OwbKulVR6pv/SLSLUOtRZ92vKqvxXRY2VTKdUlxwSZvt
QGxGPtZ6FEXoGPXMqNgHxc8eCfkG+yQusrFBKks2pXTCIIM4Qkfe/RO5icgKJi2w
RgvU9NzR/TMa8JhOUa7WuDkQy9feCCXXCvo7w28hgzgGLyG04kpEubf7CpPjHeZl
ba5tiM81g2GA+q9c45eg+a+3sF0ZhOKp0rRId15M2aQTX6X9V1l5N/Ig94UJ3lie
K/iatZHeF/yYmYa7LCN8CpqGnFeWyBM6BSS8P+ocMWIR9b+hBfq8IbScpLOzX7el
g0FpbmzG1s7/YBD/PUBw91SG99qftKQDBagFsoh5gGSXplFk9y4VWj/80Wv50Doa
NKJ3L69lhzWKhl8AlKUPZq3cnaEIraXH/xMOpA4niI8Xho4eCeSUHYvUM1lgEdhM
/a8XduET2lelyZoAQfvpEYbLyuBsuUYQ8I7QAGLQfxMBBXi0uHJ4G5V6Hu/nVV5w
12ygu4+hk13FE0McwW07mbH6EbSEfLCyuyGNNHmU26OjsX/Vz0en2NZZFm3nAm/+
1pDPISfXBCkjpn/lpo8KSRTvx0rKykOTYQsZ6cP8RCiP1i25yTifG8ItdGOevH6B
ZJOWn/kSGLJl8z9BFppEQYcc3M5aAVcthAYVoWMeGUEghB6/PiJ/0xL42V9FpmvF
epxyW6YNpVH5tNX3+/S83TwqN13ZdGrOdvIOW0MQthro42Y9tINeEV8QASj5bVlF
VppNpaOwFqoqDh/HQTeY1QmnEvHeEC8XASiSf2emx5cqqN4jZHd1pPxZ57nj3T/L
nZHFy9R0EZXE2DucSWbR1FSUe72iIL09P4OxkUeEo6DWLMRL5MLwjBag8M7Sb5ky
oDrCZVC1Pm2L1hd9Ff6JgfdD5sxvlesPjHlhyIvU30RgVtC3DicDTLL7Oyg8wdBJ
JT1Mpgak4CQ0wXP/Ye0AYDaFr/NbxP7WfAaQfoj46NnXGsz2d0LvAvHshlg5wm11
H2ZxpTtiaHO8WivDarpijb3/B1Kaegvjv0Z2NQK3bygOCGIjkCT+kP006JTQBX+g
9GwpyPiY/YTnXqPQC9DTmJ3nmk7OsHvxHh766i1Q1WbuSZGmte6BondGCpjBqHyk
FRvXqW8GJO/pfWnZ86xwr5rcP2Osj27EIJr/GcqmQrJx3/sUGL+Jr/2x0wIXTTM/
FL3VSO9En8D8VtbwvX/Eig6t7cg01BzCmnOfDa/xlzHthpGceFw7o47DX//NvyV+
p1Ym7wPM7vHo0xo2EBooZq5K5LjBAW+zCfRMDukimXL8gVnBO99eu7wv7lx2mVg2
hduwuefISAxaLTa7GW2WduIjJLnGQm4XoiEGHv++mxocVfWPoY1kAkvidhcZe3dp
D7KbCIRp7OMsN32xEb7pkuLqjQWXeDl9b5SS63zFPKXBq/HeoUmPJrWQInN8dFqg
iW06L1+Vr1jQG8wQXl9zAJlFyKzWKXMPIj9THBa2kXuuTlKOkmlz1u14jD6pbVtF
OIlBaHjNrYk8t8gdD0XLV6PHGLR9XyYDK6ofIeNzPx2cNUdZciL5NcltJLDq8UHw
wKQz/Ehh5dxa4ait6AmHzQS6OT1yqDGqT80L8fT/03P8059QOUdHQqC54udxfEsG
UaBemNvWSolZex7mCjUmO3y4MutemMLh0WosOMVsSjLITX6l3qnEu3v2ryg6bKuD
+YOdFdKhIUv8FvoA/ZqZ8Hlt1FhftUDyNxoZGTDT3VKa2Ov1fBGgMVo+9qVugmAT
vQLOkL/KrGZczzAss1Z5VxUSRMna8CkT+RPBp5Wqs5y+LJx/jZGXigf8+i8Gc8GM
hDvlQaauUeKyu4FZ/9EAAJlmI4ntQQZAg3k3BJ0CGCsqpn8a4KttnkYAdO1J1kdR
sxAYTVEtp+qf/RX+g1GovlmvuMXorzPa9+BmyEvkiiKWZ7CmcVxTjdKXBILmVpQG
lNSZb6hyasCnrr28NscxRAuoDeleW4/KuDwZe4dq0Qr9Kc1hWdN9fDChXX5hSDWO
nWBo/E9nq4aVE4ZDRq7WlmgjeF55Y4BU3m2thtbTNuiEWuB7hP/Z6XMqllAYqhpR
uIp2+bqkGny+nB2PvEa30aoPNa+tbhCeSUSnXkaUIUrjmZjJmsGcQsfLynO4YNfE
qA6lbM4Ki/Egxk7CafM2pMJbMBX2lTxYvo0lmAkoNYsR63XTJMtwR6Z2RZr/WO+w
xU/NqTKdojxqwgNGQI5lEWfv4rcpClJc8KiHXMeMd0gkzZy+4FFNrssrGlkcLqK1
8ieXvvtp87UmT7MrKfrKaVl78fi57GMbUFjnUhDlQRW2wmmqxoEcGnoFyQ+bM46q
DqKGvjy8Gf5D58Q8x8VdQ/DPsuDNPI+/gPIpbgjY/NiZxhKaDpdzCA9RLPRcqg8N
wtM5eTLkF77HUhC6HG/mN/qF/n0EiqZtgB2jEsLSrb0nHyK3SUV4hyrruor1lxY/
IpdFues3sht3WrhAX7avz8cZgRBmiGO7SasTkVyetXVpEMTxHx9NTvwqB2t/rQ47
B5sisjF9xhWqogjFsFe/XfbXoEHc5Cr0A5rCuwLzG+lE0S+h2wPYOALbseTnILlY
2F2WQbfqxKMqZoFFV2kXumb3ncepymlfaoekPpg923qIHV1SIyaYCEnvbO4mstSV
tH43zj+p9DtzPvu5uqD3tZ1twwZYTyZ2I8AmJWaknH0VvqHMYQyd6uud3Bj1BvOa
lnXWbsvCb34pEHFWJrL0khSPNnuMda/DPb4HxVQv/VrThJ5AA7Fa8kn1grEGWpgA
CIaEc1YLpdVSk0cPpbWSbaTd1o27YTYYT4Njvmngh5lCYnekPHwMghABHntkAeuM
0Gr4nFe/EMUqEiX52BeNZVsQOVHhK29xPUFirBXzUnqGsW//29zU6XMPN9Pxvj6u
Ruj5PFk8H7STmrEZTmmqjeF/71Uv8SrcMdpqYQAzsQoVd+Vz0CO1CQhzVpVTZai1
FtUWFqczUjWMbWuHJouBcnuCjm6WKStQ/vcBW0XoWxaLI4Ojla1C263QjGN6vua4
`pragma protect end_protected
