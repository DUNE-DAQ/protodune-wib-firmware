// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JhSxNBt/mlFRML2KPuEpdGVmO+uwQ5+5ppelDrWDyuXsWvyWj+s0vbIqFk5CoBdb
JFNUQ+TyqvsvpyDNCHmFRL2p1RLJg13UG9KY2H2iXYirJBLc18TkW//ET8Yit91G
5nH4gcOhtZ58u9mD5CNwZ04xrtaE1kL4weys7lGSkQ8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
b6gBRtbwKZRLCysNrySGNsKGaeDTmqC/Ao3deezURaF/FwjtdxkDiHVIuI5qJcM/
p12A53Weenwkgq1VrN32yOiZMZ9gnEYSpzJnG55kgmbYR528rPyiiKvkhJYmSxaI
9MM00JE+pEAetNZZ5/rb4VpNwtdkfqQ4gDCWv7uXJCJXpopXNIHLlQJPNSHiFNgi
SrTQUMZtEGEzN2PlQcA5vIRLmDPhllwW6DYOJGVsJ2FnLu3ZORkIkuWDFRfI52QP
LuZwS0GeqbZDe95I5dked3XBRWoh032G/m2hR2SIOWlOYNrM8zhwMVNj8P53V7a2
6pFtYiYJnA4PeNy3THMWnLc+ElgZDTcVSjUblrZHCyiZBwH140xgdMXB9GqccExv
2Qu1FfH9bOZTFOZPLRVTB2al4eYJLx7K+YWc51W8vCRweEyfE2uL1ZbDBfx3BdlU
Tdnjbpr4wGl6gMtWpDpuxZ3KLvtkwD7tYB2/jsOlEQvxZrdsWldnqa2VvFEhUeF+
4u3oMk3FUOhF/Sbvb9qMYPQBFTacniVyEUBquFLWDq7DXQRAPsEtl2pvleB3rH2d
xaJQH7IvxMb2La0H1VJV+W9jYitVA6DqcO4qgOOMAVF4PeDJO2RPVWK0NhPkhEcM
gPju7ysZU0YkUnUCO/nxGUnKyT+pxz5J6NmgUpehNhrt7tr4iohNy7MJnH5HKmdl
08L7HZLp6VulAMY/5JRlP92Cu00LBzuihJxACZPW2LAEjyvGB34VYPpygnFxPM68
PhqSdoxc5U2RdH3d408ksGmZSBS3U2i+SKY0XOrkGl0YmJYOhHO2EA+YP3SuBdsy
AMj+G1rp+OVRj7nB9RdMIyRULRhFFlESVKBfdVrTllArBD0nEvMXrXPA7/nCq/82
+hG1l9SxmtAB4dGRfefzYEJz/I0FcKVrTXTwywqsvs0xnhMz5NzcP7aPmDe/LIzx
vIdrOSzw4RRvqq7NqoLDdK42L3Z+7lnNikivtSnmLJVyrR0kx94HLtOA2lK5mjAc
23EvFPew3W5ZSSDSKDITXBxg1RpM3iKyoIwqUmHPMA9t0fm8DtSGVAiXX+SV8yEz
qDej5UKu6Jki1+GamBmiFsDHd1Ze2vnthVAi0mUeFecNyvi1pAPwHqrCW/hBEu8K
1JQIhFNFtsGWK1z0tPUE0JlqiryhbAp0s/NFDq4X+dkkcpFuoPewWeeASlNF7ZeV
EXAQKW8xfDmskZAixMu71Xb1RABS9+frIZf18qyZDSVx/PIqw96098lxxvH/kRCt
1nIEqljowHJoOlUXTAlYds10X5g2OJWJ3l3Fef3WUKW8+2ZkQsNLFaebyzKPkgPd
DQa0qKJNFm+8wn67W9x7yfr1KEn++al4EoZYCdqzfIbjx6ITFuzPYR6qJx/KCtUC
CxD3yT04JDbN6aqwQvZOFhbQ8wjxLPoET9Of+aobw4E0VLRK55+1FAsdkTK2x6u4
T/VHndv1zJa1H22vvIDuuuhEFZadG0DeACZcSekiknKoShj3gCSQnh+Mp7mMJ/v7
M4Guvch0yQ+sOdfRBjBhF94Vj0I7BOML7O6ABkJ89HVKT3jI8GEA/nWR/Cs/yZCm
ZJqHqJkPENL2b7Qa8QVLSJQSF0OZSROKs4EzEJ1LjiH3x9kHxb6Iv2/lHiXWJ1A6
RHULajb6XPauV6JM/wZ4Ev9/oEbyRKlqT7ORrWyR6dna/Xp/MnaehkKFt8KrGSoq
sFoOwgkbavFaMLpD5j8SCMXq5WC7A+Wnyc5J9kljmRdr1VK/EEExd8hbG5h+GVX/
9PlEbeBuWznwbvxAbVZsgExBEuLKv5ueTTdeRq6oV0HhZNmDNrySHt+/ZQbdedpW
prI9N/tYNovkRDIz7+aAfEBBjJ0udwm7gftCyHTZxCdZcHb0Nbh5gZ4vodsQ6Qvr
SbPqAaqKbcPZVfPUIeV8mRrsyAQTGXT3voq015oEFPBRx4Iw2wsWwtujIDjDJ90a
Oq0BkC8FE/V8WSplFoZnNcBSFPfNvqtduRjMAFCX3hKWzU2xAcUbP4xCbANrMt1M
hQimeF5tSXIyzdrLbAfbpDAt+AzIhnUsFDD14+dRopikuyO3KjXP6tmBAtak5O/4
5ewio703ThbTQ5hIL5880m0FdJFbTX9P1+92U+dE8VT+oti3SQinCT35ME8sRKSc
6JvSm4HrtKqakj7tSkjVt35Tv+E1nUrUZC+Ql43m6Yz1iDUDXUAGald1Bsk3UV3M
LhmovqB722G0mGceFpiXQzOUMT6CW5NSQXAWS0TGm0wyiiw2B6MaaoPNshWecKoM
Ec69UflYqhhFaGR58l6j+OVzdsLtMAgSMkPswo89g5pX5awMEhbvgawG7oRsSazG
44JLLeDWxwlBWZg3AxP0vsuev3iYKPyHeh/Pu7QAw3kbKzM2HaG2MHT1K891qt+l
EzeEQzd7ZSLfGrozz/MpPgegM8x1nvZxQ2Xh9CLH21EnCgH1Km2BXDD0zN74PfCb
f2Tr0FHqhru77G1KZlUM3t75eAljVCg3wSVvnPNoQSIJVkPFbhKRpYW+JFT5papS
tmCRzz+oue8wSi6mHZWh7Y73DnbcDI9qvqSRbquYVXbyXs27MV6ZzYaxI1i4DCsZ
wgmWdFKSgg3CnAnOMu9oepr2m9e1t7U+YI6VRTb/KF5YNpLzLzoN1mMRNrnLXLpk
rvhkCDhowZ60SnwiytakBmpBpxVZ+ZadyzCohCXwsg63MpBZdDUk4ULGUPhz4Kra
Y4r9exvRXfsXMK2a0gRPh5dV3rSSPfV4pkGlRWR9mzI4BG7L7HIl7yNYCbj7uAZy
gV73B4H10VOgYt4EGrIIr2AGrrA4A382s9ektmrNs62X745ZdIYuzyp+v9LgF8tP
haJpT57syXMmaxmJeh/+vO93xH/jXLY4GApaVfTcfWNHZptMGR/WPiLz9xoc8byr
QBtkShUsIkLVmd0v/DzeC8mfIn5F3nyN6mcLmfvq+3SOziMAxv4dSltvHFOdfi/q
W0qsgTNXZDHcTkRXu+F+lh27hODH4rBbrmRZeD18+odresux9egBE68lm3HgQGX8
yMGbw4DxzhIjcsfDvCd1l/+JsxsVWw+AhMTmFI+6JQDV7W33p/aQtmIE+H4GrF31
hQndRcJkv2j328xum7rXCVcaXcTxACrYcp2kCcQUtKdU+4AyIbcqXQbo8bBnDIl5
RGqAtNYaKX1eKMK94HZj3gZ0E+5wcGCITZNHOCxsED7URZ0vVZ3CNI+oMkbAiF14
26OkmmX4qE0mvMUYXjmUO4609F654twZRqFUw7QxJ+s/ERnkL0qx9LSFXe3gIEaY
44OfBZb+L3VPtwVvcKoBBtLi5abvLdu7KmzfOFF7eKWfLw9QXbcBCEG0zeHp3gTw
+q/JyVgv6biUuf5hoYzhxrzQLnvBVa7K/ezEN8Lk81msHCsrBdQ+AWibi4naBIFU
WFfpPiTGiuglC9Kb2bbjr78cUebDICM0RIk1FB/5Y9H1jhmJGJei601AkXHTy0u4
DtAs9gJ0Ef6bs+664EHOKwQPPUs5jwb7x96dwjnSZFeBaV/28UlQO2E1PzfhJZuO
SX9gejpJ01/vqPc0gJgUrwHlkXogyNz5JR34RE7YRC4BszbyhjrRfexT83KKJpab
6axRHlw1JW2st0kcpS5Z33zNta4Lp2vu1KTdO/lkSCTaJnl5GOZApFSMl7uV94aD
9p7mXPOJKlMNjsaXOVL4xR0v6er+1aBY3WOxxCORpWMH8YgRtdik4q3d7gaFp6bL
MEKqIDvmvOnpeaSOL3vFMgEzHe2i9A+x89JJ3jz9ZkgmWwjTTFL6bTOTxROwuJ01
8r/XhrLOL+FfR+K/arOQBs6kz6MibgAGZzhS6la7n512BJGPPz10iMSRO0R40wA5
GoIwJqB+6OVgzMeZnlvK+/hAtv9G7osFEWp7HWM/T0B/LKGEYKwoL5kw8Iq9ytJQ
bOZU1uGQ+nZfEgj1ASreak/2mDFFULEzMbFgPZqULeFpMqYMSgrIEJ67s6kqX2Qk
MlkkHN/NQf1IwoNIqYy/xqZrJhK7E/lJuaGbGNlX3nr2cz0VPm4G1cfxozs/9oa9
33lyTHzEyh9z9apFd9n5qyb/rPqyHg/RL07qmtjGqoNGaovhMcD2yrGZFOFO+L6B
wvNCe2gi9lM76Jl9qlo9b97P6Qa69m+HQwYMd+/kaOru6TszZ/WjzxQS7CbEg3F8
NAtzK8poygs4aJnAQsVn+e9hvTKEj7dxDhk9pkQXy63QDkLYi8Y4K4sdP6LuQFsZ
wPbzC0ft0UnpeKeopkGa+j76WvpGToqZM2jgt9zyd6gl9GdArOKqxqcEfcldA1l2
Lut5ou82j+yQmqMdcsOUTdRTQVF9Zo2mC3J32RzKTFXo1lZAMjHIXcYAa1vFSrG+
I/cTVEhZNEOADSSazhNigVZkIoiMdEh9EUb7XQFoLOD52BmZK+44XnhJ8mbsmDqf
k0UNxSAQKoRXcHC9xizdllFiYcND6Eabgh4ap60Y8eNY8rJI6gZ99M+jUY95ESKv
AYiz8yXiwtFlRG+4DVzbtbb8rLI7l6A33/5ZGOKFNpGVpPlldSzOKj1S+aglDHe3
Q7Fagwh7F5j9d7ByRHvKMs1Sj2uahiKvGApHAukeb1faFetA3J9c1R7+vx8LZOET
kfQGoTY/o6xvqVLowwQ4dUVznrrSR20CRBnBlOMyrToGekK4Qdbfebo3tLHokRr+
uA5XhryhBoTYw4ZARh2upKHczso3o6/OlVr4f9dbzLp76Fy3ld9WEBaMAchrgVWL
Kvk3Mf3vUMf9yX90XUK8K0i/AlUiBnzpaYrASHPdx9CGynJdUEbpwC9RDQSkHL0q
vnp7tU/F3Kq74LK9Kj4I8v4J2LbaUbaeoGpDMjHhUaRUu4/1Sl734qPKYdU5GjdI
hKVLyrWN/z1a+dz2uiXONzrSaXGMnWDo7FfQ/M/a98fmotRKbgYPHQqJQSLLHe0v
o/nXyjqOAWWUgPKF3shVHoiUtHkTPea9qArzbfgKEGJIQEEkCsPiPyvYGZ7Ir5FK
hpIBvfzvGKz+i1zv4+ImkUx25O+PotHsx0ueUUEXELAZ9BplT3eRMso1SH9HFCPR
em+Zdw+7fWgTuO9T7iuOo8J7SUdnNHrXnOLqA8rJDV3Isv4EwLknhLedCrqq2+Qh
RIJbUbvESZP0lSJxw0XIjU3dX9s5sYAaSLaI5smRBnepTD2CVsMwee8E0BVDju/L
e8jMibzJ4bgzEHbzSnoMk4zDrA3kDrZ8XOspl3YBsZgkalF9wSRtO24oequY7urI
Vs77OspOviVxKoNU3piDt7mcwVrhs3OZThkCEayvpYo3Vc5D7CE6dNy5h0iOnkZ1
CA9Io7ixsR/8hYMC+DGJVRXpSClQe8+VOgSaILOAufCJdm/zAGXbAYnfhtZa397V
WaL3Y24ZEuk0jmX+1KOikJLYbsSgl6Rit6jfSqYBPQeQ1Dj3cHXkEUTXiJp+U+D5
omDETAd44b1PZvkNUSGTeV/Kdx1idw+Amfn/7wxdWI+Tjx+hsk24Ifl+Z027sjr/
8h5LZFgij7PXmFoXxIhmocZwQh1xH6lPR5G3pD8jKzsayOOAQfQQIHvcfLICHLmz
scL74PJ2J0I7I12LrYmh64JWPoDdxz7s2NLLFzYd+LMKM3AY2/Cf2lF1IWzCeuwG
zvoVIJ6AHUW/Ws2qujBkbAJ+vJKJGVXBkYHN9njIK1qIMlfYpdo/IebGiZZgsWIu
aTleN7ErfIPU+iqJnbWN2Pc/IqITGq5GSOk5HvrroBRbENob1IvaX1yU2L3FUla1
pI1h8BlL8Wp9nmu+HiwRoJNkSyBq85hi2hXZVg3gAFK0veOhr3lP4YPQuMA8wJGG
r6AhBGKZCQ03l2w2lGkBzrsiqoWcugSPwkoeLd3keQrLykZrjNhReYsJdQcAqUpG
huF6uS7cpbZTAET+Toa1I4cOXJxNz/VYqzHSdWhnaEN6T1VExEIlmel3x2d2sEuL
YYXVeCcxooshunl3tXn49z2jSlCEa4f6kZmPMz3Nw0sxuAQOpcSYG/KRey/VnKrT
ggjgL5xICvJHYjIbJ7XkCRXFFlXFV0JLGFAwlG/Wzs2928r7CIsOlFTEBxcTBW+0
0f89B1E/uQJ5/MxTHLfjmRREWiGXadi9Gt8Q2/5Eubkd8awYRGbHVTLUGUcjNP3T
XVLmY8wmvh1PhV4uDh9/ayYdbM06LZALpAjtI9iyf4NdcTE4CMUVCJq3+59kb4tD
GKhNJoz+ZS9TIYE0Sz8vtqO4l63cLN0w3kNvLVfdc7DSjDBtq/2P2E1AQb6i1GKk
HBjl39OvixcW3oLS2YKibANmqEnJfv6wy/xcMGpTV2jAbzd5xSI89fj0Xyn6kBCF
4ZVQ5ej2XupONU6Bfgkm4y5HwMrkqdJ81BdGQCnMgGPxumKftd9pVTgtPKRGHZ3H
2dAJYdYT/VLuQBzJfJAlAML4GPoQeYu7zPzILxjF/jarCfgIFQPy3UpPDzlVHp3K
xo3fxGhIDPhrujVd7xcM+1989CZgNfaTumOKmikTj0udPmrIDxEym6M5F22KeNou
lM5hJhzq3IDnvVYG/oz0QNivZpxmrCaX4qxunsVz1p+Ro338sjQBuFExlB0V1olI
efYEThN9a597nSiE9em6mRImjyAjPR2K0Hw5az8/3Cfglkm3tvEaMWvdHd7GCG2w
Vr6MsOA013Uw6rvJ0qFXCrS8jy+I/vEm6F6Y9FOZFq0Id9MNKp2zKldDwzrGrV1s
Oa9hVePIUTtITh7tHLgkuyuA1HEcQLnJJt2iFHqxXGE5zXq1yNAJMn2phjf/s91X
+P0ZcvxQxPAc68LL2+FhbINM+fc2wTEJbbU2OIHokaTSfTL/HpV/dJ/mLL1A5UsK
sDvJukknWyVGHr6Gzg7lmNapcL+8pCCD66xntdBRODKzmDTN6MkFE1fSzpaTJgEK
ul6V/suIZEqWxyuYkZBoKYx81bnajcTlnKtqc5MpUTo0cAXrrCfm1xFJ4v7YLCnd
2o5zBuS6CAwhlnnzj5EyStdCvjVG+PP88qVekb5UV0J+iIcYubf0niTtc+fkHfOH
gEjuZhI1UTqiOXJPIMFlYg7DoAF3VfnemafkTx39bRWvtHQe7mBX907Lfb4e+Asj
XdjhT7dLJQcseK08lemYZ0Pa+fqt8fXTzVLS9nGU7/5IkWVgm7gNKygeJNOd9OgL
vX54zGbRYfSHXnaLN1/oBj097fZ15ckNwYHBa+R8RLlB/wSYZb1KAVO6hjo5VBSJ
7+PPGH7WjNPiipJSTX7/x+Ajx2dtqWA37CvLysiCIcRVLEUHsqo+QjQUe8fZXqUQ
dLh6SGVtWCg21p3qBWCTdCpQZ1/FP5cVgbGkR2KdXISQWZGFZBxwa+OHlODzYDf1
n/JUXpWjFvnwCZhP9cJNyUrmciDNwii/rZTrho0QTOQmbjQ8IVBwovN3oTcyEMn5
kPT7NWphtQLA9z1mCnRJcW6YajhP1duLeQg2N3ZxWXcrx1iYRfID0bVKrLrAO3At
vs4Symr6yeD54/YGMK+p8FjD21SJAqRk9gIPAl+FGb/X8ypyZRoTIxfUaJMCCbuY
ScM7Z+DqYfsqjbDGpkgZKYEavUrYKAnqH0NcYCs+ryOw0SjnNlJlTE+UOjUuajjM
APT5jfyrJS/UWKcHOq4J9kwv9K/xOuarNEi7MGPKnsew1t7dqV6gmz2weLhrVkKs
K5CZBYp9inmMzlXQVu0ChzmzSU4s13rOveqa2B8KHUpMDnqioWbrnm6Qlo4+6Wr0
uB4nluZoJ5tlIXFsgv9yYyoCXPW1TQU5YBsXJOysJAcWPSijuLF6Oy7f6OjICnr7
uJpNuyLu6ymkYq3vokTNqdGA96f6UCGyNxW0t8392Ngb73HbGhaLN13CwzTUn4tH
F/248k906WH+CAI3cZ+XQYCCtVxmdHZ+e77Fi5oreawXUJYK5QQjLG9zy74nPKrg
QznkJd9Hs7ZTIWa/uCvalFw3BwHWP6dI9l35hMRid67Wob03JlT73NYnq8qbB5RJ
xN2pyqDwrcD0pIe6U49cBrOq4m5L4o1BHUcNiKjudiphpzKjFzexXiSi7GbjtIud
CjAbH50wgK2rN3xqQegTJB94l7WaVGe4/IXmlpxwiRH8fHnL7W2HCWt6Kup1nbJ8
3JMxEr4NrgSgGdqIbe7G5GETQQLDEr2RkksosuR9yRfkyJuGzNzmBNoxgPu4bc1d
DsOaJCHRTfC6WL+ch0cX/DHlYiHZlu0PIxgRcTToXKK/gY0Cf0UZJyzd1pip7j0U
WmuFtHNp0yXIjguo0meiynu7HsNA5YLuKgme4eAss8cVPngCKpLnoTIvcJQvQo6O
q/aP1dLyOTiSuXRDYHjAgx9RR/uiCYpXu8bTvN+JBkWJMi6lq9n4G19NkVhR0vUJ
RdNkrXLUeFPy7wY+Z1n/URR7D0jEFEjAI80pLL543Tas8XLkqMcZkhNCfSaerdW0
o3RT4YX3VNDg8cF0eOPfRG3KOflrtRFv7+0ZlFtyLHqGMaNJTw3mIWQoVerxWGq8
r5ZWMUcy4BHTkcgNJq8AzcSfKP9mrVCNT3FKpUQ6kD2+nCcZ+ggLTkU2GDnTpxak
AziqBccOPeZhZcv0ErAXit/RPsqXhgzvKu+pBPibfhep9riR9GtulBOEhIMMtloN
Klev4ytti6cGDt9YZunCAO6B1ZtNpAJtLFUfvM1qlOBRtE7rnEWA3gSadSe0qqCb
dm4UH8YDfVZvcm3PJ7mrws/7gO9POYYA6/G+nXD/nLwaLi8gDMEmd7bsQW536cDe
ZLqPgAZgbSuREHhlWE+qW/M0cNTjzPowtSEd5znGHs1yJIbtlQCdVnD3xQPHvyoD
CTABz0cv/JZmww8bbZnufUQuTdgU+MEkS5KiBe5OIwHIksC079X1BBb/UFiViszZ
Zq1FesGKrtIkHRKSyefxPEyWzKN3rV1zFYB0xiuQP03IwtMHjq1ruLkcnQHgB8ce
WZHjdq6YMXfljTg1gUow4xdZKojdf6Y2qbQTKG/Gg6/GKGLsxnxofjwMhpCZKIVT
jbSCWQWO7OCQnWI5+97kE7Hm2+IRAD5PK7b/JHTT/VeKUHACR0Np33kn5OREG55D
+j6YuwA08P7Upfv/xwjTFMlfx+H3NG7qvXJv9igZfe005zkNhjQ4EoWkKXHEzJdz
ztjfU8gXajEDQH8Xx0MBpRmpnQ0NxGKI3AIXGbMHHbU8Y/W72I+TlxfixOpYP/Y5
9La7UAXjAL44OoZrSEJAQjM56nDdbMBdS6fu66HgjPx48IBsPW7Hrut7M4KxACDy
mjnP9BDo5gYEqgGUvk127CWXWEgkJ6gzmWEBDYZuawzic8foWHF+iLrjaqyGSjdA
dDUpPkQBd55uraL0W3LRP+k9boidKrxrKT8mJo8dLSQR+Fu1lyIYkAcMbe6duxy5
vOp5JVZ6UBUa1WZUedXYua6GkNIIR+u6pEbWkUOTzRsn6RxXuvQdt5sfUw8RH7yL
X4yTMU59b/bgLbfEqu6hhbEn2f0k2uyMBfs+0B+RX/H2R2Zx7lhgmkPRViUXqb+s
jIwyKP35sT58/TA6clh2gI/uLh5ilXRsvTVweFp+1PDhtt1I7zaWD/RD6BdEXpWg
fF3THsLRCPZSCe5fQaWxr/U8dZYLd+t233v4rNDKB7qjStPRwvZMOS5JMVqZYKYL
ZE7xL/hAp4AZ88+zne5Ygn7b46GWiCJgco23ampflS0OMAQRizSDcKA/RwcjIQGT
GfDbBp8XbIg9BnlBuQaZq4Q9FNd1rbEI8/dmDpaAIDcph9R4432+1QeNbZ4drCSs
AYjRt0J5Xw5tZ9q3AMjAgngV5UsbOHspbvn9ykQrOXgDWqyW4afrgeIjwb89UCz5
Rc5jP10svivl63rz3CnIg4Y7xS46oEzQhtCxwms3wD6eMttVMGHCZZ5ue+rsekVf
dl1Ux5wS924M78cZVRtnXVwVJvvcFwfxIMEZr/z2tcMepDjRT4kXMALKiUw2hCHc
MF1PB5Sl0nZi1i7VGFJ4BSJw7uquHOgBXcgoSVE2mTRjhIwuO0cffMXTMKpLleuk
dDDmSeutNOZPrxo2DxSaAR1zh9X+IXgGk8A5gFAYRcO7PgHaTVaOtheAuyWIWCIE
MgYBipAX4kf7slkFYq/BZJRUhvsebbv+gPsZ09eNOflOzF0/oKlyBeXz97n7vaOX
juWEO7aK0eUXLm+l/z5Q3qMSqUHd4q893XESp/vDb6FoAAsrEWix7tX+SlR/5GgZ
bUC/GjKB61DbZBQE548g6d9aieUd0S0YY7vmXtoLijlrt5J0toAkGPICtkxk2x20
MTyOiOCLhG3BiG6528hvyy2PncnRDZ+0EORFCSkP7Bcw2013xpW4ppHStwpySCNq
Us5cgVgiHZlu4/f8lu38raahVt/NJnDvjZMW5z/Ea22k+n1Z+qR5G/26M80rPAHy
f1wYs3tM1mIlS7n2nI60WLiiTR/XoXZcgkM3SEv1NaDbU6b6S16Bq5//8SwUxdK7
iDzZe5IKcOUh73J64F3AGX9Rh7wHY7WNTUjHv8dHFwVbnNSd5ljn/2a850UnR4Dt
jJnV+82Zl1m84th9OGPy84mZTzk6rA1Jt/RskxsOIOhKd2J8RH+u4Zb9w1lYgg5n
jQ0TjIHQgsRPXwW3zWXgWgnqcZKDkJeflSf2dhgvb5J/jneVdJhW3YG49A9toucW
//GGEFovHPHl4tgfAIALRsL2n/lCL4Iheww4wLRUAXf0YvLo0vjlCiNTe253U9r6
9aG6MZ705V22YPa9/ofWCVeKNNwl+ngZPyru3pNbWDGJRUUeawT2RQGi7BOvC0pl
G91J32lJtLh/ycC7+lWOfPv0lyYkVJ1GxKRJ0Q6wYsCxkQH0aHcvJnL9SfK1ICes
dQq1A2FwBCAVjSGhP2CxHfaVPwFpBr9Qpnal8XGM9B9JZcG/vRjV0vDHEazhbtUt
aBfvuDihaivFrLVWOGGkfQ==
`pragma protect end_protected
