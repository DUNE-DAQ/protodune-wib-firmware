// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EPU71WlfOasDhHrzKBy35JoiOcYkAwCTnyQpNMZ6lm23rHe58il8Nbtp6zO5kwpn
8KW6KSGQq1Ii64gUNOmcBYsNoojA0LBe+wGd01W9PsHLqSASQhQCtUBWEPUv9Fm2
plKbaOFFWAUqmZbX/tNKiqdpYRV8DA1k9Pk9qbYWCb4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9344)
m4x6ti24JLiZasqXC4DLk/u41OpN2jAk+goteDW3ZVQVRbvKOHDkcv+HCTG5T197
IbquxbtlOrL0e45Np0NKRmSt5aPGEg86o17zpKy1Hzx3Ew2MaaQ8oGQdY5PTI5UN
n8HBKmyInpVhlIvVus9xsSjuRUwhaLr/v4JyZ2MVQWAjEMnxdO5Vt2rT6B/GB9aR
dLFIf8Gt7zpfIKPbh4+37UGzH1C4MoPcnu9GFTBpsde+ljI+TSxqBDCzEQW6LrL+
co67c8JPXYztwK7nHZpGpA5CIZeIoyQu8jzfmRIpEeMUVslNtoYwtOx1v3FBVrH/
U/3xuTg8YfsxbvdLInitQv5uj6AJEmiL1WKGAaZrPL3qxw8spXXQprwOaqbqF79V
r9ZcAKZX2p0CW5kt23MZHj023K6CSxREHuGI+6AKQC+T35hp+ykaqo2Eu/4TPLY3
py4Hr1ndeV4bpegvPLL19DLo0raqfswH/toJI6gyGrUFCG4H6l/dlf0bBiimY4Ug
yzIFskYOuDgz2ZlwNnDM1qOQN1YwjR4MVbFtFXPPLyUtsk35g2G/0SPFc+QedMjy
4B655qGNavcCdOVZme39eh5eHy6ws5fKtqdTBWvGUVxIDIwUUKqjEvekcoZBCKLF
YOeuu1IQkgGib9bOaQa8mLjdZvkLCLgTGfnl5ph/nx/uILFtI97h65/TyhdNrkxh
xHOaorp++zCy1WgmKilJjckkVVoWfCk/bqEtHmajXF1s1d4j0nALhQKkkd832cAG
Gz3kcQLCdrRNBLiQs2vh825hqwPKpsfGy9eGSm7psCvjmDDyIDbaaE/wwncbND1I
7WxCjXNDpnThscjLBPGOYI/U45YlSFNQSVLSzXIE6t887BAEUv+MuXAXFzAj+xPJ
Szzk5qJQkaNs0OYljwpySrz2LBAhaMyAzRuY/KV5Tsnh2Rf7rRr72L4tbBm1mNLM
BKMoE6johQNkLL8RiITKGMWN6vt93tX7Mze/+qzY0NpFjXm8KI7fS2NwHahBXMj3
wa+7SruNt1c6dBaStPpBB6qAMIfg6nCWDSjH/Dm4kZZBgfB8opMT9Xi+VPo4Cy4g
GFVQjckqBg9gDJtQjI99j2GBJGbulEf1LBUJzaTa3LbL8zQTmLR4MINDxfgjYLZX
2uo1sPD6rudX+ArAWbYECpv609EWDzTqN/g5XxDvj5a4ClCkCez1oB+aWmLMxLeR
VAPE8aDSr1MsanATig23Oe+AECO4zE5IogZ0jy8Ouu/1g1BV3Qh8UvQ8f/5ejeXA
iy2N3OJSSu4OvMPvvJuge2glCVPclAdNwQ6I90auqI59FlowCwGS8xZKOsOhddET
KZdy+Z0jRMeRgpHc668shnDNUmqk+FOHsfD1+Xgj7DYkaG3zQ6Q2LNQkEX+0qHUC
Qs5a08I6L6IwkS0b1Wo8zS+q5z7meCsCJtTRTdnb7vXQIws1UMLyKMOF8mOW6oOP
CqcqxCAK4pu6vNGegX0tc9EPeEp2IYgsGaX/CShqeMw8BhHdI6T4qNB/RsDBAkc1
wucCEvCYEAgDKJnKev5b/A0Wj6AxN+jQY7gn/bVx7ok0I8zR0iqUhJ+G4lE6nxBH
keuw/RvIAEaZ0wBgD+CDZtqQCubdkw/1T1shRxQHr0y5aLILR9YIrf8OLxTvRqNf
oBJjzMR5/I6ZSSYn07ouDHPC41d7G+3oF1vwCF2WzTX9sQZaiGMPHFerjXTFI88I
RFTKeFxeoAxbVQJPozVefox7pM9SNwLr0eBngwz9Wk6kyxcBYRptcf5vUz9lTycY
1qXsVlQoW3ItPOvwKQ0qj3y5Jondo0cvpzoJh+yrrgWh1Y0spNdkVRP3ANLHS8BJ
kvZURMMDfJ5H9f8q8alUqGkj8yw+hSPE1yPCqJ95j65W3YoJ6aDHp/XrlRpVeo9K
jxI8BVR8EQ5gX/EMGmx+hRy1poe/7Y9UYYGKGvh05JwmsuK/Vlj3/ZBXjURiz3uw
2BPT/+JcZ2Y2hoJCdN0wOwoiBr6WSns3QaOAxjQW9UOxbHiPQAI92/N/MT3Djkuw
7SkLuSLZ1zCvFqAE1uhqAB/WjxujHSjQLeBOSeAlW3Ujamr+Ja5l/DOHEyhyYWY6
dmdPEEqsmUCVWXZ087LRLb2pZUGvlqIij1jDAoYDr6oSTyf5/uwo0Z+AE7U2S0Aj
YpxpfxreVCq++chshlHGr9LEIhN8F5L72+R4CI3VcVtFrMAFYrCYllGxWwpAmYPB
pWJj+e3dwlt7IlEM93LPtKieV5rm+hRcTZeAond8mOi0sZomHqZmjcEWmCDdvY9b
tFe/EcegBgwPQ5wldOYRFz/Fop6sHp/9bz6tpipfsypFoSLMtXTJtEz3dnEEhxtd
G7Hh559IgTIMAOhhbL5RFaUgj77GJMWgCaXIva8YCRcjRMV0FtW5ba7DgUZtXQtJ
YU+7bz+tSyl4jOchwglyT/RBXTwseQRs6uY/gKyR8RKg3wR4dIKfrjboXYYH9ojq
1DwZAkIaIUOhWnOS1O8ft0A+XUg2RF/CL+tprRDzkto8NizmWcejEFINO1iW1HJ5
o897Hx4czv0xAyP2FzlwxHk+ttonuQiEk4FZeTryHn49zFYlM0Eh+sw0jYqNgcOZ
y+EwLN7eJ9fT/YHbWExIh+juug5EnsDMP/LXBQszNSgzdQ/2qTDBPy2ddk/azEN5
EP2jGGiUI9zXaBnMWeGJ4vdPUnymOF95usZ22G8huaIXi4wTJMkAPE00XKsNeCBK
9OCALtH3pRwh6bkOovkEep6GYsq0gux+4jlsbLZnQa+GiKrIzCWvu4kgOIZzZbyE
3zUc+jFulB4iV6gNuIOcpOu7Z3cjHgi/6NGblzRBlFR/3zQXYAglnzOfaRHBdqvc
uqFHRmYFvon2SZyxP4+nZmJi21InwluQx0RbWcXbBUpxmzLvThHWpeohJeRSiUL9
0ZhRUcM8pZJOrRkADSF0kgE4yZH8+HWR+pwU2qU7nAlmVCwVu3+Z74qtSkWTbTaK
oSMDuAaUZqfRYgjFMIX4zatG5F2NTXuCQv/XLLTWBT4CsQyDxkqlwVemJz/NReBV
CH09WBnhwTt6WPtapL7PxjNPkOwDEAfezMzYR6jFg96UH/kVqAfQr8G1HTUFlJcl
XR6veIIofYnYXIJUUT7GB2rulidr6PlfJy0r3bLlF3nEGp4sgvrtw5hpHkivzpar
acMevTi8DLEfH4PjdMZblaRuruj7nx1N7f6S2KHmLhWOD/9+eVSa1LekMMvMiN3Z
BFmdB0tQ9skAZupUjluuukCrRo3XLszF5HxLeSesdeM4sSzcE1R6mvy2SJUYSJcP
9kpvg6blmqnBnA7t2LyKuA/+fGrEBSNumgPGwWdWH1wZzBBOdfcGdRpet/X3vFFw
XGieylpXtIqFvgzNjcbI0paj9nP1WQdGEnAExDPDXIHS9vxLqPD6ZzZwQFgxOeN5
GeQoZoC+dN55Qj+o14VWRsMGTsIkvZkOCqpjkEupkjc1GDNgctr1dsW8qVkndOlS
ZdDvzyU8B67NItMMV1YZVgL0nbPT223FNxId+JZH54IN9gvF/QRAYYu5TsdphI5F
iqVbR2b3oApNv3HFbUcl5FD/jp3H5j5vtkSNa7WMSbS4tzWYkH2Ds7MF/5UMLP0E
wOy7IBRZFWRu+d93CyaYotNnMsou9acIYQBaYgdQg0mUshHW7Cv3CKazmJrjN/or
d2qoMZX1c5gftPFPWdzHG8+PFPLc7MLlQuYaXpfkDTqrxxRNo08F4iaLMSFMaFhN
B2ei6npuqUsbgIRe//QKD61QxEacnmuRdnNEpV6/a4WYaydgx/Plk0oPL2yHVpQA
jBEsgokIB6/OXIsBxXP1HwSiOzOTQ8y5VHLKJVe8N1GH7ilmN3dNa9xJcfmI8FDx
AwQafwME8hvKcZVPNCJ00Cz2BUyCIsFzcrNd03UAkEVgr6Igp/o8JqPYX+PfRPwu
v7st2ROU0qb782TbdzNjpCtVglkJVp/GloAd0sse4JckquEeEVcyRzZm+D1HuUYA
nCdCIohZx33DdshqemyMrhH/e8ZsE2Uv2awF1+tSu/+UId874p2WYIVEOx/FRRa4
sbeREeuRvUf7CmG/RYrpNTjaSWxLyiDTBQTxoPuWn4RFPoeMU9UnBvYQk7E2T/L4
9tFiT9Nm+QvH5AiYJrEpeK0/Vge5ePAK8bAL4AJjr4dMPmMetSXcUB9AJlLwB/5j
16mgnyYP8BdSva7R+mDsbAg7D/r4jkJzCvlWnW+ZjlWfpASjpBQ/Z8gls+xHqY/m
Y/TU4LXR7gHixnd9xQ8Io+FYwIGnv088YbP9KxAG4YbJkBVRxM1NtOvw5cAqFzQM
QbA5NkPFsWL+Wy/OiOa5RBu8oYyUXB1gQzTBTMHL1ouAHdRnQFR8A1xtxILAaVyu
HYHoN1kj4O/2YreMhrTUfliUXBHsQHx6l1d5mH24yWcqSiEX0Q9z+GMzKpl48E24
7qysY0X4vbABtjaKsXeLQU2qFXFh5gCa8IMS2MB8mEWPJex24qgnUxHAgk9CWOv1
B9NlryijRYrcPEHqkkE2OThZPyQAIWldt/IOeQ2raNwNbIp4Zg8ywhMUX6M6tZzs
JybewcqVwtcH7GAvpHgvSWpSmHLE/i3NOLd3q+sWlP0QW4UoTzmcHZZO5KktS6rw
1zW0C2qRcfBhtj5GnEcEp9Vj5zWmdvqwy3YqrCtMGROrxPx+4f+wPlLb76J3ULhL
4cBjlWHwvU3eRM6Mf/CRlI/XZKZBKgPUND24nOPbZyFoT/10hrG4kesutdv1bRKI
al3/61yNm158WGKJd16wx4nxKYRriQ3TitO0p8c0XaUDJbTk8OQj/Yp/7TuBh+v2
x/ksB2SrQ0NNFeXZNhWl1F48MFor/kAq7fQd0ykb3WE+dZ3lK8gvrnVpxbCgy4AG
lJ4XSoXSW2PwkFRWEkQCtYH7l94dHXXdNV4/bKF1FiBNqQzd2yoy/Uka9O/DIvNy
w2apTEJ5oFziMC2cUghOxPoJCNJosF3B/6DNCdU/rkHvxVYldhHRYj36SJIvoaGm
MhMndHFFxBp4/EboHh02fCAd0pRHbI2LBLYBriNJxEeNe4+J3dVtK8bgOf4eMhdR
4A/DTE0xpL/gB83fNNqWvodbqoDjyp/Ho75zvlDOte2Jgt+pkWG7jOdG0kT1N7ud
ZhbHICQo/rjw432B4CTVX0FEIVkzB0nuJ2J2aLx3mQgwl1eDzZZDrckLGz1mKwwa
sHQdjNSm+TR6yKIZ/Wj0sSaGaHu3KiJ7N8vL9OFJeM2v/Sm15KS5o6hpqcqimMc3
OgsNMP4np988RcLxxJg3zjNW2jIMplhfTNpgN4uwuVARQgGglmh74GWzwNrj6G8v
yR5TkIlcsLSHyaY660YxxHrUozqZxeSzTb7bbGDkQqScDYouZjL09LO7QzBT6Lv3
Z74KLeOIMtJ1Totm/6Z6XcERma6dc1HpCwbrRjzH8SIFZzkX+KirQmJBqz13JEaW
07q7nf/7jFXibrYMMdcr0dE2vMBgmn1jAih9dyJOOzQ6yzI53OnkZevEipM0j8vA
dbQY2hA3B8Qefit5k8VoeXWpiVPCnunuiw1e5TH/GhvAnoDpdbxWB1QxJqAot/1O
EWx40rWdqPfgYy37saoI0FLEtppK75ZVTa5EbI2/1es7byn3zaNBq84Eh5tWypC+
ppyL1ThlzI4j1Uapo2Cp/ocAgM/VLDb4uM6c/XIlAUCKZ8i7sP8cl5pJB8S8CCl6
wnXgeTRZepsr/Zbueuypiab7y8CsVJdI33MfBYGo0Lb1NNSVx/RtUDLJ7L7nUEYg
W977iMbvbjlPZ+LZw3uKNrCjYKcghGbKZPVkcPYRYya10Gh286JTTVnD/zWoOM66
GDyVCxlBFhTPVXx0jgeJ95gmlpz6rnWbBmisBvUdPaZIcBM/Ni91wy5daONOsEpZ
muRuM6H6fsdhiWsUHhD5N2/RjXhj5cwBZtv3Oabx1wVMB4xFElg2MzFTTLCtdT5o
VmQvkqb4aDfAF1hmgFKDKpwZIDS/Ecxy/st5IXHsv4YV9tcEq1XdxXckUmLs24jf
Rf1DItXqX6nPxFWOzPkCYGitVrQi3HSKOHIBERvIELAla6mR7vxlE1n9lUy8QrFA
uqtJO73xBfD14onYYysbQ8H/MHie9qmszSfwTSBzPeIJ8+0Kx73giJMq7bEBmQf9
9cRdpLprzWIZoStDP7PCROiLfOVtHU5KLD0FTMIxcKMWnt/0jg7fpSvFV7gbZUx5
dZ8iTjl/TueaKbhxSEuDoNlkUbsfzIJ5SaKAOdz6CuIK1i2X+YQ1dElh+fTUUQAe
nPtepUCTxuHw4smnuzVrlp+NE9HPvIhqWsXC9d11ziLT5evoP56nZdmtNXiL1rAL
CTPgAXKDdyLcR7e4llncl2Qb9Bx05VueN8SQlNNXFr+t8Tt89XOpKe8znroE8QNF
0uYl7hlQvleeGnHVZEFM0s7V/dTUb3gRK9tfTLaLpJcUNupvPldkd2iSGyasvjyd
D/0DIjh9INXyfZ9gSa6jzjmy9slgcIIrnTtUJBjR42+H1PlvMTVSNshQ7UpiaYlR
bHHeaL4H+tlf7Y5Q835lnF1zTovLdIg/Arg2hilwk/QwgHz3V9A5k4Qr6OznSARt
NYDpnfXvjuYcdVTKcoEG4JsMiQbo1BAZ8ofVHPtPYPhrDGFk1kHF2PLq/3C45x/M
Agf6/jDQRK0YtLv2/hTpigOkZQlq77TIB8oRBfh13FojdvYtF02vZFPGe+ccEWpQ
EDlGxDRUswm4F3qvS/QFRVhsek2gOZGOyz9yuiNMlVQGVfLgR8jTuOnK7/F/Y8q2
1q97ylJ02D6hvEuZ0mrb6NIrmyjIcGSDS2+VDrf/7vA1VGK+OsPDs7A84uVsGPl+
vj1/DGUQA7+mJ8cs0gG75pa+VSkP4WmzyjOnToO0vE+BTh3KhewdIpCuk/GkEF35
wQhr1oOy6w4c9lhjVJGvhhrszaKCEru22sUtQRp1jH0dLNPkLMrCckV/pIiUMTPb
QhDFDPPpvJ1HS+mdk7Av1Bv/uykS4h5YpyM1GY6YyczGvspxEiPc+3Nq7aYYMmU7
eBzLdpgmxVqvPzlwWT4HglTfcAPLeZYkncIvB7iHrgtjswIU/thi/K1+VoxWFucQ
v4P95CJeCP0Ke6gAKqxD7C6KZEqhB+nd0xVn9Imsk9CaCFr4j47eaxxBQgbHTQoF
ycphRm1ns+uhj6FHWGX8MUHjyGr7/uPgPiM3NAJOt8yPYKPsvBdebRg/p5w+osXy
MEet5mdpPgFx63dVplvbqChuC1b7mEyotFe3nS7n1ebvgUp35ClGgCmsi9nqhkjA
lSUwSwOP1d/nZIXL/CTOA4dTpoc2rVQ8BJC/VkIKfEha61Hzf6PhpoorJ090zAH9
VdKRI2WCjG+mi9YRLPmdqb98kIbMMqfM0yUZ1uwmbeSWNx1c/OTZrSPnGMqZ3ZQg
/2Y/D97Jf6OkOvVFZKY6foUHcBMxY/kITDZrEARb9BI8kZVmGGI9JezG7ANPgt0V
hL8NqNqB/jz/mM+ulFqEWDVFBprV7IdEENQSbYMMTj87ZfCzVW3+dc6F6DXr9lCG
6bhqkAnqiJHvSaZG6ZrLN4p5N013JIwpj/ZqvDzg850d6USNxpqVe8J5LWg8mPJA
UKm+Z2yDVMfaJZ4/rLogrCyf+DmfkObio9w8Km7op5muQe7v0sRvo9rwN9zq1+F3
vS9RQ+HcZYgwRez4KkVle/gW88KmlHxtZajg7K97gPTCptcvgsnB+TdzpAYO2D+G
aNLV3zJjGFQNmqRKqeHwP9ZlIG/keAFLZnbD0jo35Lm2iQdyrJYOSsvdnaU6Bemz
gXD3778c3wq8FtAXb55RkGEBrlfo6pivlpqF5W0mjrfqR2dYnWmh2vBssaIocNoe
H2fJjx0uOEogRJk4PjzS8PLwOZa+yt2ylxiKoOEC5IWQE1cK5W/Rpjk8SIbd/Rzi
O8xR6/mKckN+DobHLtvRvjxXmPx8Ud7Myr5Fe/vQS5B8IT/EuA0Po6bD/5v0+fwT
sXlNu+WepVROj8X+ShnyeBto5YDsu1uEr+kWyrBFGHkywf8yR4mLx4cTes6DCulG
LxmiX60sh8h8s/DXGsQB3Pc7t3rIBvhV/si3FIk/paG28ng8e5gKCoDo5OTh20V/
haWipFWXUlPLQAcqw2p+RWtNozuVuZYxdwdFo9Ija45GR2vfNdamW0ltladEn1Wi
UuoicJIeI3X4vTYiKxBlRutC/T2aJ7dFPUKlk/bwpHkCx6wT9+Mc28ZqXyYIOLpd
C0ZXKGfSSUgfrTet/znFrC9LJNwIj8EJFmC9WgXIuyJdkSmBZRMwUYL+T5F36TmT
PR3I+DvOimH0+c2WT0nUwwWhwkRKdVMve9GDHNo2RGkh95s0s3vs0eh0f3Phtho+
0sXJ1lsj/X49lNOfQ9nAtINtqfWK+USmPPB41e8Q9TVWg+DGSAHrCODsy2MYHg72
E6OtV2wucCpxcKrK7zornR5ufY7Q76/r5fzh7cCKD9yYw5w+llG6DiJCKl3LLgIc
REKvgoFnBEScEAHd6eO99Fzj+cNZBiYt4O5xGIxfrXsnC1Cic7asuaWOxiNzhsCS
wW83A6Z9S5qDC2q5pSgU0/TgA6w4rOK8FD2elH4yvG/gFr2ARFBZK9Du2qtrDSFj
O7eJ7AgJ20TXNifGl80wdwVzkWI+XTE+bIoRO3XZtTJrH58UhW0Z2zSEp0Cl7zIF
2Kb+eW9WWfRyKT4k+tMASxlutQQe6kxLyimCtKWxrJ5XClBM2uS+hzkC37o4wQwR
k0KqBnI3z4JAcEuUSzEVjZYPsoz8dwrQ9UK5XAf/6GEJ1T/f5F6vD4j7Fma986hf
p+ASGQhatUswiQhgG8EuqukjDY4IgAHCu3T1QJxsUpxWy2g3tHxVlN8kf1Vh87Bs
VuRQwAkIuVM7eohHv7BUiHuKy6f1Ykf0bP1VMjWD/hjdqX8mXJvxAFQZ0JwwKOx/
xYSfss9reHCCaRaH/6UXyc91OZpv1obFplj688yiTCjGxkjKzA5CebHXrIxyp13f
G58PC81ZCYO2JYrYsIlWlQfTgEJGYo/d2ZqHaVsnbpPqe5SwzvThulFngIr/WB+C
O5/5Mg7LyqAOIrmMq7uVRadP4YIg4BuST7H8MakRD0a3qbJ88j+Slmo5VrTouXUX
ylu8qwto4bBIRtacxpBzB0VZgKLAdwmijoV2+h4NueOal+XdenQ5P8pMin0YuN57
A0KWFuTcL16wL/4obHG9j9enx5ofo6eyLSXWfDi+FThJuFrusIXkyzl8hSoX9sE8
I8QdNHFK+tAj7osgEzeAXyoEFB+3yEjYGIc+QOdo6rTqmPySgvJJDTW19gzIosxv
ethwC2BSZeRH7lZW5FoJTsi4Os62AfM1ZP5YcbJfZGabXso8o3+qXmsOkqL3j1Ej
YsHKj+qK0IWHiYE+Gv5MWVGHktziYzRiOcZuAvun48sAKup3N6BMIvmKL9rpt2am
WWBIWLwMNS+9I68jHXsCtzyx22ZiDXddekwE/5ilax9qREFR63pjnYj7cxTf+2sp
xkVc1NbqQHZvxFbte1m/94Bkih4UBGgXEEQho0WXOmo9phvJJP5SHxPfoFXY6K39
SXc3nFg1jTD/AdU6/5ujXtj/jLEBObSMWFuRrW/F5TJUrqeSaU28k0LmQSmROdoQ
jPRgMzZCsT/5o/lVBkgt+XF12aUcHe1CRMwwDhS9hTveAybZIfEd2gQAOUuwWug7
yCu0xhwz3h3lBGQI2jlVitDzqrdlRQPOukwdd2e8hrdt6kwAPHgVCPz1ZCDBBicM
ieNVTyT+s64W97z5orn4SqBLANKgVCksSp90PrlinCocLWixUw7bSgcKlDBjAQ7o
1jCiHs767o/m2X2YPCuCtI//+gdmJOr+W4cU9ySCCixxx2MSspRh/d2s2Kb998TZ
Hme2FKO282Mgtl51xcG/tLmGgQQiJdltaJXJ8z7XQ0/09vBAq0avHcfBby9WK5cW
uOmhAU2iIJ7ZnvEuDLNmGbkyIdPWrEDRCdk/C/18fhKZZozb+Jxmlo3IPBbbPu9d
j2y5TGx2bH0FSlIlBjSHfxO09vuLMYx1XAaKujsynfxcdsl2tmkVSIzioSLMMSLd
DXW7QfyJF4UNhgqjn5/CzRR/lviCdv+Oh3ibpjHiIOkknmPMjx8jDEc/2Azu2fpx
8TiIn+CLcfbHzqo7XeR4n54M4pGnFf/nTx0iq2Ioa965o4uUNFbpASTWhgr9IwmI
CEtimRamR+GCkMLSFrm+9WLZZOyKi7wiDcoRcUI1FCfnXrV++F12iijXJ/oboMi5
mksnbpCMtAlk7NNm9gtLpwZ436l74s9GlxZMu7IvKUHPfSrL/BoOvqJqzmSgLFX5
GBPt9RdK1bE/sOwTsFKk/Q8C2k9R2kAWa2JJCHVqOSJTJWpW12PkJGnYBgJbBCvp
1kjBFI6OVfBJq7cZHJT+isc/7qhdliYpKrGRLy7z/kzHOEK2TdZmjda4d6SsvgSu
4bDWDd87ym2gcOa+YgOB2Y3V67QFBJUGWFrp7e9HAnmtvs5g6XfASUIzMshLe3Yb
NuQcMDFa62YDlWnN6RpfKxXmWRxYXnEYiUJMKJyz+jb9kdZDCJqg2EYXY1lhTDcI
arB7A6PTk953MIRVuaaczx9stjS5bwa8FLyV6Y/x6uJ7TgSxrWDMIzBbpuAJCVrJ
OpDjl6pV790hs8LDXa4/cD/lIbbZsKLZ1y4sDOjb1+RIl61btTD4r8S94dnzIa0G
nL8Os8vl4A45PIvMwDrsL6CuIRzvHGN1VyBEzs31FBIJphVoVU4EubeFS9UeROdz
C+EOe2bm4Ml9fBot4HLSqhWRbQV0avJhXfRHaDWL8kK7ByVCMUH0c/vEmtktwOxJ
1k3qFMDjvjSwUS3BqtDibCB3SZTtTZAacOlVKYl3FMMb1UvQRlBfzTRdmypWNQdy
GFF8Hy1bJMty2r+HN4RanYK84SvijS2nqwU0hxWj/a+e7Bd/pvwV3yVpIioBh5fa
TA/kjZ4rHy+Z2s8q4YcUgpbXW2L+X2SRxSNc/S0qVZWzpKKVwDtTCD99J0LZ2Ht1
TqAGY9qW+T6NRQoHiqEqX87Bai1doRYzlfSB209+MoAsbGJARwTzldj8DXRW4q69
8R8NPhgrYm2YVwgxvtc8lnV/f+fiij4gR3wNPvtO2Iw+vmUk8yGMlSQ4szscl+0Z
sTeEisejc3CrOhhO8XKMUtIxd3WMKct1f44++wV0GNopTU+8WLB03IOBgpALi/dj
s/XAABP0TCF9jAJsYBn72qSWaKXEo9fCxW3/i+vXgkBBtZdLDmDGCjTRqm1uRe/b
9mC0GN9MWzQOwHoCzQ2GBah26/34zfpi93naEOjYioqMD/WSuR43UU2WItg99VhJ
wy2nELQkaWZlcvrBU9OiaATk6tfRtPpbnJRUs4M9ta+yIGXGQ/8UFLMep4LUXug/
GCOB1JQiKPyZut2P5xbRBC9vt9tX4DsFSdsmgRGrPL9Z5r/Gr+avo7eri+75KxZx
CVtIX69CegqgTP9cckGO/C3Zi/ydhcXLBinGjTghjQyfJMqH1E6Uxx0yugXkecC+
mHUQDs7gHb3S+Aj3cOA2v5ux2qa/glJforyTvOItU2ObjLBYgnyi3V2k8uxA6dMu
1yqwxOB+PG6HFA92stwispSKs12P6o6Kzx4KVpfSEVHcYlu3zISr8dlRIgSZg6Xb
oZPT0BHHqeb7QljJ292G88cBVeYx392vaUi79TuMx4xrDse7tVENS5RvcsX7gb33
zkPpuOzfJE9PySCeFHt7GMHKq4iARgOgZNnwKpK/kIQytj8xgjQTI8brImZHyz8N
Oxx6RBtw08Ec5t1Tm30qJ8eGwqzJXK9v73By/s3vevevjpKWFLfYsrtR9CPUomS0
+PCq8CWf7KCEukYw3/3ScWFR+LpH0idQpUHATswWwmySrBowCr/3heNj6T2h/J1W
s3AeCZAwJfOtpLNqHrcI+Kp3NrVJCUAHnUzEwb6miYaqoT41kwPmRI3aSMopOzMh
TZylSO4iK1IyRoc5mxUIE7SDL5IP2l0VEZUxKWoR+XWuoGWBWGcpx8MnsFnZFkpN
ZGdYx329pPSbbnxvWG/TTVf1AbVcNrlXWyt90Y4ErdyqGVXvoia1BgDagqgDwlg5
aSU7akfyaS8y1tI2qg5KQgJvcq/+e+OB/RPZPDhY387udXZFOfNJSwsI4bVorVFV
wXvJzweIxkH39H+UY37Zy6wgVutqn0S0EcZOuYidDw1INaf0zmiQlK1Zmp1XxrOh
bv7zKSjHM4dmQJ1WdDJyTDFfgMonduW18x4I2PjgMSsIuztYM5UwjMAhXyAjk85u
y1+/+K9j6pBGFhuozbFeKkaUdhtlTFFOPhHOCuXa0UY=
`pragma protect end_protected
