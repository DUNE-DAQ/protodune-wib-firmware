-- megafunction wizard: %Triple-Speed Ethernet v16.0%
-- GENERATION: XML
-- tse_rgmii.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tse_rgmii is
	port (
		clk              : in  std_logic                      := '0';             -- control_port_clock_connection.clk
		reset            : in  std_logic                      := '0';             --              reset_connection.reset
		reg_data_out     : out std_logic_vector(31 downto 0);                     --                  control_port.readdata
		reg_rd           : in  std_logic                      := '0';             --                              .read
		reg_data_in      : in  std_logic_vector(31 downto 0)  := (others => '0'); --                              .writedata
		reg_wr           : in  std_logic                      := '0';             --                              .write
		reg_busy         : out std_logic;                                         --                              .waitrequest
		reg_addr         : in  std_logic_vector(7 downto 0)   := (others => '0'); --                              .address
		ff_rx_clk        : in  std_logic                      := '0';             --      receive_clock_connection.clk
		ff_tx_clk        : in  std_logic                      := '0';             --     transmit_clock_connection.clk
		ff_rx_data       : out std_logic_vector(7 downto 0);                      --                       receive.data
		ff_rx_eop        : out std_logic;                                         --                              .endofpacket
		rx_err           : out std_logic_vector(5 downto 0);                      --                              .error
		ff_rx_rdy        : in  std_logic                      := '0';             --                              .ready
		ff_rx_sop        : out std_logic;                                         --                              .startofpacket
		ff_rx_dval       : out std_logic;                                         --                              .valid
		ff_tx_data       : in  std_logic_vector(7 downto 0)   := (others => '0'); --                      transmit.data
		ff_tx_eop        : in  std_logic                      := '0';             --                              .endofpacket
		ff_tx_err        : in  std_logic                      := '0';             --                              .error
		ff_tx_rdy        : out std_logic;                                         --                              .ready
		ff_tx_sop        : in  std_logic                      := '0';             --                              .startofpacket
		ff_tx_wren       : in  std_logic                      := '0';             --                              .valid
		xon_gen          : in  std_logic                      := '0';             --           mac_misc_connection.xon_gen
		xoff_gen         : in  std_logic                      := '0';             --                              .xoff_gen
		magic_wakeup     : out std_logic;                                         --                              .magic_wakeup
		magic_sleep_n    : in  std_logic                      := '0';             --                              .magic_sleep_n
		ff_tx_crc_fwd    : in  std_logic                      := '0';             --                              .ff_tx_crc_fwd
		ff_tx_septy      : out std_logic;                                         --                              .ff_tx_septy
		tx_ff_uflow      : out std_logic;                                         --                              .tx_ff_uflow
		ff_tx_a_full     : out std_logic;                                         --                              .ff_tx_a_full
		ff_tx_a_empty    : out std_logic;                                         --                              .ff_tx_a_empty
		rx_err_stat      : out std_logic_vector(17 downto 0);                     --                              .rx_err_stat
		rx_frm_type      : out std_logic_vector(3 downto 0);                      --                              .rx_frm_type
		ff_rx_dsav       : out std_logic;                                         --                              .ff_rx_dsav
		ff_rx_a_full     : out std_logic;                                         --                              .ff_rx_a_full
		ff_rx_a_empty    : out std_logic;                                         --                              .ff_rx_a_empty
		ref_clk          : in  std_logic                      := '0';             --  pcs_ref_clk_clock_connection.clk
		led_crs          : out std_logic;                                         --         status_led_connection.crs
		led_link         : out std_logic;                                         --                              .link
		led_panel_link   : out std_logic;                                         --                              .panel_link
		led_col          : out std_logic;                                         --                              .col
		led_an           : out std_logic;                                         --                              .an
		led_char_err     : out std_logic;                                         --                              .char_err
		led_disp_err     : out std_logic;                                         --                              .disp_err
		rx_recovclkout   : out std_logic;                                         --     serdes_control_connection.rx_recovclkout
		reconfig_togxb   : in  std_logic_vector(139 downto 0) := (others => '0'); --                              .reconfig_togxb
		reconfig_fromgxb : out std_logic_vector(91 downto 0);                     --                              .reconfig_fromgxb
		rxp              : in  std_logic                      := '0';             --             serial_connection.rxp
		txp              : out std_logic                                          --                              .txp
	);
end entity tse_rgmii;

architecture rtl of tse_rgmii is
	component tse_rgmii_0002 is
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			reg_data_out     : out std_logic_vector(31 downto 0);                     -- readdata
			reg_rd           : in  std_logic                      := 'X';             -- read
			reg_data_in      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			reg_wr           : in  std_logic                      := 'X';             -- write
			reg_busy         : out std_logic;                                         -- waitrequest
			reg_addr         : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- address
			ff_rx_clk        : in  std_logic                      := 'X';             -- clk
			ff_tx_clk        : in  std_logic                      := 'X';             -- clk
			ff_rx_data       : out std_logic_vector(7 downto 0);                      -- data
			ff_rx_eop        : out std_logic;                                         -- endofpacket
			rx_err           : out std_logic_vector(5 downto 0);                      -- error
			ff_rx_rdy        : in  std_logic                      := 'X';             -- ready
			ff_rx_sop        : out std_logic;                                         -- startofpacket
			ff_rx_dval       : out std_logic;                                         -- valid
			ff_tx_data       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- data
			ff_tx_eop        : in  std_logic                      := 'X';             -- endofpacket
			ff_tx_err        : in  std_logic                      := 'X';             -- error
			ff_tx_rdy        : out std_logic;                                         -- ready
			ff_tx_sop        : in  std_logic                      := 'X';             -- startofpacket
			ff_tx_wren       : in  std_logic                      := 'X';             -- valid
			xon_gen          : in  std_logic                      := 'X';             -- xon_gen
			xoff_gen         : in  std_logic                      := 'X';             -- xoff_gen
			magic_wakeup     : out std_logic;                                         -- magic_wakeup
			magic_sleep_n    : in  std_logic                      := 'X';             -- magic_sleep_n
			ff_tx_crc_fwd    : in  std_logic                      := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy      : out std_logic;                                         -- ff_tx_septy
			tx_ff_uflow      : out std_logic;                                         -- tx_ff_uflow
			ff_tx_a_full     : out std_logic;                                         -- ff_tx_a_full
			ff_tx_a_empty    : out std_logic;                                         -- ff_tx_a_empty
			rx_err_stat      : out std_logic_vector(17 downto 0);                     -- rx_err_stat
			rx_frm_type      : out std_logic_vector(3 downto 0);                      -- rx_frm_type
			ff_rx_dsav       : out std_logic;                                         -- ff_rx_dsav
			ff_rx_a_full     : out std_logic;                                         -- ff_rx_a_full
			ff_rx_a_empty    : out std_logic;                                         -- ff_rx_a_empty
			ref_clk          : in  std_logic                      := 'X';             -- clk
			led_crs          : out std_logic;                                         -- crs
			led_link         : out std_logic;                                         -- link
			led_panel_link   : out std_logic;                                         -- panel_link
			led_col          : out std_logic;                                         -- col
			led_an           : out std_logic;                                         -- an
			led_char_err     : out std_logic;                                         -- char_err
			led_disp_err     : out std_logic;                                         -- disp_err
			rx_recovclkout   : out std_logic;                                         -- rx_recovclkout
			reconfig_togxb   : in  std_logic_vector(139 downto 0) := (others => 'X'); -- reconfig_togxb
			reconfig_fromgxb : out std_logic_vector(91 downto 0);                     -- reconfig_fromgxb
			rxp              : in  std_logic                      := 'X';             -- rxp
			txp              : out std_logic                                          -- txp
		);
	end component tse_rgmii_0002;

begin

	tse_rgmii_inst : component tse_rgmii_0002
		port map (
			clk              => clk,              -- control_port_clock_connection.clk
			reset            => reset,            --              reset_connection.reset
			reg_data_out     => reg_data_out,     --                  control_port.readdata
			reg_rd           => reg_rd,           --                              .read
			reg_data_in      => reg_data_in,      --                              .writedata
			reg_wr           => reg_wr,           --                              .write
			reg_busy         => reg_busy,         --                              .waitrequest
			reg_addr         => reg_addr,         --                              .address
			ff_rx_clk        => ff_rx_clk,        --      receive_clock_connection.clk
			ff_tx_clk        => ff_tx_clk,        --     transmit_clock_connection.clk
			ff_rx_data       => ff_rx_data,       --                       receive.data
			ff_rx_eop        => ff_rx_eop,        --                              .endofpacket
			rx_err           => rx_err,           --                              .error
			ff_rx_rdy        => ff_rx_rdy,        --                              .ready
			ff_rx_sop        => ff_rx_sop,        --                              .startofpacket
			ff_rx_dval       => ff_rx_dval,       --                              .valid
			ff_tx_data       => ff_tx_data,       --                      transmit.data
			ff_tx_eop        => ff_tx_eop,        --                              .endofpacket
			ff_tx_err        => ff_tx_err,        --                              .error
			ff_tx_rdy        => ff_tx_rdy,        --                              .ready
			ff_tx_sop        => ff_tx_sop,        --                              .startofpacket
			ff_tx_wren       => ff_tx_wren,       --                              .valid
			xon_gen          => xon_gen,          --           mac_misc_connection.xon_gen
			xoff_gen         => xoff_gen,         --                              .xoff_gen
			magic_wakeup     => magic_wakeup,     --                              .magic_wakeup
			magic_sleep_n    => magic_sleep_n,    --                              .magic_sleep_n
			ff_tx_crc_fwd    => ff_tx_crc_fwd,    --                              .ff_tx_crc_fwd
			ff_tx_septy      => ff_tx_septy,      --                              .ff_tx_septy
			tx_ff_uflow      => tx_ff_uflow,      --                              .tx_ff_uflow
			ff_tx_a_full     => ff_tx_a_full,     --                              .ff_tx_a_full
			ff_tx_a_empty    => ff_tx_a_empty,    --                              .ff_tx_a_empty
			rx_err_stat      => rx_err_stat,      --                              .rx_err_stat
			rx_frm_type      => rx_frm_type,      --                              .rx_frm_type
			ff_rx_dsav       => ff_rx_dsav,       --                              .ff_rx_dsav
			ff_rx_a_full     => ff_rx_a_full,     --                              .ff_rx_a_full
			ff_rx_a_empty    => ff_rx_a_empty,    --                              .ff_rx_a_empty
			ref_clk          => ref_clk,          --  pcs_ref_clk_clock_connection.clk
			led_crs          => led_crs,          --         status_led_connection.crs
			led_link         => led_link,         --                              .link
			led_panel_link   => led_panel_link,   --                              .panel_link
			led_col          => led_col,          --                              .col
			led_an           => led_an,           --                              .an
			led_char_err     => led_char_err,     --                              .char_err
			led_disp_err     => led_disp_err,     --                              .disp_err
			rx_recovclkout   => rx_recovclkout,   --     serdes_control_connection.rx_recovclkout
			reconfig_togxb   => reconfig_togxb,   --                              .reconfig_togxb
			reconfig_fromgxb => reconfig_fromgxb, --                              .reconfig_fromgxb
			rxp              => rxp,              --             serial_connection.rxp
			txp              => txp               --                              .txp
		);

end architecture rtl; -- of tse_rgmii
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_eth_tse" version="16.0" >
-- Retrieval info: 	<generic name="deviceFamilyName" value="Arria V" />
-- Retrieval info: 	<generic name="core_variation" value="MAC_PCS" />
-- Retrieval info: 	<generic name="ifGMII" value="MII_GMII" />
-- Retrieval info: 	<generic name="use_mac_clken" value="false" />
-- Retrieval info: 	<generic name="enable_use_internal_fifo" value="true" />
-- Retrieval info: 	<generic name="enable_ecc" value="false" />
-- Retrieval info: 	<generic name="max_channels" value="1" />
-- Retrieval info: 	<generic name="use_misc_ports" value="true" />
-- Retrieval info: 	<generic name="transceiver_type" value="GXB" />
-- Retrieval info: 	<generic name="enable_hd_logic" value="false" />
-- Retrieval info: 	<generic name="enable_gmii_loopback" value="false" />
-- Retrieval info: 	<generic name="enable_sup_addr" value="false" />
-- Retrieval info: 	<generic name="stat_cnt_ena" value="true" />
-- Retrieval info: 	<generic name="ext_stat_cnt_ena" value="true" />
-- Retrieval info: 	<generic name="ena_hash" value="false" />
-- Retrieval info: 	<generic name="enable_shift16" value="false" />
-- Retrieval info: 	<generic name="enable_mac_flow_ctrl" value="true" />
-- Retrieval info: 	<generic name="enable_mac_vlan" value="true" />
-- Retrieval info: 	<generic name="enable_magic_detect" value="true" />
-- Retrieval info: 	<generic name="useMDIO" value="false" />
-- Retrieval info: 	<generic name="mdio_clk_div" value="40" />
-- Retrieval info: 	<generic name="enable_ena" value="8" />
-- Retrieval info: 	<generic name="eg_addr" value="14" />
-- Retrieval info: 	<generic name="ing_addr" value="13" />
-- Retrieval info: 	<generic name="phy_identifier" value="0" />
-- Retrieval info: 	<generic name="enable_sgmii" value="false" />
-- Retrieval info: 	<generic name="export_pwrdn" value="false" />
-- Retrieval info: 	<generic name="enable_alt_reconfig" value="false" />
-- Retrieval info: 	<generic name="starting_channel_number" value="0" />
-- Retrieval info: 	<generic name="phyip_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="phyip_pll_base_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="phyip_en_synce_support" value="false" />
-- Retrieval info: 	<generic name="phyip_pma_bonding_mode" value="x1" />
-- Retrieval info: 	<generic name="nf_phyip_rcfg_enable" value="false" />
-- Retrieval info: 	<generic name="enable_timestamping" value="false" />
-- Retrieval info: 	<generic name="enable_ptp_1step" value="false" />
-- Retrieval info: 	<generic name="tstamp_fp_width" value="4" />
-- Retrieval info: 	<generic name="AUTO_DEVICE" value="5AGTFC7H3F35I3" />
-- Retrieval info: 	<generic name="AUTO_DEVICE_SPEEDGRADE" value="3_H3" />
-- Retrieval info: </instance>
-- IPFS_FILES : tse_rgmii.vho
-- RELATED_FILES: tse_rgmii.vhd, tse_rgmii_0002.v, altera_eth_tse_mac.v, altera_tse_clk_cntl.v, altera_tse_crc328checker.v, altera_tse_crc328generator.v, altera_tse_crc32ctl8.v, altera_tse_crc32galois8.v, altera_tse_gmii_io.v, altera_tse_lb_read_cntl.v, altera_tse_lb_wrt_cntl.v, altera_tse_hashing.v, altera_tse_host_control.v, altera_tse_host_control_small.v, altera_tse_mac_control.v, altera_tse_register_map.v, altera_tse_register_map_small.v, altera_tse_rx_counter_cntl.v, altera_tse_shared_mac_control.v, altera_tse_shared_register_map.v, altera_tse_tx_counter_cntl.v, altera_tse_lfsr_10.v, altera_tse_loopback_ff.v, altera_tse_altshifttaps.v, altera_tse_fifoless_mac_rx.v, altera_tse_mac_rx.v, altera_tse_fifoless_mac_tx.v, altera_tse_mac_tx.v, altera_tse_magic_detection.v, altera_tse_mdio.v, altera_tse_mdio_clk_gen.v, altera_tse_mdio_cntl.v, altera_tse_top_mdio.v, altera_tse_mii_rx_if.v, altera_tse_mii_tx_if.v, altera_tse_pipeline_base.v, altera_tse_pipeline_stage.sv, altera_tse_dpram_16x32.v, altera_tse_dpram_8x32.v, altera_tse_dpram_ecc_16x32.v, altera_tse_fifoless_retransmit_cntl.v, altera_tse_retransmit_cntl.v, altera_tse_rgmii_in1.v, altera_tse_rgmii_in4.v, altera_tse_nf_rgmii_module.v, altera_tse_rgmii_module.v, altera_tse_rgmii_out1.v, altera_tse_rgmii_out4.v, altera_tse_rx_ff.v, altera_tse_rx_min_ff.v, altera_tse_rx_ff_cntrl.v, altera_tse_rx_ff_cntrl_32.v, altera_tse_rx_ff_cntrl_32_shift16.v, altera_tse_rx_ff_length.v, altera_tse_rx_stat_extract.v, altera_tse_timing_adapter32.v, altera_tse_timing_adapter8.v, altera_tse_timing_adapter_fifo32.v, altera_tse_timing_adapter_fifo8.v, altera_tse_top_1geth.v, altera_tse_top_fifoless_1geth.v, altera_tse_top_w_fifo.v, altera_tse_top_w_fifo_10_100_1000.v, altera_tse_top_wo_fifo.v, altera_tse_top_wo_fifo_10_100_1000.v, altera_tse_top_gen_host.v, altera_tse_tx_ff.v, altera_tse_tx_min_ff.v, altera_tse_tx_ff_cntrl.v, altera_tse_tx_ff_cntrl_32.v, altera_tse_tx_ff_cntrl_32_shift16.v, altera_tse_tx_ff_length.v, altera_tse_tx_ff_read_cntl.v, altera_tse_tx_stat_extract.v, altera_eth_tse_std_synchronizer.v, altera_eth_tse_std_synchronizer_bundle.v, altera_tse_false_path_marker.v, altera_tse_reset_synchronizer.v, altera_tse_clock_crosser.v, altera_tse_a_fifo_13.v, altera_tse_a_fifo_24.v, altera_tse_a_fifo_34.v, altera_tse_a_fifo_opt_1246.v, altera_tse_a_fifo_opt_14_44.v, altera_tse_a_fifo_opt_36_10.v, altera_tse_gray_cnt.v, altera_tse_sdpm_altsyncram.v, altera_tse_altsyncram_dpm_fifo.v, altera_tse_bin_cnt.v, altera_tse_ph_calculator.sv, altera_tse_sdpm_gen.v, altera_tse_ecc_dec_x10.v, altera_tse_ecc_enc_x10.v, altera_tse_ecc_enc_x10_wrapper.v, altera_tse_ecc_dec_x14.v, altera_tse_ecc_enc_x14.v, altera_tse_ecc_enc_x14_wrapper.v, altera_tse_ecc_dec_x2.v, altera_tse_ecc_enc_x2.v, altera_tse_ecc_enc_x2_wrapper.v, altera_tse_ecc_dec_x23.v, altera_tse_ecc_enc_x23.v, altera_tse_ecc_enc_x23_wrapper.v, altera_tse_ecc_dec_x36.v, altera_tse_ecc_enc_x36.v, altera_tse_ecc_enc_x36_wrapper.v, altera_tse_ecc_dec_x40.v, altera_tse_ecc_enc_x40.v, altera_tse_ecc_enc_x40_wrapper.v, altera_tse_ecc_dec_x30.v, altera_tse_ecc_enc_x30.v, altera_tse_ecc_enc_x30_wrapper.v, altera_tse_ecc_status_crosser.v, altera_eth_tse_avalon_arbiter.v, altera_eth_tse_pcs_pma_phyip.v, altera_tse_align_sync.v, altera_tse_dec10b8b.v, altera_tse_dec_func.v, altera_tse_enc8b10b.v, altera_tse_top_autoneg.v, altera_tse_carrier_sense.v, altera_tse_clk_gen.v, altera_tse_sgmii_clk_div.v, altera_tse_sgmii_clk_enable.v, altera_tse_rx_encapsulation.v, altera_tse_tx_encapsulation.v, altera_tse_rx_encapsulation_strx_gx.v, altera_tse_pcs_control.v, altera_tse_pcs_host_control.v, altera_tse_mdio_reg.v, altera_tse_mii_rx_if_pcs.v, altera_tse_mii_tx_if_pcs.v, altera_tse_rx_sync.v, altera_tse_sgmii_clk_cntl.v, altera_tse_colision_detect.v, altera_tse_rx_converter.v, altera_tse_rx_fifo_rd.v, altera_tse_top_rx_converter.v, altera_tse_top_sgmii.v, altera_tse_top_sgmii_strx_gx.v, altera_tse_top_tx_converter.v, altera_tse_tx_converter.v, altera_tse_top_1000_base_x.v, altera_tse_top_1000_base_x_strx_gx.v, altera_tse_top_pcs.v, altera_tse_top_pcs_strx_gx.v, altera_tse_top_rx.v, altera_tse_top_tx.v, altera_tse_reset_sequencer.sv, altera_tse_reset_ctrl_lego.sv, altera_tse_xcvr_resync.v, altera_tse_gxb_aligned_rxsync.v, altera_xcvr_functions.sv, altera_xcvr_custom.sv, av_xcvr_custom_nr.sv, av_xcvr_custom_native.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, alt_xcvr_arbiter.sv, alt_xcvr_m2s.sv, altera_eth_tse_phyip_terminator.v, altera_tse_fake_master.v, altera_reset_controller.v, altera_reset_synchronizer.v
