// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZEsNOh+d1QVqtSIXUzQr7sEL0si6NneKE4oyfKgfV3Cx2jpcv6Urymluv8ouzGlo
YAAl7OlwcOVry9itkfbWPb2n249k97st4OXND6YMvDTh66J/6JxiKZLDQw5BHyMF
EJzdxPuYBctTJ+VaiILt2KlasDm7+/8tJCCvMFs83O8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57024)
InCRGMxJxFusfHvw9XD5QhdMTXkfw35EDqrOg0Zt89CJU5qxZuDV22uGWY0d6m32
D5OG3SG1RULl6yIJSaI87CFGd0aaQzwuYHlSy5Tf1sh9U4BT0KgiMHg/pbs9YcrP
u3/zmPEqripOn4etDW/qBLuehopoCYMq2wuh/GfEnZNViYFJOr3fcY3wHhF197kI
JTFg2FzEZJ0LWfKQPCuViJaHg+kdl3ZmE/yCtQzxT/6jPWmrpmn6trKR/ronWv1C
Dx31aGqAhXEBLaFXzHuslYg0xh/SOZl0bT3Ji54kiEnhG4g2E19BcyuLPhlzxoTp
KPJVU0rlhHHdt9vWPKffEDBurmsMeRelfn9w0ih7oc/WZNHC8+icFxb/cdEDKtU2
6qqD6U9LGABIeS+i/x+FJrBLRQ1eFbAFKMPfRYUxdhx0Z47HwqmBDGseqNalDOCP
50fdRn72ltV7dxUTXSBnL6z42HLpZF4adbOr6Y27OG7oq7sWF4q+RDx7aglhXytG
h7wNTD3dwCCSup3wGVc85C/9ghcaXKC1/JwCbuN6BkBWkDt49I7ngj2D+sweXW/d
Fu8QHBMYTNOq5h+Aqh+Qk6ne7bx+3B3PMx1xF14yQy079tb8bebbxeeDGLVIpOOU
0DXlNwXXQWwVcKj6ED8MwgoLjQkMcA4r2UryIQqZXRWG/9BzjhXfYeORTzxRlEJJ
o8XrvfzozCNPpwJQLCQK4f7N7hFBDs+RPuHiGWZvwGSaNKBfR9yrVV7v+w6fzL12
Gx/uIT31CDGWD0TUyh/CcidqMXQ05b2TpvvQFwDXTQ6WVPeHMyF1ZVQ2e/DomxfN
dlTC30+EpVnG7Z7cfVZjK2nPSP6HF2y/C8rSEUzGoSSXuC+uL1ZJtLG/ToSKBN3M
zwMvst0pDUKX6YTSg3MJWr9m+3s7J5sJf8NAXQ7pTHGnq20aAEjnVemY9zJQzd4M
MQ3PdNiJU2CTHNbx7Lk6Jb+BA0FRS2IYJNMuc2fE+M59UdLg3f8nmqn7olP29pYi
CQO+JHVlYKTFj+LOiL/mK+xwlcfmGqi9xYtXiPzJocwzXPo/fZ1ABCc9Ovg5dB0J
w8HPvkeU6dRR5enIrusekt+yK/Ws9Yd/HhcTxqWdyLleDx73zwkXyYUh4zGP1uDg
WqRup/s1W4x5/3Ec6YQFLNvdbutFtGOAdeOFeu1NAIK/XvGG+2ODYGRjRaLWOZLE
3m6NBkqipZ155oPEBimJ2AOWNttf51U8LdxVIO6hO/o1isrc5jx2q4ofQEhRTcO2
suMq4qMJNkttLl6Lwc7+dtOT5c4NRKdc7H+o5gQt3HotXLacx/cRjeCQVme66Xx+
2nlcQ4Nhzkm//mErkg5JiE85l4xTRCoduedlWHkxU4Vpt2J2riq138v9erZvtd7X
IDTrn1puc60uzlXmHKx6hWZDeUhIsgoUL5ztrA3jLphJSc2RbRqByE4mQ8rdsDKx
PhWcDl7UFWurwu7WGHfa5zWex/3XXT9+6CgLpDYGwc9CJ/j6zcedKZutnr+k839l
m8wCEMEUOMLz1FkIN0D9i+Dj9Gz2yEVfEb7t/GJeOsJCET7+ygqGk9OKFQIwlk4u
1tpW7lbcvoLZ/1YGFXDOcCCE5ZIB+b5KrO7qJIDhaRcs813v6TLkg7iXNugdF4Z/
IQlxLcboUM9CI4Oaw0ed6ksx55iV32+RjmFzKicrKr6ouFpROitmBPW48byiDYSa
3v1ZiAObhhNE/h5ZUzbk/28JLk1SGjupQRa44vFMqneokOmck2QbJsFLygna904M
da5pTEjxeyEzvovfBIUlStx+wTuem8VeNZJ+/lBbCC07E7o//SdDh0lorBiU48xk
uZUedQNJ6cdfrARxgqFF08bSudT0cRgaQcppdiUicG1cntQOoexfNlh5/SFIHLNP
NeilyVHO/j2UlkcVV5HWMm2pkg3o/7qx3u8AAAqKL6EInVIVKZ+gWCyazyIovF9m
WqukvDI2xc55+QL+W0CtUFFPS/zEHS+ZigHB/3C5YxW81IgAQ3lFqZIeKsrLB4fm
K3mtmoGkg3w26AX0gamMQD0FdD4okGDU54hzkbVlcI5NCClbDgXh8I1OGdwMXOGn
JA9qrlxQ6rGvve4SMAKFA56rgma9agvyDqtAmKArd0aAtmRfjgw9LXyKsoTYAQ+y
sjrNpPfgWlpaQHM0mTFEWQhuxVPcC2n98QbNpqvz3acEOyHV99hbV3rs6IXz2F/x
mGM1HS/m/u5TAKCgx4XPnzkYPupChgdgixRu81f99VOHt9PkP6NnDy0vbSrqDvuN
bfdHFWNW+P83k3Y9wCe0NyVZV5WGUViQC6QchOqmxKM9mzFGfCI9ggBOs/upvAa/
TR+j7kj0aYFPguYu+QKi/8CJYuhZKEqlOo7l8AhuyHq7/O3MW2YyMKfvGiWuLxo5
2H1bMpuOmJJdvlgxYhi0o4J475YSgW4XoIxRXeEjJ0PEMfWL6tAT4ZNXZjFBOk3s
XHohFWrKcIuOkqmCxoe3AOl3oDDIKV92dQrotsx5SF+VcLpmeJxAFsbaP0UD+NRq
lu87Pl6lC2DZbSj6cMOSEJ7ohkruGDmSniyMdZRvqt7ORheY/DmLLSLwUQ4ixUJp
bfiLw7VXPgDuQu442jxJ5eUStlqIbcPqXyHxZ+NaaqipTzkbZ+m9uyqkhdZWn3bc
ay6D2Wqqhd1ojr4vPL3A2w2yc9S/Ohqdwc3PSzAINw2Ipt7c/mdv6SNnjLtFxqmW
UjhJM8raaV1FpAinYfbmsaGqxdCdcFMBfZwG7Nea5xbZf9/JADCxGh7EGzGXjglZ
mgBNLbYSjMJ5X4ci/fms27GIFevsahIsZSAaW2b06vMG3OAJMeFoW1OEaqNUC4FJ
q8+9Xdkou70cTSS742LuhncEpe6WSY1PnTLOhiWjJv1+k4Lkfr13ulSN9bp9U6Ja
AjU3XNegwW3NE20WyI6EiymfYJT9AF4MA+r1X8+BgOz05Zdm2Ry1jW6SlrjEQ94V
RCCD4lz9yWRauRbP5lIM6WAvs/1hKBwyuVO60YjeKi3j+2RfbdW+DzI4yUfjor2+
b3wm/VKP1vm5xzt6fg1LV/6qrp4SxlqW+8eT2jqm2EYDuqX6py19rRF5l4vtRTvF
4IIsC4ZnfTK6gs/zlyR3LJk0wwJOkc+hw/g4EvfLPf/IlaULpy8xqfSkJ9OFue60
8Q3Dp1ajSNK/izKnnDjvTN0c3YuCKDqCsO7g2iavpuZneNPPr8s8dIiwmsDqI55G
2lH5xId8LAQVvnbbVop9YxDyuToexb5dfPY28hUExV5HyMaQur5dmi9WwZjycYMD
pC7QCc/9jRXckdA71kf+Uf6WGI/th45vvHO1hKcZoCf/5Oxx/z+YPhgHZpE8CQEw
Kwu5KwpotCCMjPZdopaLATR2ufFhZCq5whiIc/7he7NLJcHdAUZc6wEeoE+vxUff
H7tQpCl0UuBWfr4K2ZO+USXLrxRgbRZCSNrKMNrH78Es4dH1XI/Jm1R1gtHKXJSb
zb8XUfZlovPNQ0J9mat9hfvUOwzIWqPJUqDRUSqhSlUBwB25ekYfqKgah1fuIC7K
/CVWie8hJgZlnoJPb3QFUB2sMbLYVxqaaug6QgPW8U4UCqAjENkd+By61cMgODTB
C7aSD6Xk6fVbauT+SL2wNC0L/wHNMgvxDUuuDww8tS5VRQBwfDhznkr6lIew5q4K
UzzPwx5gVErw5Wt/Chf/JhN7YedAyjVleIavw8F88cKLgVRqUXMAVlJzepZFGXqz
PgWkxLjXeJSaJ6Y9tDNwRQkZ9JapHdXoUM/kKUylwX2+ASUhR1ynHNWf8ofXPlW8
JG5asIMQJSADuuLUs8QUFTOuYMdWS+3M2wliq1ghjFyFr0dTYTkefnrN6VI2DIGk
aF5YDfPMHO95yDXvT6DvyuMF2TCxZgjSfgOuBE4/9ur6twEGhxhEeKt+9PnzVtyq
PQupl0fjrz4f4jtryVK7F4dLBMenh42guBpTcKNnN5BH1eVjATDNAp6+evjd+Tka
TRvIc2nKj9GyGRLgILvcFDMyfWpNKMooPThe83qbuNQ20uCpwuEeL8ZqE9x/WgIF
f9SHvdR+3vbdUSlCXIPVPjYWliI2pfaxzq5YhmQ/TyosnduM1s4aux8AruGtk/el
97mGKB0v8lyvXMq++GAYmqvWhaOUziPNjhZqhbkmhMiOEjwW86IqzIY3/pCOFjrh
Vn2gYAp1dQlnuqwgyz/B/APwcQyBYJgLASu9QopL7ecy+YrdLepD/33d1d7WYvJm
kkfqaQpdCY0fOhcRxfaanAqLTYovynqR67Igxah3GOYfjYD5saTHN7yuqVywelHY
ULSJCL/SeArbE5EOZvrAy424X8STFqQc65K2IQ+2Q3yJH9rkBEnit9VeFGmgPk6w
2Ru5BZk/N4dot4FWeSqojCc9p0x/yFpw9zNaArVP7m8h98aIHFVUSPmXZJvULpsB
vZ8JTfZPowvz6z9PDx+L8d5n+f1lYmg4I7FTy7c1TeFDr9BtZMfoUzpNANJxSQG7
0DOXQWSTeiKlJreY4RbV7pC2NFX28g98q3BWQSRnxvrmmby68uRYW67qUJ8wCeAP
UvTpU5uIep58fsqF0qZ74uvOyeatAxKqF/GsJOkX4mOG8S9uFUmcmGByV0TzJDTP
iHSs+skdKmDqQqndanjcIUL9MZaNxxrDPsGIt6qRj3TbtZMNvQFJBwG7bpUGZXWl
TSsa+0WN8r5tXK7/THxWtlW/SgJExayF4agcTfd65scZ5OYTDPQI4lvKcp44fWof
8EaENwBUXudSuDWNgVcjKNK2znDL4kx5eJPQnFhSK39d7ewzpaEo+WVkjMTDwv6v
VtoCvOR18yM9TQnA1gILOCDEQwSIHp5vgwnYWb+89h2OGnPm4YihK4jX0hF5Yl6g
2VzuUYp4AJdmi9YDhu5aiEDHpwrrXIUuxlhabLC83R/+Jvp3t3bydI8Vb4aEogoQ
qjZx4LUHAopO0Ics6dxU3g13TCBKURperrYe49/9jTzPbELeiL6o8tcgl3ayDVOh
n5dBbvZqpBdCrVwof7SgBXIc3lUwikG7OUomjK4EeRRi+POrx5HMKJ2rspeVt3ub
NVWrbCN57Ma57WsPhCWH59iAy3oy46tDMIUpwTPfNm9He35+leeo7vfwR9a0ZcmZ
TdIYrTNw5H/Sr0uIBhhXMsm1YezpAXzrQEAT641GeGaNReB/8LFX58hH/4Ryz1qJ
MQF+LhigfNgmu+qi/snfXkUEhNO7jGLA8zXZbRLSH2RnYYqDPtDjThn0Iarorcq1
A1C/U2zDIL7LnpBnJPxfC37zt7EvLMp3zgC9mQT+H5Orhig9wXY6Kaiubx7volVV
mI8+swhPWjFX5pwRybpxBQ2zYlFaLDbr3Oh180hAIx/t3BUNZYJEXzxXXzBFzaiH
18u55NAF6/+Q8HXpGlOtVMGlJqDQ92kw/PkbBlGdbZA+mdjwyPmWhDd1IuFqYkRM
lXbedAs9/B/GLVfaPgenluJGL1cvttmEriuAd8AdBwqSFublUe1wKN0pNWcFnZy6
4Z+q0LNhRYKZ8BA00+vX4lzVd4TYmyJDwlzqZeegSAKfilPRkYfBI4O9aGuZwigL
cAYhq4aqpHqo7LHi7Za8CsiCyp9D5Qk/VNtENep74QikqAeIUW5JBqNtIEMEJC0G
l/vwCxZcB/cWjmZMz2GjBrTeivRCF8oZwa364cPfm6rIjSHLVKT4C/CGgl4Qiugd
CtYS2M5u1I6AjXBjRbYZUF7n8zVwm9mmzpiCvAx9VFFodpep9Y8ocuag0MQ4BG5U
RxDpP8P0/cBHrXd1xeKmxSq5pLN6rKk3989t0u+LWyl85NxL5TrACmcLFmN7TEYo
++CFxcQLS+GE7BrrjguthB8oyhqCie1Mk1it0HJ/QE1gR9ZDNfkCS2hfrpscuqkj
3jHrSh+Gp30KP6Y1DSWkDqSSnWzHHqUpdY5HgFG2pZbHE+mK0IXgQKVtJXc7a1j4
hihrtvmQ2ZwcN37mah5iCvp9veJ8IIyqiTrMW88hk/N+/PD3xfFYlnW0QAqkBhzR
sTSmVygT5RBRb43xex3UKH9U8RGL1rrODw1V7zCcFkPC6fR20IBt/oMmG0/L7Ojf
mNbymig9RGbcu8gaiOM2IRN9I8eJDCNzL2UgMvGlVppEKIHPyRg+/bfIwM3MOUXY
MYQ5Vlm6++FRIVQWyFZAdbmzGrn+2oyxUr4Nc8LmmYm7iax6pbpa9/+hwXLCiiRy
1qIe8rNwrWsSP9JLI1JnUW4ijMurwZyohyiKtYXlVpp7H36tQ4rxdCZJX2UQoqhg
kt/8j+mQs0lvDgFBRa/wnkCdpDlOwTHHcibDekI4Vpy0Zk22PClx7vGuTM5LJc6c
i4DLx6sxB3211/caU2aLudlDHFSH/JagC38Ol1J/1i+uOWBbrVYu21uWaWf4rxDV
QbkdL6utu24wxGSgMoRc5wJvmnr3qXajN0OxKtlqN4bHDLvoX/qEEV8pmqpXTToe
Rc+aXYvQZ39p8wqCGyI/U9lGSj/nV3WVoZUFYF/5Pw5Hj/VNC+Ip1mojWBQZshv4
r/bdXa9zV91aeTf6VfIf0fl5cDtbsqxNbHycOh0FoJyKKiJoXwhaH4qX/6Urqaj8
otDajxZOZohcQseAznVdJHXO0rnGTri8GML5V1AoZPqltJYa7wVS+sxDW6i8ulOh
kl7mxFEg4u2q8LE9NSvoCETLhzpewb1/lAWlKKJLi3dFiRGyOPF9WDvffa3t5nWi
up1qJNvuthkPJfI2Fo2KC45JwjS6hL+eJPu4kjFuZmFpanZEIuKci3HGXUbI0jeW
rtEjxxppF0PIZOrcEd2rsTcEl1NWVDdAxgOPYbOVvoWhb5AHgK0AqYSdAlmGvENf
OOnhyX7Uvuq/4zSG8cGtNQPD+tGJGzuRtj0Z0hUORBNTmX463l9mJLJqYg2blrvo
/JMSPxRZpOEO9HnPi9YXCxXkPdWHnFkNXxYbWWIUZ5WSsRfaCEyE1icUB2tsh4GS
OGBCyoafWgXANzze4VgIACygi7Lf7iEftmOUYTlx8bWcp+ctXUPJtKiHkpYdtk9Q
zgzFc9WPq8WvnZ8S3jcLtSXiXH5oHrcJ7l0TbZEkvylHx1BHnKo/e37cYKfo4oal
9mW2QY2twCWypXw/SuggpeS5N8jfV+NHaYu+HgjQHR1WV5gZT+DHta2ApHv/iQA2
5QncTRVcCSTBEad7ej3QmXqh5ASnAz9IlmpVKWmoSOGxFxi2YZdVhCZk8WbgQLyL
moB0WTD4+X2k/VGvomxXQt0SWrArxyIMIY9xJ3pBFGGcERh53LQjdJcOfepw+oT6
1xsxVU5etVydBD/B3CQoS86QrTP9cGv2ImCoE46BFdJpQxmrgylSbkLIzEBrH8nh
R3FNDrC7NWL8+CpIejaelCuo0bB6pkTGEVbLlGGDGSMFYw6lsLl3GvhWFt+bX34f
58+ePS4UqWn7Hx0LzqkSgmvCvyO46FSKQyuo3sv7LKH5qtwLzTCgOjWxZV8RAc5e
w5mUSHz8IDtUFi3/C4EAZmLIik2wqf4BV48qhZps7fPvC26Hnj30rzBJK7PG6Rzz
ZUR8/kFjU0MwGUu2r3V5hcZBRFcpCeiuibjjos+tCXNK1AgsHWDzrtP751r8y5YD
IO0O2Tkze7ZO76WZzq17CZzGXHiRnQRpcWe2V0LQ9mbWkb8d4uLB/21fSnz4sghD
BbCHFtMejit4gMFOe9orywgq13Y97t6W122TQb3IspvP9bPWWsk8b5QePEK3xBIT
yp5l/61/RA4CpDUlwuqMC0CagctDdNnXq0uYRV5TOv4cKFCTQ+AG70/3eJyKqRQJ
VeVpfK3IjFjg11LFzFv3cCrkuaY5vo8sNEQ2+UdSnNU7O63vqi3UATJ2xESodNiw
7BN1AUyK52CWn3QE4u5BaKSQTOjFlsLp+3EpjpKCMdMugmjt8lie75HEesQMml6j
7TS2Bkx2dvQFYnUWRAmfbViwhfG2V5uurYze0VSaj9TrNEG7z8DfY4m4M3QODLVg
2RT+Oxgm61zm04WARmddbThMUxGo4K7OLTH0LDPcO2FiNlyOlGO9UReG0SS+0rG5
NHp64MZNp8Qxs4gqJ7CIKlvl60I/fXjYrf8TMqNoQ+BPT7JaLnkIBJZ5VkLew3X5
0l0FISXdgbSqMeVsN7aVNkVKjImXoG+XZrfpWI3GwUTi2V/NKbeErpKms8uJiMsR
/pm9kYDgQYDYqaM1ckNhuINkOPMYSvEhacpGcBqDTSqRdjghW40kRBItC7ZweR8U
c6l7GMoxy6zNP0iIaAM9AMMxwvCcqSDW801r60+QW4sipWFB0kHWhWrdt7sTkeyf
uAIT3iDtuX+1ZO9h4C7w0bCXJu82sQnVEA6QzLbMVHqSLZ48VQb5mPUiTg/nobq6
ur3jiFgP9uwBPO5Vr/pcrXpyl0qyjLVy+0fiZdTgZnZ0baXlXflv1uRyjj4crerU
NHzOebyvHfEQQ0FRoWaMgc/6DvzTdaxJAwePYnre6AOhsCueJP6lZVZXORvGKFAa
Tc5EySt3g+zjCIKdTpDxbH739PBhQT9OhgXBq9kJs6SNBgbpsxL8hL8q14tiUSje
sPfw798r0LWwu8G2PxYv2TEbdQi/+C2iALgPAzPo6I4aBpT7Jr0FhW2lIY90n7yM
934zsmRe2to+ll2rhooVmQdTkvjBU69FLlaZumGxs11JbRZMnGVlHRMFQA7aw9Uk
VdeT5AYsDUGNSiPY1ymFtMhl5FGKmYYAbVZCf6kIGg5RiNupXY/HVHwcy+r64E1M
sweRgpLOhPu1jbb/R+Ze5W8XV+BLez4NYlxF2kbBbyoNTjaWITIrYVvQ+jmYUndP
nWD4Tb+j3OeugKLgnYAJAbqs68O0Zo2RzoGfA38VaKgsO2g/MEgEuRlgvF4vgueB
mAxamUP32v1cPoDMy4G17mLDCpq6K/UFAtODJrHrLckTTkHT0Q/OMH4ooL6w1j7B
hnpWPaTmrQgO+6oIl/QbF0RXB0yan9MpA/gDqxWAdNO88BiqqOtEY9bjN4D1gsj2
bfgS3itcjJhJoCguHsoV+xpR65fPiKEYB6+tL+lLu0DsWrJue6UeUhS7vY6/iZQs
+OG0yQx0RwRjWZNWgAh3DfO5ReVt3z3gSxw+EVL/1ts26xy1FYn1yAFY+tVakbrH
aSc/9OFY1AbgwfviSTiQmmpAUaMrMuU+RGEoFjvC17jNxZpKBgXDcXCOs/V5w4ek
CU95W7z0BegCtYsciQ3x4G95o/0XP/QxK/8xU06+xdu2AA2PO0nsuuiUskxHtuBW
cyhsj0fyFo8PCOPqAx7s00EIlnhAEiTwOwlN8ZCUX/ss71SjhcWx6HumPlcN6wWL
Z6X36ja+h7DE8BDRZNg6oIfO7eQvAEboqRGlCwIthM0bJUGT5ifPOjpphYchOw8L
CgdwgGnLEMB2AraYudVwmC7SEq1pLJsDKKLwr9a1WbhugO2vFBRozniqZfCyjYBj
3IdCNkObMxWWXnW9tWDLwTJO6QpT8sdI057E2A8nhh+hPAsssJin6jYBYpG9AuWA
NxvrsgePDt6Kf8z6vXfjuioJ1Ril8RGRYNEsrYCkMR6uV4evYozOytH/GKIYolCT
9EFC6R+Sw70u2Oguym0Ht61D0rtwALMKFNI/96aJKiK1BeeRqQ2zE7AqBG0nNh0H
c1Kdyt61Qv00M3jwI5EDwA76Gzes3nlvXzESwBVqWWkeFYaYjuL8CPfGQznto5QN
3aHMrNGaU1OCn+3EV0tewh/nv6y9ZS5WZrcXMJ7f/UeDhRCSfcu4CsgzrddXtMRv
pEnqq+O5YSEZXoQ7gRHAM08MRBtEpt+jL1COyRPUDzvxRX6+sXYsjGVQZS9nXd2H
YzVytW8W8LyxBdU5GIJIFivFRce6LUPQQvWnIQsHkAx8ePfSzwPjzt0G+X/sk0EJ
YaFNAmy/SyQHK2m/OSzmmF3jULHEvIcYkNCEJ1ImEVqmU+75VmUw/Tn8FatIwUss
qbIRFsZcXLL3CG01u/OTgpJCODbyEl39HwVGFDz6aq1GjjLh41ZnraSpniqBc5o3
eHVkkM/76lVV4AW4WFtCP9HN599r5LueV0rGZRn1pDTL3kfuUm3XfegETxV/lGvO
Zo/3/SC5ArDdtwKd+SaCCNegu9dugqD791AqWcNz+2LjwI8p6DeRbfrxJCo8QqKP
ViEj9Q6x1CFTRQE2nNhn4RpNR3rBRhPq0EoaT+LigxmL0CU083MjlfStyzpJLi5r
XDj7iUsvAXHgbO0/l5Uj4EHm2+rWX0gvpar5MloWHezbfuWwev1FxVYGh3v4UY9f
YuKx1Bpz+AfM+UlK8NQvbGExTZFDlZDq6rOZ+oeXoRRAbrIcdda7bNNyJztKTXBb
Q0nd/Ar42PHQBy63Dd4ZGNMT0wTQdbg8zu9QX4yWu4l/x3qJPgC/MMnAbZrMFdix
Io4syYNXPaUKvMCAWw6lDAQrMdNJsoZLb9jTvopLawgKuaGUY7ut1K6JII6adtyS
nzDXveMMif/ZJL5hKlW2roiZzn1o2eKCwy8PlZB+kj+nL1hdr8g/Dzc7uIiR1CEc
vbqcI/2nG6cggk7FPBBSDQLzvl+jUtVhEk4HAcHg6A4GJOw8NFjzoKXM6TA9yrND
O8a6BW12Gmvxx/c4ekhDNNbBUUgDWMCfEq69mOYn9vOaQs7aqs3gtktoL08hwQ7C
Arj7iNZ6sYXRgubTmSAQumMu94FidXgBZr9h5p4jkJbMQo4CN/FN4QDA7YMVUlJH
Yar02LzuHXFzPkxwdROqo1xC61KWSVoT2liDjDLYshv11tsyitf6bA/AFU2JOEGY
XDngmfu9gN6Ov7dnNc3wJMp7rcjVtD0OkCkNv7shviBjx4h7G6FKLYNKaLKVaoU9
zigP3aV9IphNkjSeI61sYSRP2Ja227cr5OKi0j8fArS9/nBFAtnYYaS7yhlTPy0Y
0vV3Z6iAWoCf4fd820zSW8vCDj+H5oKnR61CdnE5RVCTGt0WSQjpR+u8VMdxZkNh
cwtD952rTjeqDBAt5ZJjgsz+i+vErgk6rgl4whwZvHL2RrMKwt2E6NyZLWNzufKW
ftdCrlx90EKdhmIHvUqj94PUa8GKdkVaSKTwXqTnJF3dyMP4A1KP/crVrDXwETlH
JCB07+o1s6db+ZD55QuGC2+YbE85FRejJUHu3MMTbsFGGt18cAzKMdBs8ft0XmTL
AumlSgp8TOhLs2CCLmAdheWFD/iD5a2+BKocPV6AM/dO/n7MYlNc+PqhXsOsGmMF
8PYrI1Q8gTjUym7KVzzqnkoDV1+jXaTfwDOzBSQTTCd8u3N+Uu+yFxUEBZAuFUBn
DCAM/lo6EEI74T2FFmI0tVBHtdiKIXit5gdwualpGs2/lV8W4OMFJxDMascFQqVN
d2WfuVV2H7yC5ofQzYzh2E1XyRY1ulkFCLhsfCE6skFCjAinrZTAk0OFTEPx2bUJ
q6jrWC21aHyRPtthRy0+aj32ON1JcM0y2f+n9ipcwmLkuQ8GIouasy7wWFWY3ziZ
yu+aqMaDbOqANaYwR+EhZFAPxDOahvyaHJlC4NnGoDPmjHDv+335azjGSlqWeqxQ
ayfdVc8jTkLqWxoHqczZV7zJhUShSh9+5ZiDRFEDKSK/W1lvXmhf2AJ8UVkMigOi
4ezxYIP9J1eP1WS+dzs2di8iWuF2KutrzEi8eHIAAXGgGpi5cLN3WKO2Ym45Pkby
fvovH4hJLMu+zkcqFpvEb83hZqaji1q5WCMAl2QaExjeyg2sADXVYZOwVL21qkPE
cHqdt+Q95RJZR/+SzGGvQMuE6tShB9+yqE0Q7E1fxD7IumdA+hvrIvixS9Befx7k
E/F7tagZ0cmYqlRFZCf03vtqYj9DeYaw1n/A5+YRcX9zfXxHtg7wVZ7IMZu0mjzA
Iv+T9kxd+Qx9cVO3hnPEjs5wphtV2as9wwBbr+C9Ir0M7OFjLf+KRAafcE0dK5Yq
ZJTAkZj+BOteTojzP5h9DaZCUjSlyY2VFvbNvKJkrveteHmsw/smne67WO8SPTiL
cMT1HKdHwiv+GjmCJ095B/X8vbXmVXFZYfCgzo3CCYEIwwkBmC32aLr1vS4rZZR/
9G17FNPa0LgyWmgOROnDaJORI9DDvlaI6+NdcfL05ehiDLZjlA8P3L/zMcLrM3nV
i6bYDgt9p0JQnbO8sbhLJqfXs31QKje7XPrJIRZq59TUAgZD0UFz9sexhq9soobp
XNm1W+nHUbhOGFBLgxpETbN37Xlen+/1khhTu0ZqPI34vxI6xt148KDOCRJF6KrO
VP3mVNwZqaOqb9Za6fahU5FuhcMzw7S3eszsdBmIB3MARX7FDdO36DymH+a05x9W
9NstuLxKZGmsMX24vJ1t6Asjub1ozirWPlrWI7c6gjjZGKP2NZs0wNoX525H71cs
LCB4yUTIzLA/p8t4AWKtYFu0sLDnF7mIkYWL0JkPZ3NPuaKZmIB5f+StyyBBzEis
H7SuH6TFEVcEOZfzh+x8hJiBI2qJjkqZ4IWCUL7+joDmaJchX/vQeZqOc7hHUcIi
PI3rWrF83GvI1/UVrmq4qy0WywSV7CDnNRzCUbVNPaKvNVNoNZquCToTh42yKMCV
Jp747Doy0eUlreHQn3HR4YkMVnVToT7XTl8WjOJtjDBcrvHxCcRXpSjcxmeyNWgZ
ILNA6lZRIuvE4JHZW+L3yGtjoOcD3sTdOkiX04hZdSBGql08/UQidd97ML3XZKJO
wxGcCOGpD4+OaWhbJmVkNGMPnH7GL8AR2pcE9Pkm5FBAfzHmd8GODHUoj8WIjlXf
D1yR5M/G5vocoarScBmahDdJOJwQ1xLVmm734XZi8nqAfz0BxR7b6PLU2OhHXWE0
19cLUj1NAnSUoQE2eqGy7oWJCYEBtEscSadafFvLFzvJI8JsusFn9uPRjflKMnuE
19qsgTAJyEtvvaAkDPd2ZCWHV39MzwyR/kU26k4XshWFo4Ri+ChP+fCUwcFscMtS
ZAB2T8BOIcPAxqa7aHJR/CdGUfefLCPZNwCtyeceOHXkZOYDv3g/pANulfpYAD3R
KQlBJBUv1hwmzbW6wZCJWfJutaOJJK3uKhoMRmqr0dKR23Pveu8v/yH76IQC0OB8
QxzU446KByvpr9ng7qT9zpeaW6fjdFGwrxjLuIAUFOKyj3FDNhQ8LCfmTzgaGxyu
3FsF5m8GO875bW1UvGqca5Gw26xsC0g8gIwa5GG5/POao74E2uo9Q5rYbkfJ+/OZ
V1QtiN2Zn7BFj6N7sHrkvxbnAWGIJNtLDPs/VyJlvWSfhB+WaTrNfDr7zFmilEk/
bwuI3jPOugmBw1spkB+e4CC6qoPrLb315iaaWkwu5ErYGR1JitZS7wRptybwGqS1
ugITdisu65YurVyKSEkA9YJ98Fzav523OGg7VdHr4aq9oRbufPJw1100aEw08Og8
pvC/w08HlSfypOYpNgv4GfHFsZWn3CplmWkDJNvlYHEPsiEcUNLD/k5X1P5/w2Ke
L9/yV/4kWzL/QDl+DPxHCR1G+pLrrdP/KvjzeFv5xHDWNJ00BysfAhK6maIqVf0P
aC29QC/vATd2ZfrYN47EiYmG/sDwSYMj3BHGPEJdX5kDs2r6fbNU3zsxDbX7apui
lZ6ylGP6RERkZ0ROCJLs2oQiWo/pV5gXJXbsgAaeq3yAjPNZsus7xt5ZngFjT8OZ
qXtf3gZeVoCLj9WBM+FkwxCFQDik9ms0WbLc/Zb1X9bo+qi1HNa3hAnIZWIfnjnz
fl2XUe6w4rCet5RkRSFL6cnTRdTMhXZZeTEJgM1rPeHJSEd1rr71G1Fc669MpZoH
0J8GVgU3JjfPDL5+6GjOhH97xWjQaXZMCjLDJ/spnYwJZ1hlJKeEwSa9x1gdKvzq
NY6QNjG67I1sTPrlIHuKmJngrkCmKGducQU9/iajJKxsNIv0VIKVVrCMxqPXWsEz
NPrdS8A0MbMsVCSgNUdOTRBApYl6FBJW52SkcAYjk2/fyLc3+JpoZxhc1l8RVMr2
M9z1cQv1FuWyc7tDzQP+WgLSX6HLcosu3AMiIVkQzJREHNti831g0cK1dF548fzl
Jo+5DhwiEBx2VjOkFzz4cAdGj1PpPa5/D5dnUlZaxEnFqsQVP1jZzwwB0t+tJE1o
Dt/1FEyrYFtg+3eX0UrGkAsymATACtm0K62vfshl/5+2vpdIo+8kQQpNC3R+Wx0c
hJ/HcclznkyFMPOcgh+nhHa3HNJy439LLsspk3EBokrNHiSyBzHu050DUU8CzSXw
hE9f7uDplerH9JAangBCB66Rh1qxdBclfFoWIUy3oU/Hb7PjpKfvQaTONEYs5teq
otdeNW82dAQ4v3901DD3f55RdRxYRBIc6EETMPy9tdDQhNOsxWw/67OH7t0UblMa
/EMT5aJ19GYRJRDm+5qEdH+zhan1D4rnF7Hkfr3DglM1lM6gIf7WPtXvmonYfkEx
GcYGTCLHB1KyQ6+nepHXsMV1DQy5CzPahrREQ1hBYYSjbn8MitldGhQoQrkskTn9
qhbvoWdT+OuK/UZ9rLHnKFd/jgIzNZg8cL1u/j93eq7fOXLU4izk15NeuXa9F4N+
NPQI+F2/YnL43q3zmkbxxrgsQUbXdJ03LBznmzL84YlANWUBaWeuYN2bTG4XO3ow
VLc9yVqZFUVccZM/s5tBwNDIqGkmZqurPVZgiEYjldkQOgnh0L713/KDHkIIo1U9
yFen4pCyH/j4yPLuQFdrIpmyJO3xAOXtP/EvoZIrfSrvxyWRwqLAwXdAiBH7RoJS
J0/wdb9wa8QtYNWavc5YWPHBGF8GrSE0/Nq6hktRRkbGufm1/vuZCcKFCIDMDwM1
+AFwadBFGDRnp36zepI8qB2Jip8Ndp1oDBxInMt85JGv4Dk2S5Bcpk9TlS4pI3aF
qyFwJVlLmJg87PVGHTmUGVaOQVan4KCr/ea7j3ld4LWwAUghhWQfuDATu3xLF6BO
gRojwzS0oXRGlLiuW5+DGpwptajEJUhr11U0u+3qgS1crq/Zk2l9zOmsBlSI1xxC
wOa4Yft7gqS4o4GgyGNW/qZQdqLsauvbi5k1ZqVYh7X+0KhBCeIpMcl/E5prB+7X
fLjsEte6Ib0aH/lC2ScyDcfDMUnfXUXdLAvCd46rn75RiuoXUQyOA4L2IAnM6Wy2
sWRA3CRFuu9sqnHV9bsPpljEIEWDZXpN7dAeEU6mPt/GCsEvIl0Ddjsag113tqkj
IV+m2cGLWdn1zcTBkBjDg1nUI3hNfy4n5WKMVCFg9YWn7LCbzklTBjQmGyFdgFlM
5RroEMeqDeSK0BNkVyg6UcbBnmad4VITK2uY/v2Ysyz83wNuWJzzDKe1KIWexMZz
AyI7TUP6bdO0SApLRvE1xz8ZtOxEbkQZtqddiLv8Z9UsOILl5x/6+BdhSfpKsA0S
wBgtzitwAMm2hnzHnRpn5LhWnAsowhVcd3IME3/8pGBegGbafVfYKveYZf1ITWJf
ZU//JzMbZbP9VVPJsjFDjkrVMpcFDGr+kVLIFFYwiny8OwJ2oocE2xjTWaY+tCA0
HaxGoS6PEuI7NNr/x+ln08sA1x8v3b2AaBOjoSZvWH+wrSmR9dJH+UD4wi5t/3dj
z2tglAXpLBE8MrzXzo8ZEdPHjr6frcF+hA9W4Xei2+ScDEb4P5WMuJIkeku2yl4B
+ME3Ar05uYHhpH1KaGzr8mF/AhubsuO5ygRN/EmBalSn6+AEyVlkhkL9yq8/1ZoM
1b78mNwFsvHlZQ+UXqPoN08kdKvE4uDtHiKxMuZqS03BqVYGBgpO/0qOy+wUoqAg
bxNCF1oZRtZYzeIsmUQu6rgA3Z+6OpwWe3NCySS88YYa3xLRTiHgmkk5jmhVDM2+
t5ZUBxJynuwmXB3D2ziU4Pa63so/LuGDX6L1z7UvNkl/wVjeTTTZiYGRNu/ddPOi
Yh18dEXm6S2VZvqUBHJLISA1rEt5gV76ylBbOYsogdBZvtFnbDRoV21gQQMMnmnM
3bAQPGVAPdgGGXYejLGB7BVXQKedOsERqco9LBYHCOJCSZurgBgcHA4QutVMnWA7
tIQ2uJHEL0z1iGzEjwATX6P3EN8f6sHBhyaL7aQTsbYg/kC8kC5rnpeoMi5rpOLG
9gHPfQKrDQ0ljYw3l+qnnya9PuPB7+AnMNJcuW2MHD1OCjktQG71Rqb+2V3ANQS/
PdMqOEhHtbCyUnBgxxKEtTSdJtxgX08EJxXdPCIHX+yiwYb2zMO9kBT8Fz5qhUqA
PbgRWGOz+1f3VahYqBex9FZGixypEGZzn/R682laywzncTCWfBc/jVRJhoyZ/wU3
xPI72j17jYcRLW5bSBgiFysSgkVep4hk535ASA5vrsILBd+m2uptstux3MKyhIlY
Lj9svAZzWRepJCvCpUEQ3jxsYbEibdsEAT22Z18uFGA8tjaJGQf8bxLMg0CxmOeM
7/mUtmYODyvdnvHnX5XHfkt26t7l5utJH3t3lkoY2S7rQhXsen81aZnj8wn4AvUV
vv0iAdk8doiSa5ED8GfcCsDX+V2js1d40LTD+CojNoehafdvlXqYu9WH5wUYGl27
tCtrvp4Tqa7TYIpi18CuR/sNcuSj/v5dIzFeZZP6VLpTREdrHQjCLodqPSM6wvOx
2gJZq+ADSLqlcrlpxChVhRlB+YcCNHauUIEXTWVUvB3Zqvjralh68PFdmhhHw/7A
ajHZwhQsw0palkPeNSYs/HibYvhMoTyOTn+J885y0AaD5LfXsDE1LGFgI9h3UTQ3
Cx68rM01/iIPfuTtRl/dPMd7wrI5626is7bosC69DuKS7BMZE1cO1M6/ZYx8u3K+
alt8mNlGYe44fxVtZw8k9oWUTQkZALS1oAQtz3o58NZ/U9N1bSYNvTalrnm5Cl2T
ht38d552yKhZNAoXim3KQba7m/bq+PHjgxAkvbKpanI8yNvnte5WPxoth/btB417
f7P8+cKn1F/ciiVRAFFEmpRh7EG12DPNg/sFl2f1CkFANTgTvt7+p2iIoJeBiJQ5
c1MmZHKr1Xl/W4AKZfvvUmULyqmmpxxYXd1my9V2wIQF2ifFxiCL4/mhsuy35MXo
RXTB/i3SXSVLUTZr4K9ocrlvkwipuVxo9sNNrL4kedHqW/4h8tQTVQoBowPY6CkW
75Vpw3dmTm4tmZC60d/pT1Kxt8ixWGkV39vPR0pb3AyG1j+Rsu+RqO43sr5VJ1GT
U0rkmsnamtoR2LGdd2yjwLUA3NosEFfThmdBbw/e90MHFWUuzQQmDsDOg0VUDYWW
4FnDKSyvuFvei+MmxPo9nJ5uiB6PThjl/i6PHMzpsTOuVxP/rg2g42TZ+vURlVb/
o04YiPbOs7ltVdoUGr9vnwa1t8ygZWsDuzcIwI4m/gQx86/rd8piqXRMYUop7awp
F/JK+eETn40GhedbGLtwshVT/fgUVhjd+PgKl2DfJ3g7taDAp9hfRu4OtPsjcRHi
gI1AuLx1WIEZGH+umMHwJr1Oo9aimmtIwQ2T0bwq3cgI27EoFatoT6B80/Zuza24
GmY6pzHCjM0G2XEYiy7//E19ntVQXUWhaR558kAfysTy01oCTUCZpeDrf/nIA265
ph7XVfCTfm/5YIRT/VFTGR5zaOR8bCW1Ubs5uU8otr8RZXOkjkzbL+9U4Y+L06D5
qEJ4hGudy6qoKSU4O3CWd2UDk749nJ8JfvrjvlV/rwPpkpCKYt+3HZcqpgZawsCq
CmCp1HK2hraEn5kUV5UDWyGGhEUk2INI35UDOaV8xL1oK6THyCUuSKbjimHptZNw
zFuoMZ2U97rPLC6QkWG4frV/rGhim3oumRq2kzBrbNPzc0iILeU/X2VZdAp0tuHh
Flkas5hHhUbNdZf4I47XWQ56nb/h7VjEnOIe6am62zsi27JE7VQ2NvOTck63QUTD
+QOYnzU94GrdsEoE8858XADjPUWCenJEdOx9JncWAfXsd73H2yThLiauzNogRKDI
RZmkz8P8QfiNhOirdwc0tfjNSHkJLvAjSR7FvXyc1z2fPBjmrnGhVZdt1ABGzamz
Zd2FdtF+Vst3AYIRMmvIKCh7VFKA+Z2WG0dubFG7A4+M1Dt8EpSI4iq0MJ9QmkCh
NT3ZRhj2tN+fDFqSxCXIITFMT0Cg7tyeh+AbtaPGGGvzuj8CY7raNKDS3XWAsN+E
6TdEf2sT/XiM36agrf0cnUEF3nTJoYAK+kjOSOj4TUeI92BId2S+rUl0tN1zn/KZ
qnuqyWfvZOyPLxnIHu+CwSm9t2CmdnE1LD1c4aquBRl/GfNZrfWVT3vVWOYHAZpP
MDCPfnMwVOUqMucZhPVDpe06s6kZ4g1Bgvyb6XLj5U9+wJ3vhqdMrT0g16ddhyQB
b3iM6TCEWEHpCw6Yum++csgRMKVyH/pm0ZuY08bqtHoo3+Ja5lAfL293jf8S/Smn
TapQmvVOwsrPHWQdP0F+mOwUFzAJzyZAZ/DD441BSqlJLBtzxu5SEfVBFk+Qw3H4
RUV6KL9xNbhJrXJAUZzVS0JTKVd+6L3/sL6w2zoTuSZTWd+yj1F8SAGpeQjP+aQO
/QWPrZowUzWgX+QvFicV8P1qIBNw87Z4+YweZwGBaYa/5w/CHok6uaDfV2hbwj5p
Ndw3sywlxy30+8698R+m3TBZAdqADCoI85UI6VIZZUFJh6M6ps3Xfic7OfDPOkh9
mwGj5xlny+S+K8oVppQaZXMrk/LgFIpf0YrUALCQy8/cmU7xJYR4i9PJPmtRoxwd
NL0hnzqS0G7+WjbW7JFBsbokMM3php8aBz7vznQHHTctSkhJQdRQSwc9nxMVjn0B
nRb4rsZLRQ7xSQvuB6JvEchhtGfRvTl1R/BQfZIUAaT2FvSNzlLkMS87rI1UDFbs
Tn8QXnd/Kr/oKPauKMNcmF81lKbgjKuuyLc0HWGwyc9ObGfNni70sCiX3RbWJuZs
LMCYFIPebuAjpOK7cGNwpC7BLk+WZ56sY/k6dK/c8B8A/Kl3w58DGWbWjQHx6WI0
dWauddDuyHMqqm6gfHO1eX8qTOLtQij7ifZTSCOPyYSiQy4Yza7o+dAWSK50T0Dx
W8pyBnfBjVGx7OzJ0d558BNpXkv7C8sAUx5xJSOfhZgxSclxed3vHhJRjAGQ7dXu
N/8Kh2cdswWQQVX3ncGJChPaNyAp8zV1opGDf2O59BhlXEMvp4UZg15cxxzASpZd
zJMg0FG2l4WMOA+aCDWRYNiPJ0FJw/0aj89e5VjOyAPZ/KB9NBJr9jdfC9S4VUF1
M+1MyUR2nG3lU0WOeLrP4Iu/7FIbft8s+SzVuTHq/SlX0gcR5jdrg+BKIvRCXIEj
8Ts+J9Blb7UaHqIlbY/7IN0bcs+hKb4xhnyWcYG7Lpbrhys8L/KePkK/J7CFVDFU
h8TEcYJo8vmGTtqeXh5xUJcCDglVnegHxU5JdqfrbLM9x/n6uHwzfof8UxLg2EbX
dxLXwgV+Dy2wgiI9JAcc90ebiwI3pvmYlJRNeJKPnjc/ce1Du9A3RlLpIGWsQRLa
pWbSop0bcjP9yyyla2F7fSQY+AfaMTdQAZ/6HlsyG31ARqt3tXSbotgaVTkQU7dk
syXv8fAOP0z02YYeSYt0iA7EKYOfaa2Dg6+79BajdXdVOwxYdsushn7dCYURnjXZ
NFrY7WV4FG9wE7gynBrpn33D42c+PKuRDTAjafrIdsU8kqXgCIILJkfhcwLpihJq
04JQQsetZ6Aw5+RmXhEo0mgSmkQc5KxuWkp2trD2oSIKd98110CgieWASnHoBCi7
48t/dya2O7lezT5KmK9Dk3PuuCUy+h9I12oS3UxD/Srkb9cTIP+Jg44lx6cyzoli
DMZIm2XGWFOekq8cIVX4l4+/8GT1H/D4m29bwPbzqvCahQ2MPgOf7to9b1kgtdsy
ml+BfR8RZKPSoaQpVXNs9Ixss6RvO8AF90kIJeOb5poB9XygSxBmrgg9wqIXNlxp
7QaLRDmKtOamHeq8UCH+gHhaoxsgbX5Urmb/Z2Qeniezvogjh3gI+r/g5yhL1I/K
+V22im8NLsd022uWLM+OTzQ7NmIcg3L8sHRQki1AMDfT1tG76F3B9vwN1X08SIoE
lQIKCrsWW9s12wbYswTe09LdforfdvJN2e5H59MAvD1FP+h/OXo6+gVLkwfAG0k/
sqmlfBQ+GrdYwh4RkYfnQs+bLEQkn/wP0y+ZX8BzHc+JWJKeH/e5SNVHCNFWl3Vt
DB9O/zNC+65iSyvq8EmsVq4R0EmlY7HNH9BHdgYTiKPoFb38E6GFa8J5IOmj27jY
MZd86d/lgKkJzMRscon2DqE8f89Zig4y+iB3EolIwjeTPQp+HaZmKz9HJ/xsJGKd
Wvr1A29Y2mTuGANEBopOzdf1z97T7ACxsN/Y9iK2mGHPPsxT7Kv1P5tEBwGgyTHN
7aHQ1nnztKRR8O/yfUYAWYQaIimoRCVadsLp+iHQ0Jn7U8pMntwnVtteZSbuEBPS
oZ1yBhzTdKmrGdQoYW1rWDq0RWUMSKQSIMwKOhkZjSlcYAHGE/utpdTg+XaybUuJ
Z3jAt9ngXouX2fV7/fsKCqPM10lN7Y0bG5ylusNc/7/pINZQJLA5AWrVs8gSMtvJ
bxy/c2Jhl5vcUWASzJcCVGAEeA8z6kCNrylLB/8p4VjAr9s8wC4502VCGt7hAePA
WagV7mz5wFHojRT+qjjBNxn8R0D1/+7tvQbrFaLC++wBNFMNjIIsKvv/x8Dr1FK0
nbgYUlLxIFAQ/GmjTO8TxzioLaFheycAigC4mMD2Lua0CAFw2EXvUr5QQfgiEO6l
G9FCWWKEWo0bHdWfH7oTL6JLVzGV/qkBKyz1INA7KUZbNA9D7AVoORiA5v9QTACG
C8aRw4feCbrUAlgOYkZxLIjm2BvvdMjHGZQzHlqBOVz1W2TZp7HN0tn7wkPUBOEJ
0pXOJTYtqJVShpdXiF39n2Jd9c6B39Eq6PPPitoM3U8eaWfssqlmbnuSiD2hMHfi
/+yTITCPFClYGsVldxZ7Ci2Utrtxz55A0OEvlDdPkXZHj48fy19dM9cHD8NytsIz
4dynhZpqAouimNF7+w+hxe3URkSDlfE0xSq7raeRbCsd/j/OrYdIQSPuq/XzwyHC
4ICSnHoV7h+WZxlqWsM62DtHbyJKfoZ4qXfklsQqzNQv9z8Uej8qhV9cpoeU2Efv
HteqxjzUb10zafFFDPy05aHGTWGdAYz/POGtc3Rt+W+0LDqHXxn2irLADQp4uBOH
CNHvudyul6qyWj14IhvA4JDKGWWV8RJkDm0ci68MOicuau9swjGYk01D/wKd2p4V
Ua+WNiGQt3IFceHzKsmSz0tgphYcPQZ6NulFCtK7k/UBE50qivDEHcK3mqKNNckU
tASYhS7PulCwgZoeTdvAkEacaHs7UtGS8Ee7gpPP5UZKq13flYR56jNzs83W5PI6
N0yJEPFhdZQWnUkxNGIJxWaSO+jn+YORAnB4nUV1YdBLFIIEfSU9ZrPLtK1kR5jU
oct9JXxgMyZCBdXyqEsLJfh2PVV5qrTNeiGCmPjWaC9FF6EUePJjcsAg+GKfTWjd
fUi4v9YFtS9A4qfrYSJKbea7U9agcN7Atyn++6mYzjQJYlOASF+UnF6EgMmSBi70
OYv2YTLVO8FShO/vGl5s6LaXL4DA5FmBZeeCi0WRhf/S8p2iod8tYIm6yyzX/1z7
O5wxei1rcuAZUt+GHtmSgO2bo729q0oO1rOP+ZpNmLVn6zYxXQV3YNFmzWiInDGP
JE7qZDyfifUvm77u+t0Q/mzn/BtXqjT8ekp7DKMwW+o3PPnvno5unGori32TqDf3
NUSsM4zgLzCyaH9f3p09370d+tKW/J1O/lqIliKlDLv/umA5LLOCGzyaNcY58ApN
8CvdQcuXYpYHA4CqDN+DYIVLRByZILYei2KKcvLvZNSacze4Fsw65lfeklGAjW+P
Ogvg809c3dxKTdBs8LcKB+8Z0NQAx9ozhMtR65fzJTy96FQvsFZiz9As6OxJTKwT
rJHbLE9NgtSKr6b2lhvoTU3j9t3QJ0d9h7uAOGS68SQi6O7g9xgy4PhO2omgFYhX
zjkekUWWkA+cCHUV2u5hadNykD6l1A8GkW365+qDjo044yWmhbV+lIRQH1cZlO3r
Qb0Zo8zynYPIBeWUv1NOaLQbqbXeKsqAh9Ylq1uWWJotiCmjWE7r60Q0lW7e9l9o
s3rOHK1h9g19Jd+oZf5+RQyvNLNrBrNgr87kcxmSvATow1au9VThFX3PHiVwfjl5
ZnRBj1m4mpDQ/IkLryVexRChzUechqfNRG9N3hyHwa3+mkYSc3E2PgwoEJm7Z1DG
ErN9jI7bjAp0yxYYmrMedTgeO8bzeJpRhhJjhAJQRUsA6r/5Tm8EOK1AKs2siLlw
YEAqYJujG2gGHAuUbzRjObsMVgumnJvAQv5lu+euO7czOG2UaGITVS/eYnYpwwtH
j8rNKUmUhPtODwsPtx18M6xtdW8APr44y73Jx/ZwhLVI2zyEkNhibGLjhg9AOpVG
wp3Mk7mwJ+XcYeqiOY83+ItRkyBtmmGc8LM3GaTNCeIhOkjCCTyIuxginJRZtSso
Ln8dGsgzg/wl7wMMrIbiEGqsttB81UG3wb+AmnPER3x0yI0xH7IA1fch/kYIGHi7
KUPMAyk6FdBKf2lLKvyygAqGPBwqTWh0sMoZBe8mTVEEve2I6V+plnLfzdgKH1XQ
l9tTIKgIzzaDUsnstuLFwuoTmPZYi23zXQ6ZVrnlTzL6kj3paMkcZkPY1WmIc60+
GiyvfcpqNFHlq3JnEQnzFRPmutHcV7RM5276dZ8/NRnFOhPT+xKlU00Dyt99Yqjr
2aPnm/dsWRM6a8MPSCqHzR9f/i2FtgTHvc111smfEUm+ZNjVkKxyox+QuNaxZkZz
28NjdceM56iJr2gcET4MEYPwsRrJxJGAZAxQHCemGPuE2SLGxDkEeE5Opv/yjCfI
tTjvr9gh94lrgE1z5jWvVazYbHYAFbZ1KGPHJmPMvutHj/kdY5M8RSzHLa0nMxwc
KsIWcPRkVq5EHE/3RN0QrbhoeWkq26wtdM2rZgty/1g43tZ7ebEtUUQ62FH66dqx
PLVMe17pr+MqYGkauQNppSXOYz1+JVLpuw9ZQcm41V1ltfIXPjTfukmimkUmwnnh
P5cVN92QPTFGdAVUcQeBaviERxcErcDVphGK91i+C08jRrphv3S0Vw2tpdt8x6wB
xLoPTquZ7CtWu5cUZ9KU7RNw049CVyLaTXDM+vcJxnto3wfz9sItghVqjsYZ6Ydb
pRFdi4/sqhERszC8cYkQEcHapUWahLiSCHT25rxH6lFrcH9wEfVxUO2HncCv5MRp
iXt8mAGKvjvaLVbnLfmnVaeMq0/uYJi2GJEM7n2RGtDBZgpIhE+pfzhDo6XUMgsW
OYV1Zt6RT/iRie/eyZsXtR1cTqPrkegTnjlHXJwoR7xF70c6q953pulAkj1baww9
2vcJ6iqrw5g80KUvSvTKsVf92mWfectUAhX0LZuRZCrWmfSTNcMnQRS+EFw6qzJr
wBKAC3luKrJTNLw/7FmB19LepYkRQlWopMDHrFGxuZw83+bedE1GAJQ1KqE5QsQB
ZbQaTzRS5sZp1OVzELOIS5LmiMjuFwPSPwLmDNZ/2xoiL4/iZ+q9LgBXgGYmYf5/
1TeA5Cim0fNj3Jmp7GUBBdhmGn/FnyXQuSmo4JZtGb0i4mq1/NaCLteXBfvYz7Mr
yBdILBA9rmA0g7zkBgBAq0pWV60hIaAbYSwrnYZ5IhiJN5x/LCQ3MY+1SWwPPpT5
WENBAI0d439UVM93mIeAy+2GnQlTRQWaZME0tjzzh7MWp7FzylW/GnbhFn8P/WEW
rA4ZTVKYjl5ztA2WHEUI0qBzHwiYUWVjEhkEFlQkcYRfF3TvgwgjZhMuJfY7a+UT
bCrozgzQ3dY+9Cn/ZE+NPlGiXgHB2JQUVFvB5WPUjHzzmo3AjYXy8Grb6+pbbsM1
2k519QllufGuhDJRtCMMNbaO6J6yUynstE6ntLKmpk3MPFfi1vWxv4xAHv70LfAg
aQmfqZUitXz+jgzwz4K4Px18d/EoBUtVpDpPYTIWBUHK4PTo1z/zUZnpk0Az4xYx
Xu+EfWlW5FRHF6QPLkyESCzxkM5/8kC5WN0kVipfOReWebyb4ApIFqiwxGCZ1qhy
mWBiBqmSblqGyAfNICegQ3DFLFZ2+yU+mijWzTf9Yn0lziVeOcA4uvlmh9dYdaom
0jPm/77+WZaVTsOz46ZvvW2gbQnj0LRYEiCrJhqHMAfOGfTZGjd2oPGJO8ki/Nzb
Ny3h5brZZdKagrdLbBrMmdIOCZeo90PY2ESN3Hh+ZaAXZU+E654GQZgrkIT8N4NE
1lv8HwRaSRztDLkGA+uMpM2NwThWhjqefO2EaL11Ms5XSOY6f9/BGTOpTRi5aO0Z
GOCPQ399+UjGsJbG5lT5kvALZapzodcEi5elXfIPRuGyV33uZGBnePmZEOdHHtMo
hIjrcy+jH4hbAF6HmK+7KXGjFk42dSwOFxLDYJsG7tRp1m4LC0lBhH88S54Owyk3
uGiCNtDZr/cmT8eoovy7wBu9BEqnF5aGq7DoYc4xyjSU3h8BuUHC3TkmW9QiwGHi
1QRWweh14ZHY5zrHWLVr1w2MM7W5nm899ZIK4lQ8p1TiegDYqBGlKhw6Z+IZn/Kt
5PJT4qp/yKeW21gIEPMtwKRYn+LquEPC9UzJr30SttVse9LCCOwTEUTCDMkmgQlM
iMDLRpQYa+JxQPJFrpImtOsgUNQ5Z3l3cqN+0e67/ffqJvSPoR3V575hgeJoU/kM
5zUe/qs2zlHtRLT6Fx+7whTOUVU4apLqsXtRNBYInNnn3Wc83D0RHTmoB87HY4vE
j62S/D1irtvi7DEM0g6xj9N0MXHWYoo3q/INxrkpk5MP86PNKtH2zB/6nW2lx04v
Mgc7ITYTzporSCOGOID0KgiKjwHaHX4Fbz53KoeLMR9LR8P9F8XEEouBCsG4NGGd
ACkOHb8JGyUPKC79lcdXlDC1jUh+YHSRY2L1ECjk4uKtF38OrIkcgiU+4zCIWeoR
0nWgAWW9QG+ULm+l7MP0vL4vSm7ZPbSm7xeDJBzoyTzaCsKnOY5Vy0Dj6RytWgii
7/iGCNUSsHMoOitN5JN6ye35+wafpBx99ei8xpAnPTk7FaDoMxHzFA8cNCkVbsop
Ak4tHv6Mquw9gSM8U7sEc4ufETVx88NwrDVx6nsfG9vL5ZTB4pyspdy4T2YIG4vQ
JuqsfvIF3knS1p1IDfjB417qI5JZsELtzRvB9Tcf4GLKi5G5RL9SZZTcJwBSHhZv
DDptYoa4LQtcogAyP2RTORCoJ5D1oHqjrrjIlGYSXgu0A4PlRQeVO21q3iDJfLmp
gtpCpvmmdAovv28q0A/MNRy1we2/FLJQXfU4QLgjT/Go0KVH8kSAH0OiozquTgMV
4Qq2XBC1XENnNK81SeqAmepPrLsmVHrlo07xBD4FaPUIAOM++hmgYtgsWZXivXxJ
D+pn/PIRBeeUpaSzmOQmf5vcJHvLb350A2LlsyutlP6DL1txxfBsQD6rjjgBwvNF
z3tSnIZjIyQDRJXn2tPHSoLct0eJpgFSVRRH4wCVpyruko2alhHc/xJM4pJbm75t
p7NS/RQ5/HXAD039b52OJK/eC11z7tPivEPM8Th6hoeZXMYOntzsbM2rRmhGWXVd
hSYAxnfVqLf3s5iL6Oe+160hv+KvS9Olj8RqrHUc4NxL9oK9L9TzwpEY2Dit8jVe
c98HMJr+K52mrHjcDb95HtcHF5XznEQ0VvO2l6Y7wV6gLd+M+N4muskA/rHn0MHj
6139LiQtdYtYfRox7JqWMPltliGmX0YDfCbANIgvoe3/AYQhocBb2hgZFZz82lNr
dSP6VN3IRkFDma8V5mWNZXIGhmDd4U/mvuCnRZubaE5VFTq/XPc9g7CJ77zh3kR7
xNbF9WhPemSig45LaqSuls/PmKJ9CL44cT5EiBx2NN7f4SYzVkR0w7Rffw764wdc
YPZzOnkeVhfdi1G52OYhKQtpWYggbv11rpj7l2+M8d3WKBDXqhqB351p54eWmaA1
TJfQRizduiklvaASS9rh3B9sgzmboRI5s8rhTGuOBc5+PRqOriYkEUb7oQ09tzSv
zPcw/1YjMnn6eFSfh2SY4c27cnwCgcK17TRSu8+Qb+wEemawWI+m/OpR73flLHzz
4JV7hoKr8bJkwQ02ZvYhnhKEzvPzMrTJ9SIMqf50C8LHvxi1W9FSRLdL2Nh+bL6e
93LoshCTMmiDYuEu/5MqYdBHu//6BpBc9i7+aX1kW+mT9Ov5yUg07cFXv4oZqg0U
0BbX8GqrK6rYRRizmozqUr+/4I4se9H7DEJoH8U7jXUzp9r1jFl7EKaK9xVKVavo
rzIM8zzMOxsX43HtMTLwoutlIjx+ztnsKQz5+FYAhcf/3kbqLAIqpBA9ChRbZLQM
1c5H6C/IO1v5/caesHYQcDSajuJrp76kjjEd6g9NqO7daRHvTllcBESMlxT4GBkD
Ov+Mef1txWYjkzUdK/5xXQuAwtLHlJSjt+51sBqmlC8pqVgqvEfogA0Zr04fIj3+
v2n6lVBCzBl+zPYjX7Sb3SGMKUrCwZPxknKCZQMXvqme/Lg6dn0gSkR4SKs8UcXs
LLGrvcQd34oBnCBHvrnenIt+qzwPgkkDjvujF2TtLVq/BTyDigs7Z+4U8Wd2bHey
O4gzGaiPraQiUNhxjKVAXzsbQcSRHNxCxEm0lIzyecx+qhcqes0uj6svVrWONc0r
h1WnP1IQW1X3cxMPmGn7LktzDDnsH3i8yw0/TjfyLx+aLNOkF3jN6g7Bee+aAYls
xUIolXO39W89pCBDzMDFJvE3f4yTcayM5haTIsY3qtFBCPEsSf2JN0e9HC8idPoU
DIDUEXPagYUVlPRlVQv001+ASsc5rNj4GL0+Dw18co7PKDP7f9McxOKV/7MIA0DN
by4cmqK3mfNjek1C8hMdDiDFk59aMU1ECUJTGF4gnMAzgcz/G84bmPRMD/zeUpnX
HEZRKyf9QpeQc8wMthZrp0NEBQ98rCoDqLkt+Qz/1INpTBmn9qwt5hv6ZBGSsTw/
3MBT7yHbAMoQNy1cnTXLhrogGh3h933v+nxPxpPNmbok9w5u92sWe6lRdUl/VxTb
M/CVHX3eS0MzrQUrg7dyz+jADwiDpqbUhFqk6vV4XH6HVEOEhiWwsjCsEPT+KTyr
TX6w4eIHtDhyyFzHBtAofJpm4tDhr0KJ8OyfuYpRTQwnvX6OkGlWJ+2fL9akPYTX
ap4cz8L9E/W/+hcrGN/CapIc239b/PPWYTTibYFNuPNyl/RuRNcG8xCG0/TPWmXw
jUQoCWt5jkWxwmZsjhD0yagRaEuwxpvQv86LflzJM6flctMu8Tusai82+hSaKLD0
QRlzRhsvnFSDFR4SHc2aVXjFCDSavc3Ex+R9AvqRUHvLJAVNMdm34s4UpNwzqiUM
gmG/VGIPYAwYuc17e4BigO7xG8kyCGAZykTv/ZLQHESGvteH4QSPPGfFA9yiP9My
zmRwcT5CfFmhuJGlCoZ1pGgm+fgR2IY5dPar678gQhdrjX/Z0s5EUVW05CZI6/Oa
uL/kP1VGrQ9WnBpHfR9skN31/IqenlR8xPUmz59XkYT5W6DiSUGGHl7DNPOqQgNj
B9PP/JibqX3Sh65GRFHP3NkynAd2Q8BJHqZtAsDR6y3rdZFqVaiRnliH9iYWozjA
sWgsinz+AV0WOKlWtWoy98KxJP6ItZRpudDZ+Mr1trMTvRKTHfTW6C9CQHo6UXQX
qquGTOKNEZFYPJw8lb17kr6nLdSX1faiG2C8LMjxIz3nf4B08Ep6M/pZn0J07hp6
o2MEUFQuOdYSxjxLJZfsjCs6o9QonioKKNqvYn+Ml+nO+bGn4cYoxnXwndYuIB2d
M8/FS7h8AIhYWqQZNb8XoWBI1yaBLOqGEX7Mo8HWMXm+DPqoqV2pR/rpHsSKjrYV
4EWq80LbFkD25BTkCTFOpHEhJT62pxsWGm+2O0RPI0JCeMAQ2HY6cShFti/+4vBS
H3OyBECmWRcDz98NL8ixTWpWUXbj4hQdbG3z5tGPjKtka2blkcvzeZFVV0FKo+eR
fD0gWUZrRYtIyFAalvZuSDpqsoegpvH3IDFgznjkSX5j7p5DJMxXwxoli7xOi/qR
q0lBohz+2+hJutIFo93aqauRSBJ1rMv1Kd3crfcVhGEUprfQLxiaqc4qb+/w5Lkz
hsTUlvsO4n4B1hf+9xR1e4hZRRV9ZFss2KkW3PpznuJgXPBAj3AcG6CWkLM4qjG9
z7mb8JIOa3QFwXJYxnVm7JSB6qUHhUnlJB4yBnmcYfir+t64B/0TLDF29XfJPRjD
lx5Q3EM2yhfccjEkV8600wTmzxnnHt2wkORiDuUaRhqErYlao7dh9/0a7pYp0prR
BlMrxuOR6SqYNQErTUn89B4/UoFOD4PcrqEzLrEWxc/QJrFtM2qEUazILWDO3Bar
OVbwKhBxcBKbLliV2GdXObjq1BKUYuIPu/Uz/oJfgJgP8OUiEDoiXhPMUDwcbRf5
S0qFR1xRRKvR5CGsbwcp4wM0xe3KFpeLhnnCm80WbUEuv1UPGMUPyku7Gm89hP/X
NROSvjtcZG5YqcrW9hVJWRA0qjeR4+oRDAIySxYy5BWD4sXNyfPVeiSJworTKjmM
fdUhzXwli4fcng0oOw3CwF0VZ5Qo6JpGPrxH7iC1tbBFcDoHUEbKpzwjQHdtQaOz
ntRSqdjEfQlOYG/0FLIBUmgio7ibd8Cx/H9PBA2IRp8zOSxMctpjDdX/el+ddU4X
HW3SiUXQTzONnqjp2P7j3liI3BtxPbteJYCFwBcOr/vpkArZqQXHY084uhpYJLVa
PZJ3l5M4nYHDRTCc9QlY5+8SmxN/vA07q9Ei8WIqzmAA2gpyJjADjR3al5+N6hAB
ZEPmbwTrtwNu/++avOvRvrxhbwidzJFWhF7ZWvMwzKgGwZXDppYpPeCN+5SscOyf
LBAGVl7YCAimme33XtlgAZQDvMtYDsVTrj4OYu81ya8wPFHlE7SYzrgvlM9qOjoj
4AXwof2xI44Q7+Svl2+3oNbSZqzUTGY19TmnWZWsFl1N07Cye0G+pDg1WqsFAli3
aI3tWpvlW4/LVbFaOO1QOa3t0LY996NP7lsfpXQynpIfkSsHnqLrX59CCehGbIJn
J8qSHDPIAqFjyi1TOPrzu85f5c43sgnoM7NwA44jSTXKXO8+lMyKZeLKgZ4+qQb3
Ga3L++n9Uj4W9Ox+tTtwh/xdetEbG/JkuOF/XNODgxmkBWwWtOwNhB4iSxdTMBFb
gFBfb8fnT5UadtSSCSTbQ1G62eX2TcQoc1JzU1wfwkw1OI1LBKTE6bX2DRKOBXNz
h8HTmVv3OPPZ6DcPzeTeCzefqvnPSpxXCicT6n8fWAX7vLz2qWk1CYrHJ3L0gBKN
46L07juDteDDRu5IRPPVzQ57J1JnXU8k9s9ay4ht8bCPP7aIFk+e2hqEOiozpjuj
5bqUlUh0JIFAQelhchs641oGn2FePblI0LyEjFIFY+5WA5UCr/wbVClQo5286FM7
D7BMRJVtmwLq4jH+iAuoNkC2c0r5tLGP/ezqUc4EtgNA7iAMxmlcg4tGpjhrWf93
E6kQtAprnDlhnt4n8cVNbnoMiq7FmK2sqLZXQOt8gBDed3H5Pifz/r4wvXrxrxk6
C3SXQ7m5/F2/9rQOT2oiEYMm5xmflCo+tG+fCqjHDSkJjIXFErWVzDE1oU0i8MNz
/kzvo4Ocb9xJXgVNP0F4gQMJyKYI1LCdP62aziw3Gg0QrvtZ9A6cTjdFtwnijJZ0
VnF8GPtQxtPQdOxGqbZRzlcy04Y7y18a5pwCTWf8+NgO+eOF2pIuJRn9DY9FM5H3
FpATp4cV4BTGQZxNh8Jv961CO4YXYcUnvku+cruESVzVuv4y3mdOhWQ6NCnvo8+H
U+xtsuZ7WHj1Ox/3TDHU/iTUO26FjlU8pzCoSoG6Ep5lMU/EzEF8WO08BHwGMdOi
/X3LtMBRW5qIjZa6/4Sz9CJ0iXjtxIgKpRJaZ5iKpEvEyc1/8Kh/gsKxP7bs6qgL
qJF85mxjY3apA2jxw00Q/PL3+ShSBMJx3ai/io2xJyL6rq3yx9gHwZALnAmgKcyh
As6+9rCE5nRhB0Msf6BqyPDyyFyIPrts1ICe67NyOTqB4NZP4Q0piPpHayhsuDwt
Uz3n84qL+ol4hRkOVhzH4Y+dcVLSckgP9qMnxffft2bJG+Pb6xMyxS82eau27VdZ
z7E5JXIBlsm3RdXpXd79XYWOmNJ6Lapkt5vO1wlx+0ABAI33saka9HjdgmJSVhlA
7ZI33uJGh2ZMe5XZKs8CiClLnLC/o2St4rEv1wzmMleWUiMwFaovlpA87EOcSc0C
8ob0pcoBv+kiehw/RWG8LxQ0RS8IFjHjU9ejo6WzubdKKo1Oqo9KtxVe8H3VaBFu
NgMobLSidwNmk6AFNRzcYXeYJGkolVrxumqieMzCtonq1AVXNwGAAFn1HrRWUIDy
F1P0XRoow90F8TLKJHwpReAGkz4ScFZASvuxg8BzstiWWEupYKj6OP7WLPaSK6Ne
bdeGWh0flyzvTU0rPFHGydejwE/NqoSlxCopCRS54NQmQJ8eDTcpX4u8k7+8p+Cc
XcXlbv84J8q/nI/o14ICcMVIBdEubQOxVMj/vkgqBDBun3zjmwTgBSTFOmYdp+75
wGxXzFa48+H49sB+nbvWa3j4te2w/pwVD8QzweFud7E1YKCGSRnKJZGrrT3923X4
ztUmrCLBcsGiydT4y9P52CatbK1KtEd2+oPy//wEOxwhEozKToX9KH/fk+nmCdbk
tCjusto4ziq09+3BijG/m/O6ASPZF3S+8f3SWyZz5JHKLkEAFdU40xOI98LENUsV
lL424T3A/EHsD3Caae0NVACukiDTfbaSrpWVKRLQdMk7NefC9iemyWvrkRuJkQ/4
A87rgGNUo7ufXe3m4NR6PDgr0d/zTs+kAnmS7KhO/ZOUJg/vzYl5hG7AqAgyX1Pm
4CT/5VhTvqfVee9djj5sIs6tb+uCloc2Zblmlx4nsRKeupHnHf5l/nQFGExAlYvY
C68YD4EWdUa1uCmzqU2eOtVe+itOBfl70Faq9JaU0yINGi76KrRhn08/szsmmvAu
erbUg424X4psjZ0/4+ZSEeEWoLcDRQJ+tvixuNfQC1sAVhWbKzOHr+Xb3JN82kJG
gHrFpMNj01DeTf+n0dVCCjmqu5uYz9tQjbY2EUeIgCHvfnouBX2et6LsVZFRf9wG
W37J4aIv8TgRsz4K//J43RuvOe/DRAPDb4c53+Vxfh/G7EC/GDew3WHQBtRTkBx2
jhth+mViA06VB7Oi+FmVG5me1D2Fc88NtIcOjdr9EreKR52lYeYK+iAmhqZfO1cj
kJdtbSXA8EidszY+pAHcryhtVU85ptk+iXhxIZlbL7AdNsGhcHwdw2fCqSIH1Tcd
7F5c1bZMyAItjDaU5tpLHzIkq6G34xgErzXXX6X+U7XJy+C6iS+qzcDOTnni38rv
brYAybK8aGeeJvlUWl9r1ixFKwEK0HqgG1allwTmjbdWhpND31ZTUad1VZ+9SKxd
tweyGDLITEylN1XRG7vCppWnXZALmSm2r/K6jJ5PVKFswCUUOKCoWNLZ6H9YtqAw
J9SPnxtL9Jtzt43MOYPC5H7FIVUEx3/CJ+46fmEo/ihrkZyin+PPm5PqHEsXdKG+
2shwUAIeTbqHa8bVYEqLTqchkuAcn6M3hGkbCCPiCuXG/bUPac9XKKcsT4IEDW8U
TSswsXrwz+Ijy8v5gkPbJqmyDLPR4KQnkLJBRAVdjYe6vfgffpViBro19dvRHwba
xuW1VgmoSdE7LYumTVRjOGzBDJYLjMar7oEXAy6j6TAM59hcNEEfY8sSES3S20Zn
BCH5rLDbE2s7IAqUdUX7FeKEBbBvWH54WifcKWN1NchysajtSeiv+CoFldZLqAVa
0ubLqktKtJC3XIBRHKG91b+arq+DNErXmLXHv8DVcTkM0xcKOExo8eOMts7IFyyS
BJTiCfGMz0I5cRBaqgLLUxD59pWbTn+N554V+x8YJE03DfCfngmKi4c+sNFVwPQB
GF33jL8DCjOlYQq0LA5uINiCrHZtJoCqOeYnYKdB6lm9IRL0nJHsbC3LbfIG74uP
xYc2SX3f4sildo9XEh5Ha5wHb5hG3z8+JdNXyZe5qZ6rSe6DKHBwdQ/KyJtfJ5mW
eYfbl9rwMgIDMpb7rJlJEtU0/H9e+rirzWiiIYJc7rBKNjafhUTN7ClaiC64uzdv
YEiKxNBlCVlRh420cw8E0hvSjgO+ESkBY9P8kddgpCGVxi0RM322UVf00pC0ZE6O
2h77hsM9DqDTLK9oYlQ1VHHBbhdg3i4fYUSv4IVvN+Q7hwmAXvZXqyF6UedpoOpl
QdAm+/3l89wJ9oxtGAviIGYSQ51xLTonaBN8iid0anrAZ1w9WGQcfK1KJ3A9KMWN
reZ6i8y/p9YQiAC8CpCfMTJ58ho/H309y7H0AMBKdltuNGsNoeEEuYRjPGKC4337
2IYC0kQMNIrfJEy77+J6Oj3yEgg9JLlZ8+y81iM+0ImprCmw5/ojiApn96XdkcGm
OsAD5gRek4USDSBrS1ZEzT0Eubjb2H/wkrMKpP405mCKHObHd71ILS3HDTwgpKXL
kObw9CPST1BXnyb7emVi2NTokiw+wmwbcYad2SjNGGGaSEa4OFPFTZm+Is69UE1+
cEZGVZAKUTuU6TNu+4IPQY52Cv9fe4XKvJhUrm+2VdGrBA0voG9//1COnOAn8e1S
R48bHALhwc08ryYkDBRVO3efbPPu9TtNPEwW4TvXXx9qW25N1n8N2bmpqLwZ1I8J
OTKJe+3KrneMgCgfFpGorjdFhTGwIsId8viU57gcDZEFCp8wh3gjvYLuP71lrQy7
zWvZckJkVhzhZpkJiEV9Nh/K3qWUbGSsdYGdN3aHN4GLCNP4kV1nSjw9EC1h421B
u2bKE7Vs4784TI5WFfCHVeqWxTvneF996DMNkOoMGpNfQgaU4SAm4idyglG+Ft8n
rjGoJVHooIW/zJLlw5YnUI+LYtjZqzFDyi1EvdGCqYV2lqMWaxVhCEsIB8yK8TXN
TJBKGJDYImMpKrH7pdNVI8QL/ekNOcT6pe9qAY+P7VA+H98HMSf1Zgv7z0+ZXRo3
tA3i2bmJxa1f5ImnC6tBMuOzai+xege2ku/3ZG1ORaJK7T9juMC1dlc2s/n2dswp
jhgZVGAwNRFeAogO4fzYDQIYpj3rgvTc5xRfe7bLdHr6OJCpw2IULKjXaqhVdIQg
urXM4dwl3nZouuKPsrlL8clwxYyGFPdeVKKNukRPba+BPnHo0f6IG7MrYdND9MpP
ta+BqfrIJoYy6If32B6J0oRD/C9uJgMrCMhR+q9N7zBQuLkqC+Uz2+GdI7fEgzeu
KrWAbvPvonCgBjpJsFSXwrSYMie40P/gf0bZ1FOERfUCofGEHNTpPlAwm/Ppjxx8
1/4ffNhGnEw1MTRq09RUgVpJc4W/lZZcfgYPOjQwJHuIPfLdsfbaMcDppOpV5GZ/
9ArcTqiX1Sq1l4+g2bMdWlVnGrwJKoA9DUxoYoxqE7gX1AwIJukBI2TSDBXAWsEz
vuehtUVgKwWauqezEdKY7YtEYGDJkEvD7m4ODBBCCzQq+aWCWsOr9vI6f5kEeanT
qWOoUCKK5XvE6/1xRVn5E+HS1ghfz2Scrk3mK8quOnqL/pX4B0e/77Bxmc+ZtIJk
2TwwW5ReprAfX9pu3VXcshAZtqJ9JW9wsuV4ub3ll3DpEM/2CgCPVc3MbKJYAgal
2EzgQCXnQeeLvOJNqDKGqdSg4S7zR3vqJMPBEC5yupy8o2u5n9Jc30mb/3G+0E5z
C55jroeIk4V3kq6wqWU3B6ISAr2Oz64rYnEhvMNUdFA2O+ORSUqpeHbI+oNGWMF4
bickHy+ufFNLbWssFTqSLFFyduMtqvHb1Qru+g9PCMogP9yCevspsXmuj5D8BD/n
FxS0KcLpp0qBQ2vDefzahZFCR384LuzdBwR4tRJtX2BL23fH+lJyzUbM+bhZpPWk
57kgmVePsXMt9aCen2c0Xouy5hcJNwUJekSBOfijPtF9l6fq79vpNB7e231M/6Om
2nQIZgRKfJY4K2Ep1VVyVyfMNU9aakPBDfFdWHEqNJVSMCfxG4lny8pZM/Ne6/mV
N9vfTp6tf4b+XydUwjIunySHHyrMjgw5zvQvQrtZaQzhrIdxqzONQH1K176C/14b
54x047a0huqmy3FILiPrMgn4ixf9L5sFN5wzf2KWRhkBH+PeNEr8b5XSEULGWWE6
I8XpuVTGI21m35gMsya7QEXbG7TzcOc6W/zwEdBLkfGWRvP8vvt+cWFgzP93ODC4
WgWNATcsMVdqTDTmGJq07RYvWwEo/yty/o4vuGE2HGWKYD3h6CmLlfdrafeyYn0g
hF0M9qJQKy80Qn1MdbBia5uWCMECcUtmEKiaSkCfmdfuKOJ7wZ8372uiwNiVkNVm
Y6hfeIokWxx7rFu5q5kXHi/vDOWUUz6WMp6JBWDxd2tXH8C09tzh8cqEz8FXkpDU
eAjjbNnIL1y8QLDuYYs5s3Sn+XPKsQnw8+ACvWgxsL5Cp74fWL2s2kvjoc6KkyJL
YXRbmc4IYS7H7hftldhPfKE/oEOrjHfqt3aUDZ4ekbbA1tiKPh5G4A9WLvhF8hKW
Gp4Ik9XbKxZP6eHsWH/+9bCtZR4gSZN9j78fId7N0xMcXiYFJ//SF41W9B7fNWPX
X8W59Wm30HnIijzQ/6iAv6ah+AX0u43C6mbdHc2HNi8ZGkIZdZcoIlcMKsdCew06
ztv1p9N2DlB2IGRUO7v/Js/TRAzXKp9rkpcWTEO4GR5QA7lhvYgHrbRoBO+1rAFY
mcq7XI2ec16pE3Wg0cpAdXewDW4vO7FuFAZ4tOtZbWPPMF/yp5D63v0KObw63SsA
h1Cu5qK81uAOZ8Jx4IRcUVXPbaVGaUcnSlkw4mHXHoZ+r1C2jmxqp6xtrG42Hce/
T012eonUNC44PHkvED/XqloBxjU6Udfgv/ybGy5XrDIcKDKdHeK1pRenAYsFtvnL
GH2FqYVozbNo5l0uL4bjIPpGdi/OEYSZ6hpS73194ZJzkCVCXJlr64MreLXabT8W
oPRNbRe5fGPKhg8UxW1848eo4m5rY34bZ+uGwI6MMlInqth0wW791E8MzRNfLcqd
RnIQZ+jp+uey64rIY4q21cXWYZcKkqtW/roSpywYuDRoxJg8R3InW71QzbdNC4mt
5NO/6L4QpG0su8VG4OqTfHch6bMSzZTgZkltjnke0IO/dN/n/aCHkQ3zxWVxxD0/
sBKsjm9h1UJXKvZf/PmV/ZgC0N0vJroBsCibq1dn4qxpPNUNdB/WyIe3sZqyFPhJ
TwNgsnD1f2MzrALY/MVugXlWnJgez58a1dNGn6B6qTWW/Eo4C+m4iGbx/ZzaJhHW
oglWM7ycQNBRhyF4im9nHn5Z4fQKIeFp01VsadQWMzJVrvZwSbX+nSwseZ5jnGTZ
M0o/pbvEZPL128kaSIenX4FNqL1dl8i7FuctJ7BZSLHgHkjBR4eXYd2Uu+SNDiCx
rjHv679B/N5+YT28q7lIDL5FL0GlQfRf2ad3OA8jtcWyn3DOXsv7UEhKFJOpsxE3
X7Uyh/qAoUq3Uw9DNBSUrAaamLb3Z19BYySSG/KdMwyQ7CuzTrouymtvI3F2geKX
xF2eqscMl6yUXR882u/3tX2JOGItKAKc4ZF3sC7OhMVyUgCg5XEyBK6CVBACXe/h
9UEREl9JBQKybjx1A4xXampEoo3mzrl5isTCVWrC1HKFQQhfVQE8APmxWpcs5bbV
P0MR6Z3WhqSKNug+s2S9ypJx3xoT7NKO8jv5SKXrMzcY83bH51ImeHAvLiz7pzvs
Opvtmk8t2/16W96pLt+o3lcDyusBATrP7cTSSiRebRfcLQZ6xQwMWoj0mAwR0C2t
BaAw4beKW+RzrafTmqnxSLU3jQH4+3eqh3pAzP9VG6pvnP5rKcvK4c6CpJsLNiyv
92qHY8ZtmTyNCVE8xjZIz5BV7oCWe+/AIrQ2A60ZwCrh1buIWa4Xdq0GjIoUCxw8
xIIuzvEEFPjoFeQRTw1v870+ot4DfscwfRQQlSv6P/+rhXtk05l/QoENH99fkgTz
qKHs5kw++axQNTzwiu0n+a+xIBAqvlouEMzXNdBdqRBr3jZ8UeVIqn+yGpiqBQCI
iMrU50qnBVzA+u69sJi7h+VKBwV9B25EsWRKmQzaNShstkpZMQRACdEMyfB4NhKO
bGjPxjnguvPGbAsQ1i91pe52kPoodYpdKIf8WKHMkqNBeT+3Qvbli2ouZgbL0xh6
GGO42IZDboyzSq+kuYBhkejOVHGzZ25q9m/YwunBqxyElEO3fK55AJ18mvJjj+l4
e3DjfByrIgNDBlmxvv4mcQFEKhds30IU3RyJt1W+HX7eXq8DaCIYtKwmLWvx1HE3
JIF46lKb7nDdYQL7K/Ebf0zMF7s0mXAkAz61o88wempb8wLmJ8Z3TmEuB1CAQz3x
Ybf/8L8ZpYFjFa94XE4dTzeQRrzKe4n88lEiZpr9hpcRdD4T7HLabRScjZsQoNDO
RrGJoXhy7+pNxNufJTAaBl5rJVa+P3uYZERbwikJ7KqWKFnF1/m9AdaiRw4V2VT8
yC4NzB1SeOo2DQ9Ga28IAoqwISQxVS80CnNakcY11MPT4bhEeVyQ1sExLBAQQ1BE
MTtvD+ZugCheS2pUyURHFxELZN4OJMX9Eu53qWtKbWOCfOC5l3M0OmjtvUzAJIeL
yjYgkTyaKmSQc2EvBPqd7z6lJIXrTQ4Rm6hHbc2EFU4JVsu4OxIqNd21Sp3uWlai
w2SlfJ81EMNo4ljGNll6sqBI9MAEXyXENxjYRcEIKKTvDQGdS//gByIDm8COlcKt
Z71JpdbynrdYGawjsfEWZocQ+aRhsr4mS8axoOjvsrJ/sLmT/axQYiyjNq2XHEdc
U3vvbj3bPcfXVyuGnp4XK8JF3BCukRzgvCh4kL3SCVM8yaiVQHNrIOwKrw6nkyCX
jH6tky+RI8PKbrQ16BbhfMVyZzqMdxF2+4Kteu+dmKGXyMHbwcrqRJYVo9axR6pn
RtBhhgzCihDGI6dZI04A9wshrzP4svZU/0AYA3xcVoEBkax6AaKhQGkNIt+M7DuM
Pkd9nU14/rvWGPEtH/0VuYqiTV+zc3qY4Ss0O7iQxwply08EGqJi2OMc5XVOj0To
BcL33X1isJcuf7oskbzy8JgdFQBrrZmbz9D1uqq4mS1Oia1BR2Wmz28BlB/rqtBD
yqBh2RyjKKrWyqpol+Rjbe1nmYvsyDIw8n93b5cfcdgSmWdOGhK83rk0c/pwjvRW
QZVLrjOsgXoD3H/qHeQG0FLebTwhYnimwUPHazY7rzhv/28vdaEZhzW+hE/E59Jh
9ilM+7jlilYJi0EU1LYOAmiUX3X6NpSzQEf1M7xZIi4BVM2GX8dg9nyONZreCYh9
v4tBOtEjenqxA9b4GpkznpwAFSxPTScUlpM5geKJJYmdGmEyhejgjCAR/2GG/EI3
tns2u6Dp60UsT7bWbPP+kXYeNEeQFAbRazHphrxKichSU7a6gvUoXY/cm7QMJ92N
NGnFyVb0ch7ttMcSuBXWcn7nAmPHlcMbhsMsrEgvlC03tKxQxWhs+9ieN55/MEhd
aWXvAcxhEOevH8Ii1qK9zYapFdm28uIwt5LZ15EEx2rwzlwShC2ne7cB8nf7oBHB
BqR2gWkBAjOVhs2NvBCpqYI1IzEhogUO4wFkBNkRth6xyEQO9FdNR1NjbiAPQ0Nz
MDo0CotRa+v8Drz9Ldjt0/vNa+GsaSbzr289+oMiFHMwE78KaqaMObf0dUFdJ89t
A8QSPDtOqJNlbVHAG6HoM21nnXf1pCWaEG3/ZEyS7+FdUZOglMAdySZJLWhObvCG
+dL7gtLWj1XLgm6GvZWQT4D653VG1vCTMtMu0aTzfKPm4csc+uiLLVEP3mC0qfyI
kcJXxAVVHI2an6yhxzclkCeOfR92nlYJSEAjZAHvPgbcCLKuJz8GICwAZ4icdV3B
JbUa/sraAQrvwu10bwsWEUVp5hWk10u++qHDlcad/zKhOI9XlAfpd7AvZUYmYYtg
jJ0TMsJcKja4Utr+/zUNLl44UknVLh9Y+x4gaOmRsfjSgldjanxAlPkxfbgIIxVG
nvWLGSeWAPdmbK4s92dh88bihqKcbfk4w0os3LnFd6Twcv6JTHPq1qxq8SwxduIK
x8SzYSVS2jG4F16d//X8h0qZpYxFHczy+lyR7JzmZwQIS+cYRu/jWrRaoU+RTTbU
govmT5Mt+ZEtd5WOz1q8ZRaaLNXxBoZ03ttHjbbndRsh1BM519J512oEU9W43bZz
3rOpEiuMKDhnTwYve3/9Sk1/SjanGJpdfmzxjmwW8ZuDVHIHlHM4r3BTn/kaECJN
qzvzDoHuB9+T51F+djm6hHSC8i7rCFY/SlC2w+DcidzVIjm/Ddcx63PwnF0PW8y0
/wb1nEjX1gZo59W476Ykqr803tJTMDMhmmK9N8XVZENTBjXUSNE1rDrRFloF5kaU
d+XMTmK6cuEmqzzkxWukHUWYTGOt93uta7X8Uz/vZftR4CuqBokiqN9SlqYtBZyZ
ubigKQjLtdc9XL4Pdcfp7sSMnIGFfbtQmkkcM1fAtKaRmnyB5ROmNyABZhXHRYzf
pqgGL3P8ng6IL/MIVb5LAjd1U38yN0MqvDc5UxjVhI80E4iKVHRvKLn+OO/X22bD
t0Uif8Tmp0GWRgPogLuCXlHv6FP3nx+h0DIzr/FX+m0dNIxhz1m1R6sF61x3urIz
M1bquOVKqTK/doJu/2x/SKIfBOXeDp9AisBCjvBpRzKb1ApyRAJifDMqQyrZkKAg
lMdmhhqgxLbz8udrgKtSoEr/XVw7YPsLmLd8iZYvcyK0TKfYSJFgmPrOKcj4wBkD
+J7VlzmAKaUUC3TaszF2HkGxNF4FtC7O0pr04j8ChtCV4WrdgTb931N79fsU8UGB
8aONQVHYwsO4WoPRdEeccmosWkXEbzJMChOKDi8icavj56mBkcc2ZHAoEnxyeRIG
8sDELeWK43QuKX7kZnqdsa+fj2xtSRDMM/Vg3Z96lwLli+PrBPVwIex1OUuO8xYN
4uziwGepxmEMJp9M/OEbgPYvdqp4PwfweO8CLo4aQ60p8LdA2fNhUKwccOLf9fr7
vQp4YX/JYuXG0UYOLmRE+VNxlJ2KvXEwcDzP7o59CqbZ5iRQ0A9Nh/XM/NUKd8xd
S4VjpSsN3PtnayWr1gx2OOHQfBKh/VnHPe43oZ+bEgupTofwWEdBE++AFY8Gx9xF
gq8ezWmkYetMOsQUbUVUBfhQfP5zc+XAPQV1/rqDgaKiWNYR7bdyc7qnzNQynwq/
OkkX+p8LtxN7h2R+hNMcF7NDK3pLJpzyJKnTGfEsb/mHhJmVY2VlGGXv8muv323c
Z+CRgYsUOuKp/HUSMaCALXf5E//6xhfVDfeCMD6yitfTgKDZYO46nrCksmeuup7T
d9GSy9j2fNOJNIa8JW2I/FrM9AU4lSFQ3MmHsW7N7jVAMj0ieC/yM/q55wfUcYjt
J+4FQG5MnRrh3YVNtSNzPeF2s18dPxzsFhskeq+xCDsmEhZXOrC6mLUjr6ej61Zu
/vir3Fe/rrL1ONPDqVo3C22so5+pKAYV5CxpMOeBiz7wkdAb/ElCAoNh7SDMGGi1
e/lwgVe4FVhUvhpd6nKgYCVfPHyJ6sqgoRvlH1mvb77OgN8CvCrNN9XTTaIMAFWz
67InPV3xjxwyX2YT91qHGPVfq6NKRp2dON5LYNjdTsy1f1Tp5A/l5mMLLO6vv4Bu
4gX3zMWVcWTm4pPYJXdjU7bV35w8xImEo09P3/mm/uEEyhSfGRGTdflQy282OVq1
kwUc7ToLJBzHmKGHtafl9CEsz0L4Qs8upnHVurK55xhYBswAlWH8Minte36YDhZM
mK3XvfO8unkYFL4FnFTL823tobxXuq3A4M0yMtF5BqHbTed7GaxfBezPryN4Le3Z
c0E8g6DgW/H9MsdhRODg5/8LBpoePKgZFNm2I6QjmpHIBmXuY08lEVzdmf+nKgnb
4RwDwAZ3dtwEm50fF3wSXZuB/SFPfKaN3HI1mhNHcLX38et7mTlul0M1avpSWnKX
hpIz8FtKavbj79UZJ5eBbVMvtuT/ehiHIdUGVmBYBAubvozfyFrhRmEFHeCAte7Q
RparQ73X2V3CUJuqMsgktBbOsBmh2WUf5TatRn8Z8ttfi5Ski+5kajvfRbummTna
PQfwgFpRIkGmK2kFWBx05VIw8RVIlrKAcTsaElzbYkF12cZGO1iiDO1KOZvNO7I1
+NQ5nCURVo++OIErb0hubMM3tjNSqvk7VZJnkAxlH4Nai0eqNzR8Z7g8L3M+qaiH
z0y9rdL6XKfj3WMViCz30sTXkx/7MMt+VXaDvfiy3VF1Rdd4NpRCQEJLfGIAntMz
lGUYRYOPvuZ/3XRgyPaA5bkWE9/27tWlV5Tuirk8jFZqyYX/Tp7e5jMjeNxtRz1g
DwCW0RoJ0MnDJ8Pvtv66EB+gOTZMiFTen3/paI9e1Ge5JS4fMW0bfYlyZ5R9gbyo
yMyF1tAVwfLLnNomSCZd44CVvFm1FNs60Sp0TtEkSS3GItC2R5QCzRaTYjcZPGIz
NVc8zfYKeKPw1sasBojdTkRpzRGM6TlR9B/c69Z7/CdcmtGmUrhrP8V4uFvUhE2w
zwnCaWRNkMYINw0fk6OSTnVGUGOJjLgeAAaJL7H1FpU02rz5tJeAuxNEbdIVGJwU
NxO5R3kftiDygZuUo3kb7W55xSvOTUX4AvIh5cZrLSdhJWZZNzg7Ed5brGxmzwkr
D6O4IEpSmwcChglQlvIzXbxSF6I0jpWLJnAoXYAg6gvpXHB1eDeu06NbHlqRzYj8
qPNBULX8bmYD1VL39X5NYjPOfJaYRI9WxmVgjH14jZeu7TwXZRRlk3sShDr22u5G
WAhUzD6qS2dFQNlzVdklZTr1rmImxW5L2pXPKLFT50zY7R0m2tJqk0kVe768V2Fi
1FB9zylXY5u1tk1vWe6e8M0CwTUrtPRMIRBr/ijyPtouQ4Lvy9O6OyxglJSinX0K
8gfiCuHRsTU95Qvpic1NhdoJQ/kXpKdUuHTUwZmNyiJ9jt4sgsNfOqY423ecB7+p
3fe45FK9KpWsf63pxiWnVUlF/sR1TPB1AA4q9ngT87kbkrECi/+s6mo2TY75pU/h
2043ac09LhxwfHq7vc4RuWor0TrJeWtBYOsu9DLZA1rcSkmovR8MwCg0Af3kphJF
lc/d5PPJzIeIPAKXoKKqUSlZUkPNhj1gGO8XdSEr1BmiI/n+RcvHFBy2GeIOHtZO
ODDydsOv6Qvnu9Q0k45cpGiq3E3m9w/vFA5zELWrxbfMJVN/QjrlyK2WZFb1mNE9
DFHHDJPni3HzmBmbPS8vb1Uld6MhSFcCrf/gFpLEHaKoSt+SH9FDJ6gQw/zCsYbw
hPdymEbPF+XH/X9uPn8qpFpCMMy3pAKbMIEM5hlFskHV8uN4+gIvIt++XDi5urtB
upx+wpboI+/LDEIN/val6ut6SMwYo6xw3qISAvccGJ23wVGIqftESLS6Q4IFaHRr
ZHg7bcDkCh3L61yLCseFh1vlJUQAmWToVvipGiHoBcj5FYWBqjynvdhdvTZK2cnX
LqGtTRYF/zELt8zDHwYyA1BhtjOHEA6tspA8s9yxjJqWDcw76/RI0b4sA5lZoi4b
Tajvx1eoATHH22mXpa2n5TXB72SXcKgmjg4FTXoClNHAszopIQnFJUzw2XLlVcfy
RZPTwzwvU+e7rfjiMx4h1PdMKDJkcB+xzpmcDd+KUA7KqFg2pu4feXshqp0GPqnU
XXxCLqqclqobcpwQ9F8tACRgN1Tk0NomfGZ4gCD3Nt+ofDte/Uf2ggPeyYukqiHo
Fq3lNTcEP66t2IA69QxoimiCgSLzOrAxqRNHkkUxYRy03TbvH3pbxxlC2AKOT0I0
X1635clCopJOiTGtQdWn216WtVSNJtNqxHPmW0mOkNaqO9l2/asR7LpNr+kyy08h
Jt6ca1Gcc4K408jxiahfXmGPGth36aqMZtZHaAU2Epxs/7JSC3Nim7nZQXoUGQsJ
v4jO4zgEe73lBm7xluhOhg99XtGHI6+03C71MXEqAdcWtE9XN+3EI3dP6ISPZT8o
VqA7CCEDfH0PnMcKZOSp9YLLSP9N982we0p70WVb4WAUDiEUGhlgYkKOcKNqDnW7
BUhL1HWzzWBgfNZdoT22yPba6Bfoh8JzZiF3JVsMINYBm6bIjwianZs8eO/HukpP
QAaVqPFNuD7PXYi/FH1UggEymEEBiVCs6PycI2on18OHjMXPI8XY2LWPVJ8UatXN
2RYHyFqvoLJt1Qx4UU1eo5sZPdb7dExfNTN8wc7tLggZqbcfTb9lU8Wjl7X3lve7
eohmVYWFuX500dEey+xu4JMKdCqEoY6ZL84MnAUwrN+PnREmUbcbzHJX7Ny/F429
DH727nmQg1xRP3gkhJ8+vodL6RYvw3txhQrPzi0QpWJ3u3gdrkLR5TSCn9Uq6qPB
WC/zzWVB2AoO7X4ArjPG+wDewJ1DAfLUqase7ZyujiaeG3cwionUk+XDXRLi5czt
czyePHHl0b+sU0WPf55d4XHlMRsx7F6yQOWYdFk7vPiZL04dH3S1kD2menFdNlB9
dtvofU0dwpOBHDM5YniKGqxMCBGIUaRdOMnwMZq26AOjGWFcUhLRZTEldQCZ0fy1
e9XbpSp+l3YQ9uJkfVrn1k8IXaQH2uWmSgEX6KeqPEL4CLFWgRzg6ruax1JIyMlg
WqkGgBecEERe/IJgcB+7SqraghhT56fxSucGyLovMMCe3JMb0vBSPtu5cKQqw2OB
6FMBunHazol3tUl/rbg8XGVmBxAfVgZgRb+UcUsnCjyg+cvD4wRAoD8/7KNZRKri
Y+nJD7cf1iSMwtH2nt5j9Ai/dznUL32Z6fl2IB/R5LlXPqb+261409slzrToJp1+
wyHzqIAqtV8jT27YlCREsOM1CQzJlZ0j8XrMyYyyU3h0Ig+p5b+C8G+8E6Do+Aag
fW6OWk2faQfpED+XDiN+bBHLTue6nIsO/0xRtdO/Zs8L7BNAZ5pNIS7v+8J9IVT3
DoCKth1U4CdjE2WzTuNuxk4Fy7mQ1k+wUGC+y4SHkGzl7dIdXclbbd9F34IFIvwu
7x3/4OkeQU75qroFNinRhzeycBkOdMBhcr3DEGj6e60cVA/xeUc8arVK45MH3A8p
UjTlNIuVcq8qCYhtEiGVNLvZvy/9zmFb/V3j/L3HraI4Dy+7YDS5za0cU64Dxp/j
YsTz8ZmHC2bs8rtZDFvVe9dhrNUGXIzMJtkijeA6YFaeZdJGH/YzdBlrz+IHaMDX
y6wNLL1wDeYAwuO7okiMCfDsqpkWrYtqepPX5jY74QV9NZNpUgjfk8JLVRaCMaxc
9ZGIdzVgwWv4zx64+8wRnTFoHLkNDGEn12Zssmizo8HxQuGWZmMKVG44Xy9Pnf5J
i69iUlzmwXiBK+8KUlodsW763C3c8KInxbZA4Fydis8i9tFU4ljD20460+bBcWCe
+NIuLmwdak6uX3FpTpx5aN4G4GZZf2pPqPCvkT15JVtnlctAD9XIaxydmT9RksL9
itj2kAoTxMbSL4DKWuKqsXdxNpvWCObNhkz2VFJIr+p4yrURn82ltFwQD4irbG/E
mvawundu/ArwAkYm7fdQvlhSABi1wiSbNvaXcBKQdD2UwDtU0kVBPBZDWCCJuoaQ
mwfVOS5QtqyLzuSMBKvrSCyXYkWyqVVrCb1TZM8l1kDABDAqo4A5BRrd3L0tPKVa
lMaFnrAgSvFwHLv2dwDzh/MENCNWRopQWmENflK45EtmIDjGoQ0CKpGJubb16nmN
tnOo74q8l63I4GT7KHOnt9HEiZEnJVYIaocJDiuBAaHO8I14x7pBQ8YBp9BxA0LE
4sd3fS1tWprkOJo/sb0A13jux4E/5YuEpiqcZzkm8l/1Gs/ye3if2DAfD3X1BlHt
09GcHSvZd2XohEh2SP2V+gDRqU7+z5fIxzb30FKLfJd9LGm+X4lW5jvlW6VuDnMy
qtqn+EhKAtc1LrZiik8bb8sSfOnsbWSP2yx5cRw8vEE0GjCjYZxt3OkBbqI6ITrZ
tuVde9jc586MNYp4ewdlP2cMgjQe3FM1RHsKfAV9hu4yAaJdWx/Vby+8G9TUsNHY
nyMIYgHwp4PFTRQns3WaZRq7hhKesulG1+TEAu1Geh7NbL2TXMEUDMrPLHd4nSkE
JbSrSw4vO80GM7vM/g6epIJICWU7RxAcVvgIOb4fl0szNk8KApODCiWUh+gM/cMl
I5QJEzvFYDmBjpjyzaXTardktZLZFMpPil3iysyz7eJebUjVmMj4MHVjfwPd6PO2
IhVCdgidAOFs34W1q5JdMsrqdH0w3VVXKBZstrPP55+sqC3LuvI0vvWIDgu1eUGJ
DY1YKO4uRxMlcQoOxR69+qd9BtN3BNeMQVnCaOOSXYQCHJAEQteBX9TVPoAdWzHa
TmsxvktsPdg0zgaY3cdCLVgLHZ1jtCaj0wbQhx9P9cc5sTMeUUGOWpoDN3AMtESS
f4BWdIfGOE1ytNwnruT0YD7VxLrpWh/JKR7Ggsob14MGw26aOzRQvQ/2Z4Z6+MSM
81dgrgjW0/FJv/cZaBADgdMLJUvi4hmvOfpAXCuaaikMuBuCJW2ZYqeLUP2ewLMj
Stp2nbd8iHXsgPRt/d5lcVu4siNw82yz/i5RLzOQiPSaH/m2ZsBJ0q3g57qfS4Ha
3x2R7Dx118LxPvQWwOa3/5ot1y7hd30hVw9LnfMW7nm1Bg7e5WISt6VuxTZ1dhaI
At5GotO7EIaG39oBNlKy4EmVXp8uZkFDouQ6CzdBWkqacrUe7NFZIG9t+8fzzZOu
JLO63GIYJBJtAtcq4ixC2fPTuFCYsL5lesc9XJIzMXQDGJ8xq3YBmSubIIwqLSEH
YEs356O+u1t9pEuxpqiZI9ogRvE6cNz0/WDwLs1cZwjyDkfmoO5i0MlTuXcnLi7g
GBieJDvbomJ71AaAyCggDmhpW2HQxPf88wdce5HNaItBeOVdc2sF5biArMN2DXhp
IDPcjHNd0maENIBCSqu1TGHpvsQmaKql0/ujn8S36Ipldk/4WnzzHgXkgyN4MToy
1holMQPRHCZzX5+47ZPWl4zRNbjHZU6Pc7cqhSXmuRB72H7NuSPSju7Spf7ujl66
EjeW1r5BpdyMyNyKGtZOcU1WWoaf/vSChlVs+JwDjKdVb8XrvEriG42uzjRPWjgF
MgrI/8pdJyQ7UKD+dZgbOhlW/tsRxSMBdEA1T1yR4bO5OphG0Ggr18KmdixMJNDG
i0EuoTp4CBTOaAv1fnK2F3L1WTmq5kTpJ5N3k8GoDz+L7Qbj+HcFyNEGWUMI1sVP
3bSpPkNzl+iu1A0Wf1wiHY/krpcyHzE7cYGap5J9h6thHrcwJ98+31sZ4C3xaEM7
yDMLBjYJLIJnuwMwW/UveWJ4gi8R3L4bFadV2lpUVxxr7MdsJ0pRBk0p02gzc1iz
MuXHEF8L0tEzaKE3VvGvIj6DGPaLdDJknd7WVErMNJu00EMjfjBPNGWWOXr9HkSD
fF6Di6uemfvXYmmlwtmsaViTGawwc3UrnWn+/6Ep2KTKzXBR/nG9kHNF1JEfRMRt
Duyif1VeonWlawJfpg2dzIpVAMz20cdHeXnamAiiErfVtt+Ob1Vmob/+whihwU7n
kPC+62IKi5DVLVDJ3yxoTAUIiVtoPJR+dbvf875L/xiSiJsIwHBwdsgqgXiPsv5K
WQSpsHTB4JLfQgW7cur7yBW4msz8fcwqq0ITh9j+gdGKI6s7/1S4yuJ2mIk27gPi
zoH5UHN6ek/5gi49LCQjPpkwawrT2vHd+Nk1rRSpsUKybXdAfgSFKVipicHpKxWO
Z4F8WoLjc755a9gvHb7287aHrOL5Gy9SXm8+IPFpcFiLoX+TXb/hZT8nA0lnDB9a
EiSFYsvQusX10MiDPFOKc2hftU1Fcqb+zF759NY6eq++6R1amhBxocp9kcUNZ9NE
KdDYUPlWPPymwS7LN+diu80/ugemFea2u0VVof7Is2EXZgXO9puoppkUtT4JLIy6
EhglFGAMjRhh1wWG+OK4gypPvUNObQj6YGac2HiSttgcWxpJHSvyaxeU7Qa/ybob
ZYZr/1Dw8XWV3RR10vJey/p7fY3WwqtBfxOEGJMnmo2rRAfj0CUp5NZmvFW2vTvF
SCEeCvXKDt7ilXE7zHu4VG7rrGdHvxK9uqmjwi+VjcIjsGz0YFIOhAxln+seonWQ
3bytS4bhVDnPMgWWderwxpLfRFhkMwOmHil3RcRR0lnlbf0qbtF0EJHL0WkXVvu4
ui8P3fAuSu1oml9uhBMYRPiTVJz7C0LBOo56LyrnhVuTKGzlhe7GFEH7TF6PdaYR
0XXmsw1Wcn81v46qitfT/GMmmMUQ3y77PZRZdWsqjVIVeBWUOnsWA+eX9GSTYF/h
tveUBEQ8COYeWzmy1YEXEa9T7bZAJH6era/lXeUNW2Z13yXrXIuCh4+RXhLodwgG
sdIcnZvYUP0nYM5X/9K998CgKYGDPFh4zDpuFJGO5yyA6pCO9QelpXS7Ot4zFXZw
Rnr/+BNKFqqTVRQvvbcj8mNronYqA9tzYgjZakE6/eVxxn3UCsAZGj9I+CF7b0tQ
dwTH8WY/vDykXlC/VJHDJ8v1A2N8yBGOKATxsJjXaY0vRaqIp5UtCJz/UN2DuAJr
liyHGUr0Ow5bC++PUZigoQTxuPEBzaj6ddNL9OQRC5Xfq04W4nFpEpfxqgaCLNWQ
72bTqjvKMgE0LIRZ0H7qj7+2Cn6meeRee2Bm0nEKXTOUEtyLPz84QR8rfepbbnLv
QNdWun8RefUkV8GoHEtEqcR8lj1UY1i9dXD3q5HDXQ4jbfhVLO17QqK+XoNtatdp
gONWr1NCt4G4hammONYgKa+xA+LTAxnPd0ucn5czhwPItQQmCZ/r6loy4NrT4adU
5smUm3GHX3jCWmjPmPNOiAMe3kJ4kwt/41MrIT/zfy9Irc7jrQLcbTAv5MqQETvX
OeD1yLN5HZ9fFkZzz9hKaWSBQvSFbNBPJv7wcHsyLo2jq9XNtDDB9ta0ofoh2hKG
BPv0w3aa5aYsHH5AvNZTSotlWFzZsLI3lnxhJ14gDoWZdYUfYZuJx1evOFaNH6fg
u+tkI3XQB7bNq1GW3SUfEilBHryQHtd7i4sEe8IuHuW+NMIZRxzLY+OLTxXwrgKf
CicrIrVCom6ll2TFzgL/Q5uLvEy1n0/cC4Q//z++nrD1nVHBcv0jbDTE4Sj8YTok
qqWVTu/3G+ZmFGJSijWS6CXmmVqEv8pMJxzRVz9nCMnVspkA1EIx5LRghFXKBVO4
VWtJL0SEnKT77VzUWTTLhdNXtJiCaLxiFmWVh7iiEU7l32+Cvq7UozRcgEezXLac
faB0IVO6pvWrvITw1G9TiQeoCOvY+/bne8ga522htUbs9Lc9w7NRA2OoA8Xf6nZP
c79tk0ZPWCp4meUxQCvNR9u0vcE4rY9q9p/MZEjv8WlDaNKPpkxw8AT1EeehYvqU
nc5wfK5xGFJ1Nh/0CcCJdWF6KLfRVyf7TzGaTpLjlxCInPmEDNj8/HGB6xfiji+5
7Txbdn97F+M9rokLnTA6ecifqohcMmKC6jmowSCCa9C/4zQzZOhPc39Y8U2SGReN
bkr4TthzX+yImOEuuDc8/MqsAaQpvqae7yYiFJhW6M77K2SNvCIU4LOp9YAPdVLa
1621uL4ky4hHzX8/A9RdpNVGYjuORQU4jf+wJzPzWRmY/y9S6fZLUKP5i7Eo3Ki7
d8hiHsHznMZKASlSym18qieUwY9fgeBPQQN/zqoBwdesYN7SDsay+9Y4bUWp1GVQ
qQGsx6YLLygbR3s6OfJrBWhKJdCs0D2anusJrVyXFN30rxmzIcWinnth+8moyK+Y
kaPO+i9D/9K8Is7e1hCHiu+RCqcnIBqDyNVEl5jHhOPqKDIF703tirGF+6NCbrPr
bxxMtyL/XjIvYG4nnlJyKGKo/L5k24Gu2oLIZggHZqZQfmI8GyPh+EEu7G/AzTcN
nm1SIxbzXW6mlpUegH2ZYWZbpP43eR3Z4rp5LVXp6wPeXUBismRACPxN4qgHUDjn
724HXBSY0EkH+P3xn1yNRzoDBN/rkYq107k20+k8e+6OTnzZ62uLm8sQbVObdylp
ZFkr7vn1GHp3CNtcFTKqZ24arBGnBC1Sc2EwTuwY7jsTswMkDecvD5OztgjABWkI
r2Vup3Zxnd90aWBAEPMO1L2T+QMOp2sK4+DF9O8eCz9srXYnB4eWc5GBbpex0iOe
QpxTGcdxPyLSH8F3oKZDRQqpC6K2yH+w2BAq7RZxUyiSqZ/QCienYQdxJl6a+7sN
G8w0yfaSeynoBZrs0tWpScbVlyS/Ug8wxwpvhSox7AChpixAEuN7XOauREkEfLch
QZZX9PuRQH/yMkUVbwYub8U5yEvneBv2xIYqixnotj9X0AXsnvKfZX4SOccMo6Bi
fO8Co9TTgIlYFGy2fHPcPqOeN8FFtZEWkyuUfCDOb1C7wxp0RBVIzJ9swHE2R08R
7g0kB/b8ESr2m1T5oqe8BoFEPiAbYNPeRkfJsAUlgpY1172hPV3BC5jkJaCBqK9W
tGevxXtf7xpVFfzq3AnFh1wELz1BD6lP/LeRPIdzEmBuOO7RME8ipdefRQ4PMSqX
JfUOm40ajOSu2urCtGMiK1sCBmuvK557hj1evhBlMHLRpvnM7L8kVfy0Eont7Ex5
Oa/jbOyFE6uMTXi8yaaoHESQEFKRUejWQornQ2te387p1aEaZp3/5c4QYNd+ifMc
5/5keT0e13PrVcgtzndOUg0nA/hA3Q6YOIJ/9kvsW9vup9gq7zcCE80hdWtocQJq
jCOisU8pswzeBCw3Kn2Jw//Pvf+KyD1KUZYsgQPO3I8uETQ3dihNSBzvnwyXudht
4WhpNEK4FuppBWVj36Hs/aTZna8GTYkn796YMU7+GUoD1CSRXRimIHVGUp+1lbMq
NPmGdBnMhORO97RJCg45vnmj7+xcid49pIO4SLGxMteCDIXI2cxGEaxUhzY0ZZQY
FN+dAnA37YsD96jNZ5BmS44dTewAcMY1bETyUpsv5YNX6yTWxnQM9kiS3yxv/gnZ
kNIfmn6XqLxf6giiLgdqEV/CsIfiLlwdyt+LwNE8NcW2zb45Pfx/HRpwUY1cZWbA
EIp95Ozg5M6VEkmxPIZR6XzwIi0XWEvCUlj2/hy3JmLuGrshY5Ira+o8vTY2SS+N
jaaUiTcqrydzYx/rtwF+K1F1bCKfpXtPQOdJZPNJuGldW0aNB2rUsnuWR1IVylcn
ERvqYxP6ck4RijjVUyyFBHmxG0QPbvmBvi0C663t0Ywt7qVvVBwpJUcvFqzSfyAa
TYhQHvYB08MuCDsDlHfbrgSmrkX/eq1pNObnQiXoh9I1AU58zUZloS5rwYU0R4q6
jyBSBt3ftm44WLXaJnsqk5jRl6gceQZLhhQ+G5MI6Vnk3JTdvI+XYMEM2i3rGpuT
l2IyGN5P/MgPSwYfnTv7uRmy/tLeBTQb53hTLtcvhQaI3BhJlaIejcSE6rxHHklR
24b/rJ2TcUw5q6VAqOOCRo9cbXr54RvLuzlPUP4o9t40oduplYwhMI/+kMnJ5d+0
GlBuV11GERPDdKK5YG+ia2OkukjfHazJSjXzzngc+xtjNLdJUaEAQOq4Ui5Gr1mY
B8D1iaBhVJ3eLAMmgHENxa4JB7//gHqHhw88AtQXGSbheNRZIdVP+g5I3gBtGMHw
kSc5W/PitJDDfBwHIr4HayRHNWTHnjUVW3qDcO8hdGxv1xMvsTMcVntCFQxVvkWo
CmKXDuHtKcO/OfGkBkBMdZD92saL6qIanPzKIMUCkt47nQ323hMRJ9U3EbpCoM9n
VrutXNreORFHXJ6bLpGMo+M+HyXJTQPcrCbTgHEExpArHN4SGbPeF1CJA5XEntk9
VPx/8EZijFObfeQYUcujjijvVPm/c/YqEgUmNluD4WhO4s/F/gnAtDvYkN4PteHn
wO/E9tyykBW4fvkSp3texmpEfKtEdIBFBYmPmNvsbGlUlbEd/9iPaVif88OyYd02
W7AMZ/OpxufnDbfpBD39kJ2vjY/U5fCzJTUiOjjBI8shTWYUG8c/ytAepL3KLD8L
6LYgp4qn2PJ6uiIE7AnUeq9B6rvU1apJuYNS0glVbn014akF4+FGGbdk34OMiGIx
eZLhc6IPwUFB3cFJBiE+I/Ni6ajv1LXUhtiw8C6FXB8ARju5asNXxytNhAycP3Ob
JCc2WY7xVUt4dgSb/ZWv+HIedpNu37rb97MpUXQpCBMG9uQTgRJTmNNKBuWhyM4B
HkDN/hivSVzzn/nWPdWo/tKres11bIyqLA0/RQGmX+Mh/FDyJnLws/1soYeQVdiZ
ytox/GHQAxK7oCbMWtK5u/FU7k/qNGUP/52oVflLkFcGvj0hvqP3azqhSstDeTgu
oDk8hGFU1QrDQ90mduJWhzBnJxOXjCV4cKKp1Yhh1nBIeD3V/onRhiFqIYKdS6Kc
8T0C7F47oPO9JWVJRwl0B1areoKE6gz+sv+fzELbsQQJ8iBh6nlaJ/PRjo8mj8Ws
dMG27qWvGSMf0vvMf3CBxQUMdBG5NhBhOrqujRJhW9K7XgPHwlHY7MWUek2vzZqz
Evi6s0F8RfWM5RW6txly5JuuyrVMvdvsD1oUYGLgt4K9AkXj1YQSSgyCa/g76uxq
JsrX4dN2rByv4e9v97X6K6hz1AIQREvIrzBo6DkeEm/W63JO0vG7A02Ra8xbwRUn
HhtPVxmflgge7WTYm5nkap+xZK+WmkH69kepKD/Z5KyfrZ3qGVcmYgcKVQnqC+kY
rtQoacUPpFw5EkedaIJs38whk5L//D7JOumy2DBkmtAeC+Gj9+uQfuXslyRVGYo3
y2XJR75IAb50z38fHVX1a/GsiuKrGeHKUjB3Nf62pbZaEbbjnWh8qBg1PiNtDInp
5NnwavEy3PmzMm0MpEotpV7PWrWAToXW8U/lH1X7so8+dFjWenxfkCd2xOyfe/SU
Nm723YSN2aLzuxUst2yjT2yNoQU+R1g2rB7NT2Q/WyHAS92z3ql2wl9TUqniv7IJ
+DSln/BxjCaXRX4Oh76GFgoBH0qJu+FAPcf/J6DoA3CYaIJecfEpiF3DygWyPrtA
pooS21yIcuVMtQjPuC9xktChLVtLanL3ndpzW+svRDQ1DI4OcQ+3swG0iAdPCQmY
KCmA3KePqzM0qPB9OT28IOeHECeLcjYhEvbQunUXXc02gRiCoV5CGHOrcdrMpbVc
dP6JzzB77YwDQzIB5wrHRIGerExcFOS/PKc1JTleGGAP8/HmOIbSrhF8tscO6BQY
ZAKWFVZB5I5XjNRlznEZKaOaY59/W8duMAsBzZz8gWq5jYV2/INBK2yZNQ2v0vuw
AsW0ztD2hFx2sZw7nFD6jLgNA1lhe9ruScqeeu5Wd1yCTE5GQiEtVkIWXShyseI/
TPtd0dkAd57GAJGDPS+NnmkLmvjaqBlndwDQIyigQjDowFPFrCpF5x/9W2ChvGw3
fHdkiw5BqFjH/pyf8P61qkeoT3snutxppO4p8OlkmovJS1LQT0vDu8dU8EAErYOG
DeSg9aUlR1mtUCH2tyyDkEex1D3XUSI1JvSrwMur4ogRjG5bFvoKeLgN9/IiGMIE
nQTk8XEE3lj0Nw80ernwHA6HhG7BRHwGXttXxW9OXVW+BMSEl0U8hEXndTEvhVPK
LFFWVQzQlDptn93fxer4fE3ZT9H02nHBRI87hMpD+pnjaSHAqOZYX33CaEh5qOLn
WgrWiIR+8taE3KH1prvRhGMheYzQeOA55jI7aPH2UPf97SqQ7TeT3AeJc6UYtBpE
VhEGAKijXfyxEZAHjwWs+KyvmUtbRGDayCl4DuKsfpfDlxVvmiiWy1lCMa30ZAKc
HObtvj5gmPfwK4liXNqD+YrkXUKf9BdM6xrBLHTapRwv7oO0e8el5qQ0k2Ujj5Nv
gD3WcTcJGY2GGoyF6LXIP8QwqMbkg0qsbSM8ltCwxdNjnf/DjAVSNiU8neduMvnU
cB9w5rkkOKn7JYg/bWF3Aebyw3UX6VKOixOmHmySww8oQRJhnHimL+txNaCqBaEi
le8TJxNmWP+y7TVAtmSOB1SgXZh2AcD1DpBhEftwATgiuFOEHoZkvmRf0RhGTADx
An1Ae+2m8pCtetwDnjI2AnsnVlbdQR3co/ZOTuTiSy9J6SPObAep4Ie6MXpV/ohr
NnBWybPV6+BoLKGXLktqudBf3WY8FUjtffzRwRFiW7lCLBcmQe8ThF31Dy2QUUL5
gBr1MVQSjH2kac0wsxyodtu+RwvrqRCKoDgLz4La+bUTKahVp+XjXZ4LA9Qf31vG
yDa528fMjWQDcZQEeXATnxBdYd0/xaiLg4ejcNzNRRxdwK1WO0rJF8/ZmIthxA6Y
zk1x9SF7G5zJiBku1N17p+oxbOLtJZUDpiTnzikLwRKgnvvdfRiQBfoIRZbqvx5M
ZGS3ascM5FQazFIAZr3QsfY6lnAP7NugOVPijnf0sFG26VDe0cGOEkosKiJ+hznW
jfhLZa4tD/eERyTap5YYPqIjMEEbTV+yNV2HGt35UCOsHVM6mRq43teaE5hO8CqI
lAC5o7sIIhvWaizrfjGwNMdirEotEEDU+sMMjOyoFn6JBgFVdpIS6uxveMrG+LjY
NNvcmtCiVPokZf7YFKDvReO15Wm1NWlbQtnYzJLwI6yT89tPSJ5HrHdWaiYP2Sks
ZPv8qeu2gfob2X3VW7sZG+36tQk79quCA2ygosfIedj8ZiwVbEuwnw24o/R1qFGT
7o9iNGgG5xZRMAwNNoNx1WDBuElNk9oNkHn5gjCCJGJs1lnXVeJABZ/aCAnHaiGs
VXAaQAshXtzAq/rx/e/IQ7bye3+1G5r7n7oOqToI5zuMUTWU1lDNXnc8b0cKZmCv
/azVpTh5WMXRXZqO5ZyGVsCgVjlCPLT/0KZP+Vc7ZdPEYsyeXG8uuLXleeCDokBb
lWybyM0FnUe42QEQzAtE89J95aq5WLc09KECxfJ85GvnuFH+UZ6UlSR1AmMBZWmy
bbGmDkVc68Z6mUd3Ls4841qGYUtP/PoeoUB5r597qDqvtxuWKBeHxYpvAH85m8YZ
Yvy33E+g0SLC9GyUREs6eyN4zBvinJOGVwZL+52AYCUkfOnsdYGNJKq3rT70LQzK
a93OkFClR3oHRgiOSTPDVE6lKxnggOnUga4VEuBirFh3lOQepeaRHvz9Pi8kZkIi
rf5HlqKPTFpr6oBBh18eYL1gMJC3LQdjQAiyuOGaReCG50tU2Zc/g9NJV+GvQEnr
VuxUQ65gp5/a3dnw1zWv5AOHSm27pJzNuGG8O0LGm55zfuGiMb1XqouUfJS+zKZ9
qs8Uyu6EPBoNR1kooncWEokY0Dw8pi6ip2b0dUEuzFK7zWDTTz5lR/aW5Jt35XT7
KZfcg0uVwipY+tPlbVcKGY3HpyxzGXWD/EG0l6Vieh4C8PITgBdsSpJHj0ax6u3Y
ngWn27CNB3+X4uVzINhfNnCarAnqugbegoP4AT8Lvm4pd7Jii6yygyD1o+qgrxko
Xh7Csfw+AyNb6vstUVuqNu98TPB4MU7jU4rgvpUxlT0KIkNyGjqVSb7U6yZMgYoG
c287p6kv5okfZSGbDc2QwikTpBiwWhc78n613Tp12YcW3O9j/Hpj3qw//xTdrGp5
OrByt9AwBjlif92FOSO0iiNx6gSVRE8WfaCi3q9o5LLKsLTNaxJ5cBgjxvSmcLB3
YrK2ol+ce2rY7o4u9DmAf/uNiTS2+WTjH4NBLtu2no499rxC5r7lnPUo7DptLkWX
rF2ro66QKDuOfDRk99gC5t+RAGh1vWM2gYZM8CGcTwdQialkj0gAPVHaNEtyYmqh
CXLPs6V2I6YKso+H831H/YFDKixlnX3BapqETLyxlBi2MXt7nRcrz1qZGZICeWcm
n3XQc12Xg+76IpQ1mKznmU8MRV3jZci0kBZOFSD8Hvszr1hZqagnFwHC/JF+RESU
XQw4xN08+aM9rMFZhwNpaKn0uIOdRx+p8EVnSZWAjieya3YVHloVtaZCbjKddPkp
d1d67kmtRqZWUVHvtEsMdJ/t3GCVkBYicYKibOpUoq1c7eCortgL8bLv09k7P3Ds
97h3kS9VAtnVBI+9hHyDOwNhvQ/1VHhTAL3wSLcArXcEQbL45B87SmQb7cGZXGJ9
AatPLyhrq8PuKqjre6HZ6q6188N22OfsT1GIl1k/i6xvasz4alNCdD78BpO1SVXL
6dkuxiw3mSf1JidfLEOu9lEtAXrm626fea8mL1za96PiJ3vQgXbyH6t2za1Uhzc2
Kp5R7ci2Y0KPBGU3FpWXA9kvdx6BmFv25KfyBGPbBZdmxIrU337dKM68FhqSEAsj
hiFM54ComMa5DBvHSkdS9SVEPNbNWk+e+7INHeZnWlljOsSXXzeMJNjIJj+aguHD
gOD8LU+EVTeO0+xMQkF9EdaKstNX3BVqPYwM37+b1nltX2PMCe3vUzmwWgManYMA
KgcB2yz2qfT0Jmyn8pRGdEBeEm94EvU4tSUDIbgudMgQWXVGLW/A68MONzKi4XFj
SpbZVEM3f8kw+AGlOC741cd1nA4wYJ/5LeUioHhtO6iS1M7liDnbLT+owr/NQ3Q9
rfNROYvDkEHrNO9pJt4JuKzRtsrwsPZMeda7cdD2b4w3nhHHgVf5O6Np0TRdL9HX
GBmcbUOFMX0HRwYLMYGFM9WOMyVFp5jhGhCyoeuaktjKwXNe6mbuEWr1Ydpoh1CJ
6XBrEx4eIIgE4dchHkvSJBkKQjfQ9pGCCRV3/Yh13YSECmhrcpCrFVSlCCWvGaVT
v7Y0W7itWRC+IDjh9MM7kM4bf9aVmIOiiQu+ua7Qzk6ExbzLf4U5+Z/oYCHdZ3nX
y88CpMzYiEQKaf3SreXRDNn0vD/6Ph+0d08Oq+uN2Zs2B+VZ75Af0cry1mFZpU6A
SAnC+/J4b5mbwcRHdi72MtoVmxnxCvSYscCu65pSqbQpCFiHCtSNJ1ff/k/kSuh5
ftTXKz7dcJXYhp7ZpXC5MXinCL50dPR7PHSTFaSFI5ScYyhvVjWJCX3D7C7aBenT
D2ey65SRanAxMB5164jH4YD3y/D0DEFc0p9braB5WF8Walr5PEXcqeVUPSSM69d/
X/iDLmJ+/jGfXSXeqboeOn7QHS7BVQGegilfkp3U8AuYshG64Qdt+44d4+sddg7S
lgFV/6WoVGXL/I1DJmwB/C7rajoUOieZdzj3jhvTZXmJHsHSLgR/LlAEbrAr1CY9
wLhJyfY/MMWmFAWf3K1lqfuwObuJPHrlDX6wJ3+oNCvnHBmxRmXMl3NdsT+96jBk
3e5pDgrEpOrIlMxogoIi/qqbZJwUbwsOuJfCGuRttDZ057t4oHh3seXRhtKL98wd
6mitb/ipBPiQ1DPIqFOv/Zz4MMfqq/oJj1aa81yn2unLebyNPAG4mact+84gJRkF
ARfpHl83owDPyuSuIclpsG53aw5yKbz583wvLrV27yCtvM/URlOGPw6iCB+P81Ss
XkOHvc1OqW4Eg9uAR6TMZawU/f2KGLrviEKKdqzq49eNcvpyPYrJ3o1DXN7dkVRE
3OnGnaiPWtN8E0rDv6AJVVNoXrpbZPexZa+badS4n00CGjQvMIuTrVSO27NTwUUH
CZRXTGVyNcWsueS5m6OXLUA0g48dyfKLJe7yRZISJJl/k6oaBeX5q5TOXuRaS1IN
hoN+gFsT+X0c/MkHC62hhlWqKU43qOHiHkmzP7HvUIkQSwPhZmyUcbZiWXsmtTYR
v9lwBf8mayzipsHOs6sbaxXzxs4mKR/v2RiQ+VKm58hCpIVsqPuISG5+AcX8q9XM
JhaQXnjJLdIRsA3cKFbrobTc0Vp6k9mYd9gTN2UwZWNqBAJ7/OQesCZOTqGs7aST
hzBlTjMVWB9TezFTKg20ZRq7q9NNGlTTVdcK2ZjYmgc7RQclgB0DayICBi/j9Pf7
xX7CHZ6+edRecRbgWc7RYgHjDPmIU/TyaHzQBGavl4l8Jje2ouONLudX3PJwQqWs
Jw8m0ssDczkxYDr/TTEVXBhbauwxN6X9D8VIJGct9awFsXEB9qyPT9BEsO85syJa
SbZ6KRHt3TVqgmVP5s9bA6tRUPUtoKXRHfB1yVtBKWvcuq7uKugsFotd3mJrkfVA
Rppcbn2GcEAp4K4nAjUlqwpy0AorZdY76MU52EreLdvHMmK2hV1pgkyfgaBsziu5
RmCuwRzsEqy2UNcvZWPsF/o0Gjbx0f3p9SFUtQ6nEj2GR06G6FpTbU6zTX+JkCTz
LN546D5rHCnC1HYRU/6H9HzENEq0XNXm2RASWlnw47dop2w8D4ef5v+5pU3mGB1f
wxgdnykURdmatgKWvWNrQODfR6Dt2fy75a2513KOy1NDRiLPzbzyU3pW8ZB/jreP
xkkGRnbNRHrSHIjEsd8dkLX0clnZaL7fkbPPmZdNn5QdqwyFAZHDfPRtJ/TyHoFR
HTFADUT0dpzcUM7lR6QuqdHBhUfYmVtIw3E2aSlbqygd51YEDPo7C/qEYH89YWxh
fNKSD9xDXdutmxj/eE3qq43nyuURdaeoMf6u5ylyw8kuafjHYkoadzM3pp9s7Xdf
jI7+XLMTQPKQlCwQenTNdKvmcinQ7m4w4XAXCFwYyl/JGTqU/1DXX2Vp4diJXDUO
m1e0OUamWHnNOELtD0kRp2Gnro1eLuK0s4XKTH60bJchGcRI4tIzOsjbROEH2720
zKpUj6F5zAV3RFfheZhsjlNZfKmLW3bjD/oJ+NMbsADc4ZVG0BzM8vVSYHLFNwwl
/ycDzldZCK3FoOtrvgCvcZzxjVWTUWfRRNPtJk8052Z22y5cDs2fmcXsRmAvMl9B
IhScov0JsEg2x8pZOGoULyJkuLbrMgRu7lSmpZPZjtoUZOcuMqYdoWOc8PdI9c0f
m/jt8svSjhw/etAvgHMldto4Ot1Tf7aWqJf16etfwSA4LTIPQhXqzLVDXwsN6Is9
gIZbIBMcJ93/iEtYIlP7ESCyZgK0p5XzAvqZhywiMamNUVegcEMQkINNZx8rl5dJ
9y7EAbHRuta0p6bcAx1icoB8UMJnC3YHw+12zygL47CSdyC+PRkdaH6giRYi9gov
j4xH1L5KAPZAn620TggX00GnHiKTG3hkkDXgq/M86doNVPpH5KtsqoImqZo2PYg4
vfhPNn0OcngEfJLkaHKZDydFqKevilSzpdadIFfeNDELVCyDzwlar5qgPTccTjAN
WJqWpp6+EXWnSTItcn0nETqYeIzKELmRuXd/ylXP+CGucVAxN9l2ip40AtEv7KXp
NMEAUCHn5uGz86AEMg5mciAdc1FUshHXG8YvBbRqYPiYa2Qj5gFX7fb5YnvoTYLw
Ywi1Bftkj+nMHgiq+817kORt4WfrXjBYfrXpozv/4/frlBUNJa68x9XMdJfAqFNp
JOOm9PdGdphlWuZYlHORN0dWQhdK29kwGoFXJ4RVFwJ/o6aqwhwIa33svp5t+FWU
ubKePLSJJByza9kobdoVqHXFAHxMtTWp+L/f7BFpjsagWXZlyp3NzWbF1tgptnT7
MZeAi9GSHVb/NDddLe06mAN/JzaJq5nb3k9Z8APPLP7xQ4aBS5Eohlh9OeRXzDCj
s2W5thXfBcqjwtDWGrGkRH3uIQ4UqvHdj9IP9qatyCoWx0xM6xIPBj1SUtdxxhqo
PO3o2NkmOKVSLjUszhuP57d3nvJWociwLo0Iwi9txIbSyLDiPNienEID/asxUzkC
MSEZrVXM6omewBCRNLYcf4HMr8keM4rLgtu8NvbUZNrQXcrkLGsgK5xZTgKMD+9b
puen7xXgQgcStYOSTxzSyBOqRvhlqqnIoC+mFb6ni8IOtWDboWOxJIcDsluZLHyW
LNGPascElp5eh8rTcb+Tzl4IWX86bQnaF/rMb+nrsb/xoXkCjYvwrNoSWX0LxgXW
AkGGKK10Ef7qyleMj/NjbIn+0fDgWTWkNcxjN5Hfl4NIdoHNMMH12tmpU3Y9L5Uo
+kZSp0B38hCZg0gtA5vtIY9eUzQJEd6QpEKSv8rNFeThm7Xrgozlpt5JbZTz2Sve
vP0ElonzXti81M8CFd8RjTD1GuoVXE6tdCGNOOnZudbQvpj/30JfsGOl57d4HXiQ
Dv5btm5/23GynNgJxPQtowK3sNE8FkyLVQ+ykv0kwA22UN06e2Q0kYQnWGJCVTIh
DrL4cGwcKdflP9wi4VVaxzIVitBnHHRq80R6EruBnJ3mPFXMitW2Yhrvi15kGcLB
LvPzDyY889Sl5IPJZnX31w7Z7W4u+df0Z+L+BBpHry2qe+nMVaiWIHTOSsxhWqZ0
WuMmE1bs04bQp+YkuoEc89QCatctOjBjAmbzwSPPtk+bzptF5uOLb3e7MmFc7fm4
R4nQG5WV2ytDLF4Qf7XgsaKDnFqv26pEn41/iUxPepwJWsHQZq6qD3OQnQLAOnvk
U09+e9Br4Gy573lVp38iMdDLpkTECbOR/Ua1JV1P9KrOA8wMhY0Pdiu8D5Wwh/di
F7+/bY/24UjFC2VzT8AfsT0JtyH5IjeLxEwd1Nrp9clvj3blr+mdRf19Ry5KQJ0c
Da/00MFr3fgoy2eV7GLPOyqqnAQxz93Tgmytl2mpXooJFaeRtv64W24O9oDk0xkC
t61gYXGXOpvRjlh06OU5fkUdoUJFxUxsrfANgIYH0GgMYWp34GdSuTi+UEqaTUfS
rUeQgTvLMyRcAjpEdckvcIo8Po9clYfqgkQ8lYhkCv/OUb8YdCaa2V5922eRJWdk
/F1T0bSN6NYWbNTd8Q32WLCWarTpR0uMPdHubtS+CRMWKo8Z2i7+CyQr2vylX/H/
Ua2UZOIMwtf3ynZX6hHemSRKJjxFHzExBCkvH2W5LVVRaZHbFTwtI+mFfPTY6ULG
76s404mR18xuYED21xSQvr6YLtxAhzQ/LkyHug1GO92WMuNH/6T2JChAaD1ldYva
x8mnP2gjq3sKNwBAOhRC3uhY/eb2pmh7aL8NHRF9W3TbOXxyDZomkfzH71t5fycw
Is3wWRZIL3gxSvLjskXCdj4VTyb+pLqN6xa6aN3x7vxVFQxs7K4+9tGgo/v4zBQ1
+mMpUIWlIbDD7pVwkRoi5J5EnhhEZVci/GlGccb6R9pwl0z60kDox9CPe5HT5uxs
bI2+FtCHeBGDiJZoMdKsUdLkQSfMT1cY4sdDumabFcZMhiJW9FVpTFkhkmDyHonl
LGOdCpG+ylwpbkc9q+eqgikMQwht+OpbJ6JejPWk6REclpnWxC1IDU3cczoUwx19
eWiIEGMSfqmmziv4QmFPU9lSDZEG6NDxrTWQrjfvx7MaHI1oXbJXAXo1XWIO8N7m
i5ZDTx1hynJG/fLz1blRUY/3h6qMO+1eq56lu+cUlZR5LFVAJU6DOwvNewgvK+IQ
FwhlPsJ4L+YB0ceDawXVbF9sbp8WlA/75VXWO0vHPz0g+CavybFq0Z0AESMehYO3
Q6y18nsifFqaCAAcN6uFahSVNVy/GbHoDK3kEhLPNIViojA0eG08McqlZ29KDt+M
w4qNTrC2fy9oINbFXgqBnBv/vAneXeIr5AmdLo2L5yvSLn1kkS1odJtl117Oo/EI
ns+slRIRuZrUzi2HV3ERCEJBr+WrxsBQoL6seURai9EdklvzA2LGU6T4AQyp6NeQ
OL1thPnXLkxtw0+Ko3zZvUSSWyqWoG2qeMcEXwcznkM1UNc64+5vpljaE0ihcI9B
IqkTVRS5PN8OU1HlHKnmfbCo7sxW8wHZr5K5jdOP9n56tmQs3q9QOiOOhzHTwKlj
Uew/pXPpg4v9m242Fj7HuoCOIvHq9tHqMNCilv8OWK8bduOhPB2cZxwjHDjbrUh3
HECwl8sJb0tPA76rbTUZhhh9sfmScPeCU4UKPb3tA7blihr8WsAo7FtCIE0DC9tI
EXFfd8BQ0u3AA0I2J7e1fRDisxcchKqJbf8DHJwp5cWurQR5f9fe6l88LfSzEZ9W
fkwznOQrTLoS4yQ9ZrIy5bxBve+o0zdgu5KYYanI4YIc6wF9dYDrwYbNRa0ZVkC9
vlIGc79nNpBt1h3zpu3BvEy79knrNCNOyNuDkSL0FecjoAgXRdFPNB+BgcYHy4ge
Nsl0YTwXOAaHLr4FealkE3bO15xixxFf9+CrbGDi+z75BOtfIPHOzypGtmFzAVYo
7DR0zEpDVaM9iUz1AaFE/nooGJS9ykUcYbpClvISSRvzZbcJglMNucvh6PI5cUw0
DqPn2cuyG22+w7ADi2HOg0uesmre/kbnz0YtLg8yKgBAKXzv2AaFpUk6W/wtNUz+
Xie7+1ipuK+glK39D3CU1wGgNyogqwWtuN/P/6XUMKDQOHDLYGxud7ASErCSXjLl
eyLIvyTMWiPPEHNjJV/yYHe+Tql7yID/9NeKfyZxyHDSdBlWxDcDYL6FI4DWKgfr
Uk7eNpsrWVN8F13rRSZgWtXqh2h9I31xHGIdgSbs62/WYBrMlHo7gfIj3mGrRORe
K5jBz8AFuhgKOqIf1CDrvwNFbNTs0Hf/TWYqv8YPWjtsZDS+wwrx4rl8U15praAp
ITwY25ozkCspIxmwWlK3CFAMBSSvU9pG35PyXq6QSTwohb4PohtDUX1jJkaW87Lw
ZatySRvs9GOI2Pu/0vO6R8+JgHM3xWPvQG5i5XLS4Y9xG4QQxcyp34Ag13tEf1dp
Mx7Mf0rV+Bdb/b4lVLHT+rqBn7LohaZluuFo4DUqSSyvYCm5/kAfIEj9FBotqwpc
aRFv7DIoGgjaW6a79l7d35VpOR7kHV/vrheH/X7SlRg3I0FVSfiN+1/Sv1z09pt5
/z/dhQmnb3C5zFFhGHsOinE03vGOWZE9YSh8eJ/IJn9y7d7j9DzoCA3QoRoghscm
zDYjzwUxAfM2SfZbroCXF9dlGV3mQ+/B5iWbpTHni5xCS/2isTT3r1nqhejXE405
dtl8Fj1Erh++7jsotJLfYt2Bx+NF+3lat2pFFFDLkORtob5bwox3fdAPnKd/ArYv
UtSpQQl2bva0bpCuLzJafRdyeWQiCexmf0xeqXwVkKE17aP7pToVkwBgXNT7UnTY
gD52NUUxB+2xICYld3N4b1b8v8JogUXLO5WbPCLICIg1pn0YaDb1wS4u8CION6vM
1lQBZddQvYHnAaqVQJjUFd3/WPi2XerRtSM3D+XoYLenUm/aRaXXEa1MkVqUr9UB
W3jK3ZFJCU30Dvgwklw1RmWO91D18sUGsCMFZ4uQKPbcLO/xmyzY8esplJ6+HsvK
iTfy2wsTw1J8UGtZ3wKs+srgJS5HAO8JKxotHaqrqgFB1+mRjBqbVCDbrEKdswWC
Gs6CADx5MS+SSbxqQ6y2CHKe+z71YAim7xU9TXC8mnr3AQnp4aqeWyQqw0PYL9Nw
WunWTlX6mCnDXzw11Sa1CwUTST8U/APUGo4Agnt31Ccog4Mow9N0cRLcpTyjlxL0
TsBfnca0t9Ztfwikm5zdDJ6P6NrmmGCkURxip9RtvRzg1B86cCso5/MF8BzNkxLO
n8dSPTC4tXtrMe7BL0OxUgnCKrPN+QPudjOnvOnWCyD8Q3DmpKE7PBO19GGVPHlP
nvTLZTzlq6Dv7pT+QwgdLYSY6KS4Lkgts7fRYZ4F8s6xObsGSOUNtLzSCo21IAHK
SrmYDfFtCUUaKG6d/KeNGJSVv9W8ZEE+oc02RGrDpnQETZLpPyU62NEx1s5EHc6N
ugv+KVO9t4eJKMEVik3Kcnmc5p9cGZRW10C3YrBiieGgrJteJoypkUX/4eB+l+qy
QFLKLgIbkQUppmc4EHjm9XtglRwlCpZkwfZvHsYVLH2Ih/rdbtqshfLhfStBGls3
NVHtKzTSXhUSYyKg/uNUOesR+1JnfljRPlslDvnG77cJBpagOgWi/f/t4ngbEqt4
CrBa9bHujet8n9EgAg9k5cpnoOK3qiPHHvyQqvQLpRNziYjScruPpbW6udNDV/8E
UNK6Z8zgnq24qieZsSryajE2ZoT5HVpBoMV8kLwntvtlvqYkFWuDC5af7l0QK9zS
nbKfDTJ+6G504eRSrhK9CW1LfYyJwiHChhQE+eKgTiWAWQpwYYWSJ5RSJdahSYuP
wIrAJMqezxgpG5q6582D+UH0VVFzYsCq071z9nVZ/WlpTwBPlFbn/iHMN5BpRvO0
NMXqbe8hPGKDq+INz77ECCptOhxZP9EHH+1UF++1e7G/w62uSXtLBLyOsCO8CyyN
3jGt9EycMAkF2wYcL1oi2tL9ESsLI15PZL5O23D0y3vlrrLdFg30FkwNwFt6YtfM
T68uscSsfqc7RROwgi+h8HgY3Ah1UqNutwXVmhMbuLZfc0BYJxLP05CokKKwt7Xm
04+kwfk4RALOvyEaot5/zAHYx8711NOKsu4pZAt5Ig/PUgfLwoHZPtC9YxMykUQP
xMPh9JmN6yEP9zsWKx4nqDCFEX+Y3wae8tyJu6InwyHhaKYDdhgoLxgIU6faZYaF
mQnKrz2TykEhTsTiNrborh8QL0mWc6zdGSI9oYnp68mz5L9gupaAXDNz7tC0AZHc
EtVVjEbYaTcf0nFhjhzHLTDxKfPno5irslFnu04aZz/lIoFY2ZeLWUexKoZogztZ
BlnYDLfHKoziK6zPKH/vfCZEQgt/sdeIXIxueK+RJX9ALUTWH66K9411BJCygNwt
o3PIF5UpopmWyZNwY1erd26NwFgGpymS4cKvzKzPO7G6XLJ0AGxaYFdzzt6eHm8S
APCp67GJerV/Pkp7R1wZ28Q9eXNb+dbn5YSpfkHP3eIna+DOKdC8/q0lMaCOk/gs
UQK+zlKOTFM9afhfUdMbqWXG+FPZOOaIpilkL6eicfjCqIR5Gc8/Nl4oljdAK8cf
7mruLoo4uXbmWuS4z5zJOQvVomiUqoZk2Gqx5m2oYaKtxljD3Xd9pnOf0Eqd2nqm
RznRSCWXDU/Y/qsLz6ue4zhO+Int6lDwmzkGU/6ZmVP8wHRzGOEI29HwlxXiz4Fd
tb1Ls1QrmUh920PJePuOTxSsE1TKxs65BUB6iWYWz2u3X5p7JL+SCCHYwS92iWL5
jqzHnadPiNaPmT0UTm0MUn94jCFnhzGl8bUU0CEihkCxlYp9MSbfE2XjgrJ5FEeP
qMwrvvZ/9UaEuqKSau0HrpA+bdlxU3aDIZEgXO13nAOec7lO6UlzLM+OaL+kEWzu
rd49dI2OCMQB9+OEi/XNstsNjGIGnxgynGrQIrdV0c3i3eomr141exfzLAx+cBdX
PtzwIXMFO5N2eTuJE+2fT3dZyXvBiTe4tefr7jjRMtu9q+l/9tF8Ae7O6e3bYZaD
Onwic/BfMDAs977er8cUDiUlT1b47gVVcXrDKUaxaikztGFTy+67uU8di/VAMLeC
WgqyuQUzLCou2zLuoOmREH/ORUSFkkr5ug7Z4gOeIpki9VnDunRipMjGhNUF6mBT
FP4oqZ6ZtpeGmxN3wXV7FmYP/gnZmQnfFeLD9EEebXjdbcQWli1gvW9+GZTJ+op2
quXz6oKeVW+ivShhMi5HwsiB3Sip0psJkyM53c+ecxB0VzCUesydhr8JtIBvyQxr
8LL+iPujIRDyQkcRvfJ6Fy7QSgbkgFgS3Yku08XCOcoeS7f7fcxTIZ324sB+6p5X
DnU8Q1x3ttGKczdc2ao0QN0zq4VLGqtSNWlA33I9rCks03Uoe0VFBTuVpMlpKhm9
N0QYZwLoqRVXLoRWPJfjmt0RrEZ4fBy6xteX8rV37GL68dgSxyjN25mXifT9OLUG
ycuC/yJfzWsnJ7V06zfSIc7LtAj8H7X88dST+YsUQBidU0jB5LaUIXgx1qgM4tEz
pTypnYWOTyMpEdKaCHq3XXeeRPOhr45dr0wnmR07991+c9moe26JdTelG97TMQxy
5uHlhESNOGP+CA7CqWqIUlQd4Hui+O3pGFd62OSv3NRCG3EyRqxCDHdn5FCbRUf/
I7QQAyoaxpDvfcjmhf6S1Cedldu0G+xBxhOwF4nmWVv1m73GlFrGyF5IZyKd4Y0+
qJO/c61Grl783xkaKQGTc2OAb9sxK5AfFK+2fqyiOjbroq9T07RLV32BTEnevWQ+
9IwoD6LnWe94euLLzwLIyAiMK4bWDZavFjsrRv5AlUVOAi/7dmQmClmL8s3dhEGa
KAJ0fnJE9mrqGI9M9YchnFfyyIYTnYEDpbOdkB7tanHNTE71Vvm8bBQnAJqS2Wkt
Nj66K/Aa9gA7z8Vi65qMcvrkhJ8DSHoFY8HCcdEkAhFJcd20dpkEoKzsA3LcBa73
uZWEG9o8lBVooeX6lEO5P/N9Vj8KRZWAt0GtlzvWm7AoCusrv3al4hSxr4851UJW
pG29M1jS+5QD6yH6zPyNbMvxuMEIz5JXLedGcZsywWVYRTa2rzFm4CIBP/8LQViI
y1w0ePfYAw2Q9JGc4rc+AZoakfvrszkBDdYlHgDA3HPtlwjwEX0+LUzmxdUb7tpn
oM8vClwXBGGbq7kWUyl/ZvkIkIc/4IfFpk0avWZd7mIIXjhQLZRLF+alAggydbG8
PGZeLeCLbATHA8ofwToTRNJ/0i20NCK7q+Yi8ow8WEHELNhkAlkNFkeqcatepDmR
VJIg2ZvPwXzqrafa7CA1gSLv0ndXG7DCEJurfpCGcTe9FtCS77IHsaWwdbb9R4BK
kjDBtQgAVDMl90gD1kLr/9znxFI4p2I12sZ/2sV1X/wBcgKOl77iMeQzJQ8/KtYk
0/XrMCczmIq+462C+gMm9mv+Qp2Oo6tjK2XCVGGzy9JtmsdjVKAvt9LpGl08buoX
o9Rv+lhZNm0qJreuvYA/+SXhpHIvvozheBzQnTeu66MKlwfjSHSq3icB3E1peGic
ZgGOqis3maZI2naIJJf9Nzgx7K6UShcEF7FL9Gak2yB/71ArM9F9IJ4kacRW5ecp
VFW/jIgfZV37CJDVCa3X9aIg8vlx9SBIotWMQNT8NWlrR9ehbCesudEr7nvEPa1k
Xq/+LdTGBy45V7IjWZYuIHrNjOLhbHptbrnO2ORAIpKPWoWoyBUz329mrDsu+RVw
wjxNIOqj/n/c904HnbBGqXNIpwy9ISemciZAAJxtWUsOBRyoDpqDG9KE0oxObT7N
DpMM2MK/JDXNQpVoHLSyGkM9gOcUh4SrIdWvS6bgsXoqMkreA2uslYeHKRTfF2r/
0YAIhdzrkYWRQ7r+bF+89HdQfOlPVZxIhgxRknJfSlVlQfLzpc1Lu/fqKqAxHvjS
sc4MkQ7cvDKemBYNt93aRT8wBtd+IEHVKejsQmBAPV2gQ69yuY8JB7OuO+kirUnC
sr/l6T3JEsyccCyyobvpXby3hvyoSQiLa686s+6pkfdwt7xNUDS/RkJKh2jvCdA1
0NwJDeL811gd/cAeBOD2rmY1GQgqnjOsyx5K8X7KdizXjYx9yjb7LErJoR356XLW
d5AjJSiHJyS15shR3qvU9bGY7bZiUXUmpCNVOEPn2ucGKu2LNtGapuX2lV0/h7Vc
wrsu+k8fdn7MdHKD2qVhPDdN15QvqLHqY/YIopwEvaVB48TzKCgagTtv13gFPSNj
Gq2gQawoxlcH8PSPzjKLhfA04GUH+HG10+zBGwhXwfCgG0ZvD4ytR+qm7t2Kw1Kc
8Mx2sUggSJtu40SWTMsUkPt/Msx85hI8SYf29u5+jVolhU5bv8wE5xQRUEEDouC5
wvLDapdHA4RxEcfOqF7AYEyZ/Pe2tw+ghQfgYcnXCTbPVsJreHIt1LSWSlNx1LFX
w0tN0UcsM4WzPepZ7/7pydDaNO0ZSuQwBD6M8BJ4QaCJoVTkvHar/JIU156S/vtA
rdW/Hya7n4OrQi5rNE2Asc/NtqAcDE7/56Uxzn8niecu0a6Ssb2W7ttQb3XFe9W4
ChYumxsFiqGV+BA6d3Et0EZhBbyrO32v6PmqdSDsU1H5RT4jrxHgFdYWguQmZYkC
fDmkyZxCXj14jSJvwbHC3GGaAYobvbLaO8sgurMyYcR8CFqw+7h19mC5yKJUq8lL
hdarkffz1jN7CzM9FO9JSnHTfcXFTZizIFkp7MaPEWzgleDcuQPHzqh/vHq/6hgF
QxaUCwXHmUcQ4v4GX1tJEvprNkGa/we5c6PHtOmVt+hFflWn0FQqWE6LWKxmbIoq
APx1GQ5W37paTLYtEoTj2j2D9yg9TJcRfTQdBLEiz7xrzFfkQElEcpYaC3KFvRA7
YKEpDAoRf11oCbB9f7Ef52vOmdwHKDxwIH9vvHFgImbsRJLEEqlJX0u+86thzE7O
RzeQEyS6iHxHd7aLIpsdeav4zHT2OP4tfeJfvAypG2bek9J4XFRcRgTf9mufvVnB
mQ4HGL5vx+PpH7knhZrIXuscVM+Jy6zlkuxoazB5qK5qyxkqEfF5ep/8nkpjlzlA
DYBl2irvMFRx9t68QSJY+bqhaAhkVnmQt1TfloupO7pmo8biYdIV/ti/y4h/DUks
8GwOB8OFhaDktOIfA9iRco+XIeQIYusDwJkFGwbvFr9KqJMIXRrcSh645BwDW0Up
uEMplmgMAsgDw8LZqs1MwpiKhO7HpMH90OMvIJzFxFyhKWZpmKRL7GeRYEF5fvaz
qQ5b7hLcncrh/o6xmB1XcNpzdWhiYR0V55BB4WzShO5L9OwoKkeBGk0J7UCpKNvU
rMv+Eow04f2UgDbT+TTmLo1pg9VqMXUZ4Lw6hmggJyCaH1xQu0aUQxPumpBbslTD
cXa/f+L9HNn3jhrM/4RLv4y6F1aL8rSQVzYWnnoC8pswVJBJ9DOHjDU9jpcyW66y
t0O/k/VrdLZTbAiYffMvbgoaqPM0G33qFB2vZUR1SgwZCzeAEOgAqqsGwjd1imKa
UXYYEQmS2GIEWn6vzAoSVDnMrJmqXC5dDVLsxkS2sJWZrTGnbiTU++kg21EoP5Z3
au5pJcpB/syqMKxMU0RTkLCBnvZhcD9PRpcD0/FcYBrlBeW5gwwwTEtCOAdYNNPc
AMRYQHUEbQCffFbQ8tMN5uKW4v+7XSQQyh8Cl0B4uP+Tp3FcT8JGfmylt6nswT/W
n3hop92h56yr/EPTj6ZIqMEvN4OPpFCUP8Y/2tCk+deUI/3m5Pjj+54Y62P0Zjhd
skO1gz0a0+kOhp5UlbV4sVADFQSwUqnE0sytBizkeLMj4g1aNP25U842Mv9o1bYV
8hKam2gPLCbImtTt+5QHMgJeNobkam/8vNiLo4GP9BYzH8vO3bcnq6u2nNJtHgRt
6db244zalNZY7rRcaRLsFOqDoRAaK/GuqfZGx7kvp6ChIdxatqOaS5QaCjjt7j4F
DP+AyWLMwSZB8v2vJX1FNs+uRhq+EhH2MuPkGxLNGDcWGYRE6PczBXJuefJEKreM
CJ/CwNuUujKKdg24TJBix6kM+BouLDpPUHW6jhu/KU37m+8NmVwCljOPo0hcuPDt
FdodFbN9cFearwBdZALzqZ1wyzDFXCODGpXERUy8AINjbHhdJYbeKFFU8JBoa62K
EcJUVAVuzPthhdD2AWlgOJJtBydAUXRpycaK4AwPia341WWuVuoYC2QEY3dvJ3CJ
kZY7/CsQ0Zqzbz/7bxzj7e8kBRbG9mehLHmlW+f5YkhepSk2FmiO7hWl/zA77CK6
ASd16nnqNC/dTjg3eTfvDgOpxsGqh+NO6pjaNd7FiZ0wNNourkzvKhAQ+6X8QQdS
XNhTyWIyWFNWlACvNBaxuJaGeQGlpBWa57OYC2mDdkMSI9bfzzEmPXL4T4WyNJya
Pl/TO/QSFAkwN745xVaYq3tsTq2fKucDqhW1o1zxpfWyVtcIl2NhwCgt1oFTNwIe
a+RzuXcS/6RnWDrDvjcTsIUbBzNHAhYuu3YRxWXFugRUpK86KZ69tdTyZ2lOzIvW
j6DiFx5Q+4eg2kdzlazv22G6terpbuZHiIJI7tsHiicbilx8O1ZGqxPTvrBYaCuG
dPmwvUTjmTvj/wak47ZkFMs6CvSCwYTWp7BvJUPUi3gGa/vVYnidU3R6iDaon+iw
fIIYN57jm1+C/ITmdkbWuhUCBPNoZvn4UL4PhwLdZmcCe5cxVFPHGZR1aBuV7axV
glvDAD1aa6rzhCCE3niPFGdRDBVXOOmWiSl4BLDp7diZn+cKbLme3IYAizFz00EW
Ija23LsKZu1n1IKkgjK/Kv3cSIQup8offYaHf8CqGglYgJNv3IiHwtIGziH0WQPP
HhC7XUVOYNZbossFrcEVTAmT7N9iy56jHoEGATl/ajE/EQcKRhh1TLzDeTLx+XPt
oYS5ia7Qnl/x/ioZ3RZCPDB6yX5C9mp3Hpsn9m27xxhWVbvpw++rcaKdzEmHEsVT
KGvT8u56D1SRQRSdObiuz+KS6s8kofeXZJwHtmAmWg/dILxJW3G5C6zpqdfPx0h1
blZ8xjUfDKoZtSCzxdanBTaQ4SmVmShKBq7AfU2UU5lUj6p6YFaYfL0YdkMGDb9F
1Rtta7xHiOefEavo48T1ejO8ysPYScl7l0QhzL+T3B/h7NvrTGAAWMXE2AD1tj1y
1v+eUO/F6c2O29603+plG1/hNsPKGrFKaD+vJ1U6QgGh7JGL6/SQBtee9FjIJybO
oqi9DEpcKJ5/WzvL2/uc5HODilvlfTUNzLAJV6alm1ocCGCYJCc2qiJGDuIdLJdv
WfCbaq3L9dsbxNd9m5vUwF8gYDOLu3vUeLpT+Jwkt8OtzaCkMONvC+P0pgdiXVRZ
ryPaFOH1JmDemX/of8vC8krE4ejKXZ8TpG1LjYnwVL33jUtE7YqZ97YIAJwC13Gy
IETph04rnc8mrgoEw8/YothCmGMyj3whaIxUioOWDEuPchYzmkSSQdDSd3J0XF+j
K1a9n9tmLWHYCFwKCEnOTD7xgkkxeOp//cmMbKzRZnJFWpm8mcXBbGnM6AkjwoY/
c6NulaDzVrL/1kfV/JFnitZVOGFbr84z36SvfqB9ysWW/2cmr2Z4vyUT1cdRfGmC
XNox5a/WgOFTvmUEHcOqdAdm/TAMcofGYDrkEVvPWJwEg5UrUhE6PKzUbCgj6j/o
dFGCloQsfxUiP6SkqcB6hbTozKPg5y9HJDokJ6TznIdHIhY9NlUwtZjS3vTFLXVW
GpQne4czGYmGx/PPuRQgi7YNLaGvC06x3TSnxarlxikGRAbHdu6bdOr8oNBa2RUi
RDOfubE6pMedYXZr3CfYTMBgzhBV9rJbqR4si+YFen8uZnd382Yxvyjfs2LJEuM7
AB7vdQ/8+ZXhxyDcqJ6vv6q4hjqXRgHliLvN0KOPOVFieOegGpQtTbS2qbRreqb5
OgM0GDmwDMSmcRo2dsxX5H46YEUc/GaYpAfDqBR5KFy1I4F4DFJh/xEKdZ5Wl5Ga
8DbHATmP9aNisHMbwjQNFgR4szm+Tz3BYO2FpKlGM3ocyrwZ+HAFfczJOcTCtPNC
RRjipl91jdmVy2RTj7aYcqggYRlL0fDsFPYUdnHcO7Tqt1lwIUdb882CtFBt6/K7
Siv/wjfrmueVI7vXuUaxyU3ZwE1FpU2zeyGaKafD90qJgpHi2FID60ILpuAl/Llc
pSRzf9o0vhjYkum9vT8XBj7lEsL/xbncVkXmD0Z+FSKTcbnL/sV+NizAxMzno+5+
Cs77R/+Re13cMIa4k30Tm75CjZjhXuFq5ZeTAS+FHaABSJZzwDHYKUSx0f1SndYg
rHhnzRDaadfFSpye42O8B7VNkzG7n6f4MetECLGYuIfQ07TA8Ai4F7I909N1YB8o
Q+Y8P6OOK2r0GguKOvCqs3VU0v4lc987nK05hNBgJNAKfYf1aIbtsSGTT5dsyjJP
cLegs8X95eRKCDMp8MYpUngtsKemLrQDmA6gPQE9dXYhSopjiRPRqhU+fHmsFJbr
EpndOaKrs1FbfmXRAK3OYJkG5HMk/6w1UBuuFmotsYIKJdnB20Y/iEzh/xUUSblU
3jNvMQKeSvvW235HWV7fnyjZ0w1o/bAK6ZuA70p6vwHvNBgWtRXy/WPMd2H1w2d9
LIgj/eHYSqIOgRdSFj74POMgdi1D/EsNg0J0CCXYRqnaDcwqSCPVOK3fEcd2qTyQ
xvKsu+F9ozozbDmyE4PFZuHAA802WdKgCy2xWzd9/vWEd3Ffx0MKxSQ1Ub/s919F
nmTVe5IexFzWw/l9TlRNuOL12oXkhyCDPXoKulNbrg9IkzSFTT8V7ibiBrYuuruG
azJc240pol4EbIdXP2LzZkF73X+gROX66b9Fd7iLFk4REDEXvBaqUZGJ0TYwxmhE
uofzxiaTYORfXHfcrqUuKTjYr2trUSUAlVJv4uBb+T3fk48MPJcfsRSPPjeJ1rA8
LMeJQ1BQPJaZp2WN8WLoxiCa7OEk9KIUmAxBX+oSUV4B2qweowIOPzw+HVtOZiBY
HGqZhk1Ko9bk+BSjCkualoWoTEDt82ByvdhfD2ZzjkhdgSd5L6Fu3cgGCXJkc/HD
iex01hIhY7CzIk/8xpsxKF9V/e7xaNSfnq9tjl6Uc3D00njjxkRDPqbfKbrvsL+P
2hdUqVI88ANhOz43iW9UR1Rcr377AuLT96cyvhfjAFosO5vFpxgUbybW4RPaRPp7
YX6xbc8ZSF1znwn6z/UFpht9013jdCH7g3bzzsm85/2IABYDEs4Ui9E7A6SLsgk2
Vrfz7PMOHYIC+IvsQCTYwxUZeFAtPAfp0pGI3med6x66O/x+pNPVfAbAqU9Qt+eS
dDh/HyILQjTBHyhLlScmIw5Ij4Y4KQQ93cnO6F4ENadKKVIT25s0qMsqM/PcgXNE
hqll+P6hUW6z5+bMpQHkmJzMB25LvYSfNZjk1yEQWNjtjz3UifL7veiY35As5M9Y
taIXTQBrfw9z7aLKeRgEU0p9oUPbEGOdzeD0z+F9wAp0v+X4z28dNriWn4htbon9
PKqcqh+NFTorEWoT5o7PF6rzp/P+1mHCeYBWKT4QxnbhQw80UjnB57MABRyizOdB
0JOpGQzOZp/3SDFNTTkPJ9i1OfqttSAExy2MzsrtsjRTVxxjMyF+V9DdSWdXfm1L
W0d7NebTZ3hhCQSP/VHvsCZzSX27xwHxBAKf2NlqvcrN8zvJ0moz5HzvmPWMRP1v
zIr6Ak7QnFPGEla88NyDv3XLZ1QUCoW13LrUahW2bALhzmypZCwtyNhotWnCQdjO
xxWKQKJWypHa4wBsA9pxNu7njQWUUvM9AOmpH/sEN+99IyizPcS6qKlt2wbAqMpG
mtp1DVmr6VW0gYQfe/0ga52RQkOtOTyZ5YbHhXhFzgjIEdwrL/Odtnhhq9BWqRdO
zFGcZlG7P99FFf0ESksAKcXB7jkekWTnHqIthSr/0N52p9KMKaC/tED1cdHSdbTU
ZlU95+q2Mwrku1ejBp3S99kZuPKoViatKQe0hGLLKBbAmHnvmeiMOWmnH9aNI15f
6j8A1GrugrdVCn0omysEZkIZjPBh99jML+kQayshaXIQ9nZ5DMtVGV8j+alLt+Yk
MOcVPmxu/uZQJLDtLGZAMQPLbf1d5YV5F4ufxGTWYhdPNGLhBZoVHFrXsM6FrrAZ
zR0MNnmsRUmiA6uK/1F8Gk8/6MnG6sd71BY7SbZC1+KjDORlzzKKadg7CvdHc/Wo
RQ/a2GHv1OQvP5tq69ZKz0SCvzyFVmP0rTbnBIt/9ovb3qrLfpqfi8SkHjzCTP5g
xwijrQvzPDRUTcO2FAwDAROGKL3sCFxC641qBHRNyjnK8akKpSnZBkYqy5G3zxNQ
JwKdQ9Ta7WHvhA5OrbqjZmLVV19RiN9Iwq+n1d0uzDNPUsRXFhoGf43ot1tq4zNR
VhJI+EAyFrWLUC7vOdkXB3rdD+OucXaZt3kvL1NQTT7L01weprY7rTpxAmQkv6lS
HezLvDs03O0iG/W9v3ll9EOFsrCb/iihn0k0KklKn6kSGik/qPw7C+VvwgkeF3pR
8wbDMMpgLIiXF0WE8rW9Gfs8BqcVKC1ytJmZnGx+HFlSrtnYxJbb9mlpxWALpaj1
4ApQpYA2EdSbT7addU4vr5nbQjN8z94Iov7lUOnqRlMr01blmHZqtix5GI5abEF5
R3QTFMI1JCGWqOSQK9kPh+TjYX8pMg65sLSJnjdskjX8VJRgrEViFTmqezrOyNyF
gFzA9+t0o8Jze578+ON7kVvJe5UGC/PW/XSh9U4TkvWFBeKhzWMrPldkR/haWsla
vEBL/y0c8gmXmnN3rH7APwqKEprKoGT2ivnOnGxPyfEX0U+hlW1R1xmyPeIKnNu+
ZRtb8zJOLxt7s3LZerI9Ru+EujI+IRjl+pVLv5mT8LgikdO5pcscUR/cWrb6pONB
xiDez12zz2E1r54HaHTrXK4WbDHcaYz8qRv61Ata6uIUikLEJEosgrTRBeemyhLz
CB91+FNo7uMvzidVdXQMcwgvbvoWHe0n4fq0NFVvH6yY+xpt8Ke0zNdezEizm3Wx
g2ylNdkjqhBh0VaJ2J3eDNws8kCsEdvFE/L9nZstdLRv9om6vgfdEe+ZC68cHs9A
vMrZ3SnlzDX1wZ+PKDbBYLMNlBAv6RgKjm6yUX97mbwAU4lyVxoD06y/7izJiwW3
vzL8vPvYZNX5/8dCQGdHPFIDpDQ14+sb7paoMadloiG0DYvfcZYpR4uNaEsmafkt
pF27ox6NrSRhHQEFY3VC0SEQT7q+SIBy+IuW7XcuNzaNJzkmV+ilrvCLmgVh7IL3
5FGcdzJk8JQsLP+/5knlWvczQk4dMeWE9Iivg1/evPacSP/K8vNb21C8ot4ivQmT
8HmhxhVuj0ArQHpBAaNESn67WW0eKYWaObSBgz6pADIIHAGcSvuU9FlET5P3nNM7
hYiw3wXMC7EOCr7oHYbkofZfq7/M1rJUDvNDeeG+9Kh6a0KK+Fl8pieSCBUCDsSn
Ebnt6lqB1yRiOv3fqZmRtMzkuFHbyyJz8f4+z2+DlRO42kjtPzQNgcQaIBXeFBZg
dUTNejMG20WmxIXN/biBxnStsT+JPrJ7B4I4Fimbq0vAdzr3IZsWhbn/KdXLc+Po
3KOgciYdPfM17WnEDpD+AW7BVzAS4ExFlMt6Fiewf9j8OBSHiEvee9KOsIJHpTbR
EtabxALY7WFxez+Jp/TYauzsHZJu+SaVha3wZD5iQhdNYQMljvE8MplGtIzIK5Vh
jdxJ7l+Mf6UuL2/PmBcfL5Zw7zsH1+bBuamQDzmdzBhMlauMc77+VgHG3S48HVn5
bvfyXCp9Gzooj7aaZqdGpRDiWul/jvtZpISLD4jh4U4P5ijGfOEJEfr224xVh7vb
BWeu/V2UU5cMtrIjPuJPinMUeRLHuq7YBYMwBF1wlVLiyzuo69y4JHJAo+3r/jrZ
rSE98b7gPSJRjVdDFd9NqfUpap4sz8vy4gzOAaL8zVItLez7Z37sCUHSGC+9WFw5
rDgUd+ZdTF+i8DrmGJ4Es0aS9OWtcQPoO5kyM97HS4E9c0NHUZwQE/aHu90Dsh4T
26aIxHUTaGeaCpvTxN2ZW/vzdt3ifWOopt7hCMxhU2ihkffCTxwJEvnrw+/snpjr
8XEmSrB0SLQBb3g9FEiB30D7oCcV2hr7mW0GdZNDUgsliU1SP76gI7BYt0UNHrNn
eiuWCdy/oTiST+7exaariV9+bsFBQV5pIahHcOROiX+gI20Ps+Ja6mUKh0Zu3pl/
WqRm+OE/vIogXbNXtRm/B+SW33xRL1Qi09JtoRQ4t0htwly9A15q4rC8v5UvPGrb
8q2h+NOYL8ZbhDFli8C9LHDcvBO8JTqa6go7iUue4qWt6sAeyDAuY/p7ULb2+QM1
Zz8lXAj8jYab88J8jgrnzhpsLOoUs2OlwdiYo+fVgst8phzyRvnwdWhv/7r1mils
7ilPvzbicyh6H3LjMwtgS+okDA5/TwdzROmorC/8CiNnoBHm7RqyJZF6HlHAiMV7
LM6Hp3mJpcGtawMbuGARycLhHCO8vO+Kfx9ydFcvaWiDJ9he4bVTJsoXOpG7+Nve
2oZDNyAWfnI+NTrqg4+xOBrUSO3NeO/VeHKx0CjilA5W18AiUdEIDA+0SCQcgNE9
j7UDfTAI3BbaUCLrSeiZF+RQMWlZaIj//kG6Adx6XRK7wXSaKaufsqc5VeKr6IX+
2KmksnQGMYQGbwv7HQ4IJ9DHt1VDxV8PfPoBhFretO6NKu1zaOsMMYw8IcTGGIax
2wmhhOzEkH1flGim6CDN1c9adhBva2Jpu+3bYCgFYxzvdjXQRqpNzh9r/S3gcslB
XaDI24A8RGUsl3TILDrEqibc36pWRSwnaL2Oju1Zv0QgGv8XuvaWc7W6nhrc4yjN
EJHK5PKEYFh0ZJCjBYlIcaD7A0xxmUROZKAgILB/xS6VN8X8bPtXFHoVQXVAj6zY
PH7HzsInbOCu0fKnJtoDVrjGuVwUaS6R1M/ArN86aLvrEW78nfkj67m57qFjlOL7
FrvbYm/qYezRiPujZV0lOBS+6VtLxzcjNrysrg2mGCW1SpL55RJ/pfrKOG3LSw4V
BBA7S9Xx6ZBFbQTXtXiaszpRK/5Cm78lrRUC3Tic4aAge9sLfhjowUcuYJM/qg2y
0glpGaEhD5HauT3qIcdM+CfMu3jV9CBesWDnSkOHEndfWWwzVtkWtDOhpGsPUjaJ
Lf6FgTAhFPSICWZUMF5pU4PKtZPeSM6dihGayUQT6nESYvSNJUX4fOg7oqc+kwkZ
AHXlTJXOsKKE/GLRa9nyTQf2WbYlQab8UoZjMehij0tRuX6UC4xEPMDxbg3PxIDk
eLib1ZzRCb7Tn6ziVIPe/bWmdHXHOSGnTbVpythb9Y4PF3EESuwRwoJ/5yUHPiVt
WzjX8XP5eJu+7uvm3zsouR+eLhTjKjttbD25rkwISh7LQVkopkJzIh146C7m9A6t
W9yK881IoVoVabKEWmTt49kJ26lrQWhlTQ3SC8HUdX2u3BaRyWqqvHdB2HDb4sLn
BWIz6KNNdtDXFEnHrXLokzVIceRKKoF6QtwXDG/XXCY/yFSVxyMRXxYcEDa9iWuZ
sOlta3foQtEBJCSvz92UOkaGRrPrmS0z+ZRmg9Q0iRAtcmksG+cHOogOwPdiCAKQ
c9hCLoqgaNZRkXhy68A4D7AOlIlEg6QqUDWK2P0GpQLuzxnSUSSRnxL2TtLzkDe4
our/KpKsbIfTQ6Y1qI3e29OKfvLd6t6D8/RA5zz7LYTc4f8pD+5VUdBD1Rnv6SH0
ZeYVAavtP9swCmovDiS02uQU6EWYT6K33Vtzoc/SZJd5Ibg6H0gAZwXEWlbYDwt/
w2ye/Qm5mXb3wKpYKL//CXJYR6/L7JGfyfrJqlHdtgRCbtRMDilyeqF9jvwzSlUN
7g7/SKRQIq91TbWsqPlAcrPvT6byCD3OrUCeewwtiDvjERWB6TCKJxJZYkRtaBDw
j/7ZJvdMlxF4K4DGKxQgzywRRA5V5dT4hUNDaJVhoLd58IzO0umeFToKgZVEmedd
YmNppM2D/rqKC0HPfZqqD8a96/v4140dWY/oA1JQByZ2mRvVULzrBV/7wu4okjFK
2uWYJjRYrlf6kr6Ow6p/V3K0gQFtwiE7fWYRyIBUfSHDaxiUrMZ+q6Z1qsCBUfiz
Sktj3HR2iNwOz3JJano3BnnYUQSs1C+YJrVLb8nnnws3lndH5RA2l+yX7GOWDOeE
`pragma protect end_protected
