// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:43 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gvXldT2COI3Pf+PwpXyw4XPJYopDuqdfl2FoF66rrYbpCmmXP50lDv1Nfv6whK7H
T/yvB5tya89QX6VZ99RujCJHCS5xIo2cjoFmPQgcdu9lxEliF9QSBWoBf7UyIrFe
q2Pl3DokvI5hJ5WPI7nV4UtmzgU4+1qFzG6zbu9DJfI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48592)
T3nSokL4BHOVSyQTX3m7Rrwn/yhE3r1wnArF9dvgwS+l2QOpgIlHxqvWMz/8A1Ss
bSLVerEa5gdcjXdI59PkYyBHlW5CIMnuZIddgpFXtaeABCYRpu2klXDVqCNziPio
V/g9S9WwNrPAjJCo3QsXpb1BMUhBniZAZlfHLYdX+juyaXP/DCndmM8PvF8s4T/7
7jAjbOXu1z952LAbKeYuOSBwR2JpzGP7tysCVKFa51NMEo0WdTI29uSctFEvaCpO
FpGR/CL5guZkLZ6AOn8gyOV7P94oKIzwmMPAX89+7gTP6Kd2aMk6yt8bvaPLvu4s
LUOEYoE282x1D2jdvJdf+oOndryAdQZf1QISPd7Q2L/ijCZRJXkYaRtRat7ZlH65
rZTfqgBBYZIpyiniwGjWDGK0jdc7dINjkkP4Cm0vOX/TBeRu72CV+i87cXzhxxCU
isKxt3kxcS6oafk9ZuqrjrgDvyLiJ6IpzMeKHLjPpDmB3CsJyyYuVYsJJivurSx0
QuxNCWTbk8scG/4wqALLrA2VrPGAC13G4LJgEu7WoivQ8jm7KyXGofom3EkMTzME
gMvHGxyZPl2cl5TVdhu5ho9zMEu6I8mJRsoJe06h606kjGsMKzGSmkcxFwZLSDG+
Lb1YO9pjZ/sEc5uAzRX89oQ/cymJo4qRhuL4ZscajWA9cXg05TYeCjJ6MiFhnbak
mJuFLQ1roS4EfcvN+WV4QJXA0UvkfeL5r6fcQP84IwH02/gMieMFGiYTiv8f0QD7
nq6tKP28fRjt4DeAg4TbZ40fLeTXq9Xml9gQohNwYdUgvvnsnu48SVmCKQIOM++Y
TSIlU4/veGNgNs2q20Irtc0edejGaXp45tOIumzlJ6e5NWNqOEsZspDREZPDiShH
fb92pO7EOR51lKjRRdHcdkBH3cBUyP0lWIOS+Pr7AWKUfTL31yGve0SJzM4eqxnx
GxbusNaavOSX4myBCCGRnyeStbzrdBMNjtPMk7Mxr5aUdK4e1qeFwhRC9ii3FBji
dstwwmvb8SsWMjTK+rxWQD+PTODa+GTYwdwBQ/Ps7Ic8skl1ez1D7YPWaXdkpjEy
O95w9cyEP3kFaD30oRMnEPoXNU8saGQZMfXL+9vNjMZk3LXlYQnzvdHvKprDJmxi
viQWNI8AzlMaCOjaHylDmLzM7wxmZDNq4uADxQvLRXd53AFI/pPRIzbRE6QLFyFN
+BsG+hqnJ1u/7hXlleU32IkJWBveuveEBwjyUvgECAzw0P2qor2S+cihTCqjqh67
tchgJ8zxSKCKGs2CnH6N7CTBB/Srv08QLzyW1Y+tFEJm10Vs5Ch2M1i/DuRPhfzR
km7MqU1dpeQWPO3SVdiAffWMfAIN8OQiz1fr84319XW5rssYDVdTlQc9Tmqe30jR
kCtSy16w5ZU5HMf8TCs8PuugvMMo7TFaahK08XSGOL8Q6dGU1uv6sY3T0898jWj2
PzGWPW30xz9L+R1mnWA0jz5xOXHpX0KRWPMrt2mGnIQ1yPtqzU1Ndog0Zz9rS/K4
mNuvH01NYxBtxdLsvpUl5tUqoOO2wEWNKlVtJCuvPS2EcYltFwnvkeKGDyOxDhbG
uVflMhkDZphYDdcPM1K08UkjbKBr8BItC9Paxae5M9GK+sJJUjPlbuRLemuIOIhf
7u6GWykzkyFDp8B/qCcSGA0My6I0AgiXu2x0VVnIsbBWPrR9iqgcFvSN+C/YAtE+
pYb8lKK9vmTfufEAMd81X2ANMO9mUkCxUzfbrO+fhpv1hprtvqe3m014U+5tNxKz
N2Vy9rL6zCCW3kZkUv3TYs7679W6inPIA5bLSnFAMbk9Bxch6UIX1Uv++0Zocz32
KMwovCjGqxcwpfeWj+fMUZFHq5NSTJNRZW/n5Cz/8S892pd1wOH6t2sqR0GeFxxa
D3x6RGn2J4bR8Po5SDzvJKfZ0ofTWY2lSKKLj2EKUqolpQ/oRD1kUdTbWCPTNWaX
ByUhfb2FAVQ7+hTY0NtYzKnlNZzSpApRZ6hwicvbj8NICPc9jCMgQXGyad+A72pL
j7VJ/eUapMHDFNdxCAOAwObPwzhOPSExtoCO50WPa0m6rn+6TNwsZHR944sX0T/+
hczn27VB+6tJgmzjokCKppV9o+MTWnwPqi51+M/A8/imzgTqIpJNOXclqLRlNAe1
NzulbHOb55JySIujQ9SQnqEduJVFh4tizakQlEe2D/3ApM3wYz6W+hQWD3ZlBOXP
SSxgMxS5w3ha6IT5uyoAjJ+I0LLRO3Zp+4HCQZto8/b9KxM5lFlKwqRWfWQkgbih
Apev0S2+IatiwURfKGmgdjJKvoELMldbyQUuMGgEuCGF7fh1Nnr371Ie9j1adZih
jbOcNzVb43U9t8unv5N3xHnBCXwnFiKgWXOJXkn9Kr5a+03ykTG2oKoewsBtnFpy
8NSmAqRG5lGKppT6DyTO4dZa2o+focTWjQMDR+FzVOfvmDcdP4W1wpVa5bT0WViv
tAODO2tNI6+ebBuEaphEViI0HEXbMCp19v392Oe5uggR+fAMq4dVHltFb9IxouvL
+9P/7NzOVSVO+Do5M2et8hG91wG+1+TG7qUKxlJwl21Xv4KKARuDjmfABfnbWts+
D3HU5fYkeiR9ZRjBdCbidrUsiGh2o1a329jPwTAeQ4gU02nNcXd+klDpiqaA1pO8
vH++eqYm99gpc0Fzf/Sf5+FlM9rJRa01QsV3M2vs73JqFwiNkVc6MUjMyR0JtNXo
v8szoQqEZHNY5iWq3KXzvdef4Q4fCTpiRBZPEDHQvEQ3XV5Bj8cgaA4xTusd1AX4
K/GinCkMg0gMtNIpSA5XTh5obfZTN5unUepww7hqxfosghfPpvKxwa5lWDsD+/EU
OCNLKcsfUJ0mKiCl7+kzxv2OTYdA47VezyR6/o7yJgvTXVEgYzyavdbdinCW7l2s
RGxDIPJ0k1j6Bf9yZTIUv/YdLopemcrReh04AwrOKLAa8BymsE+XQtOjXXh+ECk4
sswlJ6PIwTGPi156CXTz7MLX7fi74BhWxDmRk4+6BUS1FxBS5kHE+ASdbftRJCBi
I+w3DdLL7S1sjs1+JcSLumpq40RKE27tdPtEhKivX1U1LnIXmSwcJjTXBAcUQg27
jSlDH7EeqPcxWO37UJXa8FBgW+w5NswcAayCKNyOaJ7y6OUy3D0KLiRmEZfwFCkd
w4Z+fr9dmBHDz/GEhuBHs5x0393HOeEGHk430iGHGBFZh2vwxP1jijpxKWBFFxWK
y6ZNaXpf/aHgR1lJMFmQsfBeHrgMoxpfZD0aatTNHMc2fOqDdtu2W2MZqoNEWrgY
0Fa9T+0OxQk+NxhT8Nz4oCJKfiMML6/p5ookfXWLPkR0tbYrT3gODhF5+ynky5Bj
zdzW6MwJDgbW2ubNMJaiFC6qQhho85aBvZ+BhyOxNZNs/VdGQUMd6WdDx6OYmcP4
7oF9CFqz30m0gJSqJNOAQGPD2JPOKnWHNyUMfjHmLCmi4TUMmIS7mZvbszwFfK9d
M9rx+qAHDwi4dSN+BoRMAVPkFdLutoolx7rR3yVowmkc4XIi3hwzmlPWjhBJV4/k
Lb+kuJfImznqppqGCz5zlg49CQGSKw6EYp2eRNss8Eb68oEGKpHVEqiYJHEZ3QxF
1sizGH0umA6sw9qXf7DSqr0eJ+Pnjd4JjPkZjHdAA96V8RPaTQWH5icVU4NCtYFZ
l0i4pwzr0EJ0agW2BLmBcQ0pVc7CICDtS2tcWNaUxL4YudPgG4YT/qzveBwQnqAS
GwFsjblvXdWsQ3GA/4Cse1kWg2uQe6Cwlid45VFjPz5/ptYE0PRJt3UcjBGBrINU
23D52Una16USKANuan3DUHfMhtoUBDXHOmC3yt4lMEUeqhhueyVu9dXpeBXKEjxa
y+YWCojNjOYOE/0oUmVgeBLgKkDRAeFqGTVSf8pV1cbD4+KfMWn7nFqtUAioeXHm
YdHQEzCUqwTvHDWbMI+dgTT/8Niazsw2JhDKa1P/OT7lVrtaORiaR7asauDPcjNb
ZzvBsdfEaoTWiFgjjUkKUN+W4reR5UlfZp+B3G4/OdhXx6GR1C6nBsb/olY7j8ry
xO5dJMgVpVZ30LebEPjNPBr3psfL33DyHEcWfo5INF6r4aG8FUPUeQSkPPuWHq2o
v3cfibDyGMMk3PUGMgkLFr3BbZVoNPHLAflE4e+MIEL+RlmtBvBGHaOcXNY6Dc/o
TCGwQUtwOTvgATGjDL/6iKiONagAEkhbwfgGV8Q3g3+5YISFa24MBw2dxklhuBSL
8xrpUt7ZyncgwM9S9zBGf156pyeg4BWmKQp4oESswmAJ6lDKsdVETCgSrhRMpvTb
Ss3kRH8aDBgv7Imd2xONUOtqYXegOF12eAuXZyinwij3GXRcFWpYa6r7YS7OsF0G
5lmSfMbcmwVFRmnBmJkbe+eF+Xx6Y+KHs6c3l6E28TxlZMkz8qVrgE1B8/pFYLAC
4X9AVylZRgRJL3gRUN+3p8T6/a+8cygZgbT7b401M4Mag3c1+9ohpFGyuQKu4+D+
sBO8NmDl/44MwyL6BKi5CyHES9DBASnp8svgh94eXHa18/rukjNW0KYzRiW3l5Vt
mwMY39YFxdG5iBE2C93m6lTstRyaG9tp0FfSf93EwmyaT80txR5inM+LTntX7FTU
dSzEtoMFn0j7DqD7c3kkm+Itahs8kMVssNGNtcU48GrBMHYg/txuHQId+6GOLid+
zsYowMHyw09xPY28gO+wU/+rpzUJWlOaqj0EjAHAv8oQ7cEG4207p4N6NwSwylJX
XzxnGBSQOp8CTovUVO3ebYn7s47r27gLhOmre7VNDA06E1hHHhGsiJRQRKUGh30r
7m8uEK/pJ3+RhPeiZKKc0iDVBNPgmRcL1+CKtBIJwlhysSBgs6Yfyo+5XjbNGQ4w
hq11G7ElJx//jx810bUrg3lo0yuss7pAq1SVzBQdk2eUiC95bHw8pcysXOzwc5sB
zOI7xrADZTDcCRktVSDS2S6K4ixKawhofNEFuHZBZ9I7e+kBZplAqhweQZlA0Mq5
hYwTgKfSenRx1t1gCo+xZb6CGVVydrPkxWTBzingyN24HNXwY0JpO+O6JOYeBo+A
RddEpuh7Gv3uZJdRBmJge4PDHlRkJ7fEbXVqxPMNl6Wtl/7JVOyzlMr4urCiNFkE
9kHcoeHL2kRjgeQo7jNDyLSRuPFJ3LSzAVkN4FPDO1Bfewzj0lTjFTx6VL9Ob68i
jkLSb+ukM1KyGr85sHVurSJ4GXPF3Kw/VqOqY7nrsq3bZptr77/2V3wPHRTy6MnS
2yNcYgTDy58DZkJQi0Q/9hA3ZgP/Lvu0RFWRTiOrZkVh5h55VlS3SA41coLNv7lu
c/5ZHOn90MG3DCTu0RsAL1+62c4R8gP47su3FitNUHzbFwFW3P9iHcm+tXXd8gIR
/EPYayhOgK+i3xgcq5CymqR2/CAqCth4pEd5oCs6BEHQabRtRCA2LZeunUmK6rj3
EMtJdQvly3CiDtLzjHlJXC2pSvIqcFl4t7/CQd6yVm7yipcBbWK3fTA6DVJkLp7R
gBa+ptSDRCY8ZQibajVcyPjCMo3SsahBlx1zWeDip0B6B3Fhne0E5IjIVPQwZHhr
olmr9Pg9S2PewuuccnXDTy2pcsOPLT6gotYpvnwDb1hRUTw9QH6uBD2Ek5qs7dwj
L40lQf18u878RfQ2LRWl/chDHrA33+pkmH8yP5GWQBXlIBa3y8Lw6PCWWiYD9mP5
kk1vPOxdw5YJV/E4XDZ2o+RbNNdG1TBgwX0qb5IxZUcujBqD4JhFbWTN0yvImR6k
58v0Nb0eQXB/W7JEpmN/ln6I9stK98UIeWHD54/ZJNyvwSDp1JfUzk2r/US78PK2
n4ADjS3ArL+INi8izMQ7qjMSwemt9B/907l9zmCAZ8iXy6L97cj1/nNBHjVPSo+1
0mId9pVUQ6uQMAEzaLAmnKpTYKP2e24VirwmCrQKQ5ZPbOUjp6e6ErMo8LFZi264
GvxbCIQ/SrMkAejcDK93njNOjfjAnmeF1BzyAmXZAE6Y8nmcH/kwOI+M2ONFSvbE
iHnGdxZwi+wgY3vJNppB/AwwDsdl2U0LuF6/bupCMYUNuNF8KRUqimMmFN2Z6Jzd
DE8xgynskcW6jKvrQ2DQAakdQZHvfFO4sFRVP6yHAPw4TOz+XaYUkbRQUPHPks2r
XM+0EIP41MisQTYcyEn2xqvl4erGadrlGW3exI5ynvPgiv/ZOQ5n/qJCzr4CGGwC
bkYDPV+6qPshnt1xw7qZ36zjTIUAcCsQLHi4Yv5Jbks/UrjmxIgffLIhFhEwFaHS
AxKgZP9jWt5tcUsuWLaqW7V+IEPsXe5DABCgqLphODx5KzAPKcYru440BmQj8+U3
CRXt4TFAMjcFt7CinVdBw46fXa9Ca8vBJKTN4hRj0AU3+6sZ0z/0uget+KRvT3nn
umVmOm/9ca2P3Qstnf8cd9qF1SFyZlExrAg7sJMql8hgacxDw0d6+2J8E5/Jx4/e
Ad4V5ySB8RTSsMdAI2t7POwGMuVAQdvnp9r4yTNu4juplGs1Q9ZX0s4KXor05Y4i
5yFoUCLWh5R+4BBK9kJkwbrfRNu7x0HcONhM/m7v3qCgic/MyYq7UkhTGQBwUBtH
K02ohD8gG5+L3Ob8qwYR+v51mhY0gzKs4q49bCF+jlbapgFPhdhB24foZOxRCHKB
nHd3pCVvxjJM6s/nTrbcZOj0ecrwuvRtwz0DX5OELVODRmrjeeaJfJA8t0/uGhNV
F7Yr//eewDeom5876V2SeoBcN2sx9zbYUi+5dPXlVIQPlVehB/7mglchcUJCfyAU
eu/DqOUSCIvX6FG0L/c4JXVzZjeUkcmF+Qdejq34T8SfGfOwu0eGpIyVa+pe2Q0Q
M8pcnuz0UsGwSzeVV7Q6JLfFWUj/p/3InwTU4LmxLTYgOvs1khrUM5uI6n469i3a
21dvPqQpUR/5CLicNZFonJoejRODQ3jIvayGX4DwC/qqOr0eut7bCIKqleNrbTpe
IXidIKnIzcLiNrL+K10KbWsLbopyDjt6Vt46t0g+f0y9EWnnCmHUUYrq1Z3aXrgZ
juQAspyNYzlKIaqXYfPcszquUHmxXGzeQpmYYoO02LYUgQHOvfcdLSEDWT0bSiYr
t0Jrw2zG9E2KyMDT2gXYwN6Gugfx86DhkL+IJkcfzfWkj8KiH8JOhoib5zl6v1LQ
BeWqlb6p2R0sGpjOmkmZXlePCXUalbJFqnd2mU2crx0Dwj2yX0nkM9/0IdiufBJk
lZ7/TO59hdarQGWKlEYuVf4y97pUXrMUhssRB5BzoR8uAmyaYtih72vbB3NfRMYi
nWJafF1zUGF8E1cgkLeyRpDalLLXXorxGqIKo/o8dwlIwuXm1IgxhdAc5KAi+C5G
8b4a3VfvIVD9HCC17WvV34f+T4I+aHLry2Zu35EZsnLi6hV8jECZWglAw8AuL3Y9
7F2KadvsWRSf4PV+CY40jQvEXsDkl/45GeDeX0yjGeg+oJWU9YxMOXtIp8/LSoo1
ldP+D1195nEMh/aTIucqHpdex1qA160S6blL0P9o9SUDX2Lx28GbvXd6OqFS0hE9
YVt4i63iSWyv981nd3Ld2mXGvU2RqDfplIZdMiKxNVeMvkpRyhOI8RHO1QL5RZiK
rhdvCBXAEklPHAGpBud9kp+sBgM473aaeCDdMo30ZgUTTfPfVUqOapbuDURvLiSy
29CSo6naXheM6PYJU7zq2CKYVibT6yo8o2m3PbReg6gSMjI5DpXCDFBhcjEPT84V
vs+9CaebTy+XYjTLdXnJB+CnTXw0NgXrbnnzWboXAY6fxOdFOgoc+MSMFwbpM9a6
FxjavkxiqKdyRWN/PLslIRkwrdX2nigZzD+Cxk94gP3JJ78d4Rbw+L3yll+FIX9C
1HHbIArBe5+33aT1c5L+QV6R8Lx9AGGMxX4Nvwf2F++alb3go3iU2ldfMzo8LfRg
motNm8fSP4WFKJMQYSZhlIe4CzGcJ/HVVigfMtoC/Fe/bKvnu2i1uLgw8KficVY7
lY/9S/tSWXIBpCWilPfU19cw+9mfw1V3coJD064Id9w7xLeJtycTscEgU+vZLDF5
1mIZw2KdZU8XbXuLid9XAjpgEGtwRtBrQmkVFSTk2M9fgxE+NLP1+8Od6XpRRTkh
KBweseWvE0djeuCpaMlC8ZYfBNT6Y4y8QBIWuX7ydS9O93MhyX7jTE36mX2/x9VA
To0LzGquRNLeFv8mdQH1u0ej0T70ouIaaWGfCcp1K8I17uT3ybXvTb7hJ/lISzXc
UUIZ8pO8DGce1N142cxddpfGa9odHd8oo39eUgSanCjGKQKQA7ngg05d6PUBOOSI
I+A6J0Kr2Lwq3D7X23UGqhs04IC6B3dzbmkbuVsHgyLwBzyj6MCeNjPGLwNU3Uvg
yDvHQjFcr3FlXu+gid7IPSsF+kYLMllah1mNa3FYLkwEldzjPwyjezrbCcz1mmf+
ER3KFxCZpXraQR/R2DuVWhucDcZOchgPC5Woxr1xRbPwDupvtKwkI9Lm2ENX9Qms
AEj0arajxVt/bgPgjY+NkSjMIwrsfudlbFa40mzRfTfcEY2X3Qd9pPLdSvdyly4g
k5vNXDWmO/0OJS7Q6rf9PRx+wb/6C+RQL+wddDmYvyQlbqNf4AZVTFtoyRPv3sxC
yZJZ6BqMEZySojwjIU56knzz5h9QD53IbgOohArv1n/EfO+whhAXKs9HdYuRL7fm
VRwFMoeJaPmvKbkFS81MlFz2x65SFHLZIOK4+O3e6wlg0cPGyEgEd8pPAnPsSWva
m4x5tBh3Op3IWsEThA6a1MKRAgWoO+x+nXQT6EM8i7w69N3WWvfWDXGEMfm1ycNU
n3vWS/i/2Lz0G6mXJZMcRPp2w6G+9mxfYy3asMW5bLaGBSVSkw75SspH2aeAFXD2
+sr98J1nJNMDSm95EdUYPrkDAd+phc7NF4vluyPZhxhRdSdPBNDym6sIP+5/t530
tI5KHwpfXq1pEovXbsgJwW0ufQoTIV2jItk8ebd40EBGNjpILufTn1s4hb/V4W9V
odloUWU+fOgvIELXACnTwFsAv8pjphVklAiksXklKgfcNzpKJcGWGl11r4YRlgTX
9vf1ydxQ2j+hbAaV8eOqc1vtMIr6MKqUtRx3S02Erk+iA1Sri47esHGV0T84Zb1Y
AH6BPpMJ4GklH0nHJY8cARri0VFL1Y0Tpu1bpEWW9ZKph3p7SOhAewgJZwfDAhKX
kbNKQXI9HcrVWvdKDb7/1k7DTMuI353pOw9hhbpi0MXWUBDaQk1+RQ6+1oA3PJzJ
VxrVJUvywCszXT/Fb+DF71JMwkJ73ZwsjYqJf4yPS6wUI7lVw16MtQpeXG2NGofo
ckuxPLIYkgmM48q91BsZcwsO2Yv8Hs9OZP/GQ8xYklWCUkaa/FCXibGmkEumpuVG
WcqhytPhSrXk5m/nSyjxhSpZPzBx9z3VYW9aR7JHHKP5utAWxqqsxELM0jP8w2fj
Wjw3SbikoG+fjO+oZwe0+O5zpAGOXklXVYG6QLv9aVHAsROQCePRe2X/zCJLOTLK
ZK2QMil3r6Bmd56fwSGhs84VlBgDH0iypWOTTCSYXS0kPqyOVrRCMcaPLrla2b47
Nef9yhF61zixUaDvCpBJ3a3VF6VtnDQ3cHZqLwI8SQaJYJ+CxLfB0rpdSTtoVIoV
vlkzRkGiUm1WNb14jYK6cb8ZJa0R+ja8XlWlqhcK4NyMAxHSeCo3b9hXrhk4aFYG
qej1zvXJjizQIFtQqkV+aOu9mzW97JOLqlDwZwD3wqdDvHplv4VagmvNFrvqu19Q
NxQBYK0WpIBEshNOlT+kBcHM8beeVjHbYzzY8cPxzrwUJAmW2p5O+51AfptaRSon
OTIivIAGKlLyHFGBlyQIFcLjGJ6aGn5p8rf2wsIQo6Q+Ax+VXrlsDcbmJ016s8vc
64ADsNdu91ribt9LrADgW332VqyJe+NoX1vTxt2DfGmSujK9pXH1vt8nkDNxnTog
Ro/bUTCdsIPtSYdkc14VncVeqvgxLHhVNFcuqjma4+Oo7biBu7lodwV4TKLP4May
Jbx9iNojRXeKEHeToc1PJsgphQCgq8dcWDOrV+39T5CLZG2T1bjYwg8dFsyW5YD9
Eb0VXeoeY2rRR6mYA+JXcjcN+zbSx4NyXjXTJFXVLFSOb8LlMd7ggDaSJylSIO1n
1/wAR2c6suN8Ybmn1XFHhCIckUQ9IvgHEZ9ikiBy0tefTFHXq7ZXrDnABeoccqdV
VB07IO6to5obIXkDh6jP5aHDq/3HbDAGqZd99HvP21QhGYNgNG8Pw9Pxe8Sf3eS3
oX/+vmhEqccRNxZMANbR3cTJ4cYwdt8nAPQ1+0XUDrtrU7O/JpnQwCjhtQQKDUK7
wbf3G8mAjjMdcY3U9iNKq9oDxP1OcTuhJZTPbB4BIQ9OSBtvzQfg3MZUB9CE/Id8
j02FD3JkcGcG1xKpxwGd9e2PAN4EeLa1uiCYGbbnUioHN/D/fxWdyCp69MQXSS4F
TosdarxJlWK5jRzdorqxWdVgl9D6+/VhzD6uvr78Lz4TuyTFmcvnpAIqddgCcZJ5
2/YkKTZIbDcG/OzxWu72guFBrPFdYE+3wtAk1Br8ATP4lbU2l7wyUioIU+XaguKc
v+TKLoIfhOKY8+7ihKh+2c0rtxt5q7rvOBXXAMrANN0hjtWgt1zhEuHncZ9oruZT
ujSGuSa3CvvtR4j8qcCfAJFYWcdPQMHV803VqVabpG2hZxyiseQzln1aG38trQ9l
SJj2Hw9sXK9Ofxxxt4FJHVAEsHkzpC/iVbXr29EH+hujZfoEQBqoZJ7ursM06+v6
aULc8x7C7ZqvG2FIZrvJcq+qydqdaPIRfkZJloyC29l9YOg2JnLZwU8uhed40w/N
Erzgnc6a7K5HotDvYJk90EetEM0fViLzHccNvtUnYrU6rK68Tg4u5FjqvbD58Vxy
MxN65I7culgsRwvXw9a8T533BQHSNdxvLxaFkIX+jHOMKBGVty7esQIQXYTmS8ol
zDHbFz5FpQlbePL9BUDFpF87ZvUpH/EQio5A42Bt4+rpabjN1QGDHRJFSgYFQ5lo
+3xGUIfeQ8RtADqXRXtmu4a896ckrnvTSiXIoX/N/IVNs4H6FvvpamNJ+FuNLzwz
oq0vwfGgXsRCM4CEwxkXDEwIiKzalA9vhgKed5F2OyXEBj2fIKSYMdHd/1V/BAhd
njTyxQb4S6IMqCEN2HG0PAjx7aHhnYPGv6qRBrOgAejL+qNnGRcZekTMBlYI8DZ0
1llM3DKzNRFTCx/tARNTygmrbUJJ2900gBWu8GqmsFJz82n5eX7LjrAD9JLix0Y0
tF+2C7kfPOnwS1P9q/wJ1jeLOslt7NY/pUsagvQx7TW5/XLgiCKTXvpdQg4WRfIC
fgE5lI+WUrIMrNODfGZPPCiyZeZPZBqDtJ/PzK8yPbZKVzV3N+BjpvU4v1NLuZsT
wS8PNoeZUP58bZxOkyaj64COhftnWI0KZbPI10CflmaD2LnbwMJc2XwVaYzgzFCW
7kV4icBtKbiCAdxdAUrgK/ThN5X6t/2FvehqUWFMr4ESxmgWwIteZEaZeCK1GalR
BNPUPzSNLBhvM/DXgjd3BI+okGnnxLgjhPq8falyiGLG/eB2CRy84YGlnP4YJ1Tp
Nz+VI7eU0r/cIWRtFKGzmC2n7AKmpUms0AslTl7kNA5VRsI0qt/ibrhPhzIAMhTQ
8u4vVLcssloflrwSa5wmsDiH9uimDjHypFaOpI4+1HpQJhvgSCuN5nIxq8+qVOYM
E2lw0i9lizBFahPbVoIvxLO3sq2J0sLxgmZgXmpj9qZYB8pbtd2k750zQ0y8Frd0
K2NCB11ddcWEl+WOOhU9HVC3a8+IG57ringngXB88LEJkSdSfpF49FFwWZv4RVBq
ytYMJFJLEZWQaaWzOH8CTi8FUNhUA6iDu8Qr14z+5tGOclDfZW72oXF7eWBjbBdO
ikfTIXaaLMbM279pZ9PH4jf8E6YfYRpJlUSniYF1gLhb8PXjvXClkf79dZI4nVin
7pcTW3gK/JO6IHp+MNv6Y+BNpg/Dy4PZW5eebGuM/ZL1pgzbXmQDZLAxcsfBpYfN
aAwStwS5vbrOiRZHmcJUIHPwICJ3t00tQmBcIc0ffCRSK3p0UcUiV+MXu2K/WgUJ
rc8S7owO1/u2ktdlq2Ph22nYyyqXCnEC9BSmxrRfpuk6C+zWAhUyxk647XE/Os/M
A1pl8gQSmORYGGGV0eZeDLZL9vZsuKPmfrMffdg0v5xdzg2D4kVrCWjJwgfkxp2x
2I+ZfSEfh2n/LAhzN3gHxEfhV8/25LTAn4tFkIw5v4Q67ur/5/xFC9pBK13MpjXr
cV/DmCOULSeJ3qJkiipesMTXCD4do1khOpIVD7JhnKQe3nk9Y25qfjc7Vu7RF5z0
bZoW5f0ZQvaEq400KP+QbXs6BznV9C/p7lTlDLF15FZLf695F0znTWQNc7hpkdTL
Ssz28nueiJWCY8jovPXBmr4bTizyaep7gHcB9vX1ecX87nVmXcPYpkDNztrLQUk0
NMROIneNUIbqjTQC/02kLlUELgAG2oAsRBrPPCed4TEkrFA4rHSNrgNdOX2kDL8B
KUkx7ID5BQ02VCM+3TH0P06sPAfoN1m85g/a30SftkbLh/dP4+N44JymhcI7dGaa
bTYUaTv6xD/HCJMEmUtUr5XsowppFKOfSIzLrymfxMwreFJWLc+DYZ0cSK70iW3l
HhiDdqadhaoMptPXRj/+31KZp6G59Ab73MVrMZVVFn6fiHVu31TKwGBWyCTvHg6O
zHCv9rChjpVxGkIVKRLKjVAvXEWxstWq05k1yqHzMQJChd9zuflGA72zc5UTumu9
NPXr2hCleTOC0buXAsHeImWB9gC4ChVfG0xgw2v4fxeszfua1BXSiIEnNsmkIrzD
WzrDSus2Z1YKZVPLrpxIg2hn7YFRJGogm84yAOGIh3fmHKCHPrRlM8VYDr7SnH0o
J45fA57tS8YwCWMxyEWayeta5Yi8hi14Sf2u6c3ZhDysVHFAUSk+Ltm3sMf2q7QK
8HXauSUUKfij/cM/K40F4EsVe2YlRT/U8vQhCQRZFmMtyNBUIrHhdujRg8TZwOEZ
q6s7UxE2fkZGht0wsW7hHMZ3IiokJoDEkzVuajagpkljTBhflxUXT+rziN97LlR+
KgphzxUvGpw9Mc+pUqBddTlvAoT1mC0D+NDhTigEQLkzBH+PzwPXt+pICahcTqlx
9c6W0+mLlauGi6YxzEW/FUEpOE6kbTPtIPQWG/8OEHUqKxD6BCbHnVCAncxcIQr+
0EXAnaT7vhjFvvAvzG+c1OGnBKrbv50ZQ4+kzs4GK2F+Y+Fc1akSOQ0SER3KZB/E
03IQL+BAK1bdjWaM2mP7md0AgXNZ0ktapH7fOSdWCbS6le8qfhUSNcnMD9qSv6fa
YQxNsahrkeOBk+dgeMS5dkK4blT20jp3brG6KygdFZ7jzUR5q/6Z3amSE8jMkfwK
P3R3J1QQnwNPCKSIXyKbgnsd8asQGZaV9JNWRJ1TjGuxQIfzUZihKi2DnY2HJyCK
u2IzAaChvzrbeoK7bobKC6EX9stXaVorV+y5KcDVVrcVIcBNbJoOt8ndCc3IKDPj
QJr0rWZ0YNtoYl8GZvEc0puEExkzbqrk61tD4kppS4eltJWxkkbjg2ky4NryaBG7
AlYLKRDRKM0ivlXOsxxXXuriUnCUemjscZkdpAeMBx/4zrnNDcaHCJBkSgMpy9CB
iIfnybRLXRJSQZTCMtIg27Gy4n2B0LZ2Pc76mvPpP2yUd7MwPoErjC0KFRDVPqgz
b7FkkS+7fmLbBsKjRo3Rx4hDfKVzD7Z19p6QT98sKQ+i6MMYXLXNtmYNAVreLere
xS+5IhEOicCPosN9cpeabEamL/bDfbpcOrgHdG//ftRWwXwhNTJuS6+/FA/gDrYJ
BZsq4bEawsM1qvZT/GdCS6p2ZzGDmQb4W0YsKkRFEkjIEaockudkrGXfZgz8CKo+
wndd2V6xBdAYx9PBNVyycihjQJzDbcMHkNIQzcYaH+UUqDLxuk3x1RYMgpHi0D8/
2GYifZbgEXmadUslBBM0JIO4SaZB1v7VFfDio1xYxKhABLKPIMfgHqih5YBb5HZe
jcWQTrR7URhUIhzXt81gJ65xIJoZ1ri9Ao8PjIybp5/iVZ58KsYSHWgnDF4VVlGm
dQUhJf5k6YiuC7Uwxuakna2ZCdVAHKVHWIZ97tnkngp4OFlkgk4b4Tzmj9nbgBX7
V8b0zZc6oplBGpklrzOU3yUwkrSLceeBFcqJ0+XJIs2zP5nyZ0GQsnj00b7I69U2
lW57QLxvlo7gnafuqo9uuWkgblleNkVQGeegXVPQL6Zg5eKdcWdE5PrdVGzK1uaW
hTfEfAvN9a4mXSHCwdx62Uq2385CBdAlkUYdWbnqNTFjSwBOcPSyPsLkGAGHLHWR
jz0sXPRVEz6NKW2JFWh2wHdlAryr4zfRY2mRPeCkF7w4/z1XwvECK6qv7Lhskxlk
T6xLmO7sTlshO3FwLGqnU4VPs70oPXH2J4B0guKNxojEj6ccVyDAAKhLeMvoorF2
Z/1B6hhyCx5Dq5MNybMLhSsVKVjsMGDmFjRipAxEkbSXg2KeWyDCu0LPP6y+V3id
KhRT+QEUkF7+j7vOgoRSUmE61J57kaJDvQF54d911eG3IKyMdbDQ1MuavnsEDpY3
KPWAG4rUwmGIjIFFb/LwG12FcCOCPN7W1nJvUU4fH89tQkphM/1r/wQNPYFoOqD1
+ajx7YXEa3CtQ+e83WhjxL13SSGKV8gif+9Avdn8g5kNNBsLSQK+ibp+F/I9bs32
MShQCoYcnW9XMalYZlkIA/Jt6JIc1V8rQoM5Dxx1MtMhxpHenJXpVcmI3mgu0rhR
3gQ6K4vBBaWHqLroIcOt5OvDK3CVXSlUAii+QRetpVW6M73k3aB3rDhAc223aCab
5V9WC3fOP4Os22JYtsRSembG3P9A/jPtembmTxIHH+H7SRaKIgagKb3eriEEA7Xk
NEFCJPhtBrZAlnRzf5MBRep6cMapMnUYsowZPtJJu+S3AAMuZwx7c8iltebkuANG
cGV/LaxMZb5r708Eu7fxwrfEiQf4CFWGxJdqyWoOe0jjNexnlx3LTOfVpr+WuhNT
Q3N+bU+IA5lu9OUUKwcXkFLBcLs/WQllCvnYZU55J76TGoHAWLpIptnRWnDQovrT
GDm4+29JFMPr0YDags1tofUAZUG9J3U+hvprf8vg3ZX8MwYkHGUIVFSLplWmfcyk
Xbu9qqAk72vhpTow6SXoCMCM37i/tr4u2kknF41RgdTLUCIrvsQH4zxGSBLSL3Gt
wv3+bqiYTkF/Md+LH3OZyGphPLAvSCe6892Xx71+0PwUODIo1RlL0KICrZAqujzL
lXhqH8rezqEY2kndwkGKsuDDFZYsITM96HhJo870JaUmOKZ5i6yt/967Y//QmWtY
9BjFbTPvq2+R1CeQ7BVDVmhLHlAqXU8EfXkTj28XD+tZO83/ObVZ7v9H2kgJMvsr
NX9F2oM8uCqcK+bHu8Pms2oCfeB4m0HYFK8QMzFmiRUHjHWgLzP3leLj85FDKWUp
YhLbrJGqsXXTb2k+H8c3b4cm+t3z64ji6uwRI69otoMmRog6H5CKtDLVldRTbQiN
7W0Mo/LfI+cEBtn3QJ352uCVxZzqJxoAA5K+jaKdCsxmiHib7x9VDTIsBB1kHKb7
oBdq+b7v+LP3jDzPuQ58LLMCju1BFuF1AwSOvqNjfSPJULalBhlo+InqeQHaaxqx
n1y0vNIfpflf2UCCqI4pVRIqnlpj5rhONNm24+pUuUwe0f2xTEvjoHqx6g4GpoUL
6XEkoxouQdkNHKPPiyOi2cm4qSI3wKkugK0Gg3CoWf/w4l8ZswEZT3vBG+Ks+avH
98tK/qGJLe/VNRf/LrgQRos/pCdIsoRdV4nJE0X/4I0gvdLeP/9B9IdWjHUNWWgI
eHOBemZ+uWTUGax3J7K8NRDFbEdLHqvPoKZdyt/YNqn/lb9KjAH9mHwrLxGxF83D
GGHfAVX27gpt1s5E1I1qEUUJKdg7pGK9wEDIMiZa1YMghPhLqWdBTX4d5INH4Meq
cwxq/iHSWLNr0NfxLixsjU70icJHgSXggc1WwK8Nt+bUIWRVFwxydYYPvIKv2/7J
wqyxUpJywKCasXgUoOMkTFr/l+0bkYDec1e/th3gGQeQbt6NwNqi8wqFA4xs950E
E1W3ZPNMQDDUaXdzgfcdtHjj+a8XAkjOL1XS3hhUVqJQqNiT79P8tB3HbxvX6SYm
xENaHYQVMnLQjH9+UZPeOPvWH1TPT/2EyeAFhibwo3Jwu4wbIibIJNWxreWe6Duj
5QKa/pd8F4hzmf4QJ8H8fRV0BbSVek6BWOAzopTMnR3O8o/YfoXaXVunwayryh9j
4qRXLVD5BtMr5QM5+HAVe2Roq+7vy3J81wHHIpiU7WQjmY1Fy+kqJgWOPj0ewfsd
V7aalQY4U04RBJtvDJ5fKqrJ4prhCCTphJ43an7dF+r+41IH37U4YpLOplOyuQm3
vadQg3Q5K85kymEPmmNdw4fZXwmGGGIbuda6QEoArlRMrYmTWgYn5k0EnxxoDP7D
YPF55cqaVstDGJ/BQ9Lzfq7BuiALygL0tuG0VJpv5/xhYlsHQptpMyl3OZSRLxn9
Q2SCbM3qAyZbfi94z+LsN+zNoH3eCps00/AARfX69A6Xg0P3+AvrqSq42+cOdoq8
L8xXezwKme+JMve2f2bJM0su+ru8eID3m6DVXsjdpX10LMlzC4//0s6qrJIPgwPY
M8UHNMR7A7BKBSrcxkRVnt/1j9Mz0UVKHyDxwBlSsdoy34oDx2u11yDCHllzzo8b
Kcsdfcx4X1V6cNtE7C//hva5Tz4w9QS0YTfDF9T7SsTldFjUpztV0w/jZU3YsZrT
GHOcTj0tdlBv+VHiDAJT7C83LwgDz2/0HgUbpziX/bd/KIHtgmlYXl5BgC3+/a7N
86R7AgdyFoc6ZSLvxBbXI8ryuZNVdcD1H1H1Hz6FH+PG7kzgbDvdaRCG+E5PT5yG
G5L71vvSugjVavKBj3Ir2ERwIuu+qLhOi87oXBjrQfjFcNwFOOaaKQmxBUcOGfbc
OGfyHKBMFkLhmde6ojHEgdOgsfrM0WT85rCGB7YyjIr+hyZtoiamc+TFrpqvGc/X
yrk60W2fIHznk6SgmgnEa7zxOs68xLGhzN7hDoKan8VhDLfeVuCEptlsbkG3/6YF
6AGciepHpUDodulMqsaYKxgkO+iV8NI4n7ieZ7uFepW5N3rxzADuByg2OYQD8bUj
tkLlHmnP/jonXExya+0/exxYLe3Ttct+RnMYGUko87joy8b+VHA9oT3vrczeqp1K
0MbY3HmBfnfGkTsXWf3OWGTngra5OtYOqaRIpTetsAV99RonabPqa8/ovo4BilRP
cgF9GmvJgzjmGtjdwWrR8w1+IzJec2H92fi51EyK7rloG1w67gD369yKmZQKNbbv
ovc3FYK0F8neH6qSryLFU5uPMUFHRj9wSR9N/GW+6CNllv09YBC1fkkNDCbxz3gQ
uCfGfbC7Ma4wuK2C+ZvRmAd4xcbWglz85LhxFPBdWYqMrVv54jEf2Zi63ksuWkgf
BdDJ1pppWCUaBxqbQSZT+7pKPxaaoKU9THmt8tky2MgaYNGDt/5jiomSHj7+w0Us
raA5HkkuUGlgR6tYIHdOyVL1XHxL5kaATjMDosHdLrviWpc6JR16/jxHjQa3m3VY
AVrWojvWujlQ5TIcSUNHcZarg341sdq3MHdhjxrCtFNLnALd+uS10rdoQkfMFpHd
SEmVyqZVp3afezM5wSSS/zJNjsrh21F4sPE5gWfBZBduXsy/0/LMu+J7Zl3OYCEs
Z8foSRwqoJIX6+qWVFPh2GbYDAaiBL/1gm16/dFnadl6lw94pTgfL3Oz95R763ej
YtqyURGYcGn7Ho17x7bu81m1/fyJqVQgHmuR5E6XuJEmfdFG/t9Ngd65VN1e7Bxx
FZ0DNd5GRul5dyk+JIWBlKr+ZFRZ6UAN9D/uA9WaL6PEmvF8LSRc+thFEy2+yO7f
upEj13h2TS/OLbUhR3cu/DQn3xeZHvo7mgL2uYF+JjicQ/mCVQLTGfB51j8WuapU
ft/qk7FQCzr1En5HNRscCaX9LIxJPPaKt3t8ec4U/vqcrHbr+iR53xWWnQi4Y6+E
BIjAqBEpEnUQ4kJPuXOP41msxdLpZJe11NekUkSP9EX9aFCkVJW8+gX3RqcjpjAi
EsslImUo7oEKDC3w2afIjHybgCL0tkI0k8XwW5U8UDVe86ZDPLo9IJd5EvxR/4Wo
TPwHB8v5UxkbpqN/ssYUV1LSLiEIUiq+rs91zHUK0yqZif2iKreoM6E30VoN3emR
ITtizb2ucfL6FPUN6iGH448wuQbCwHaP6eIcFOm107Hzc1i4L+yu02bKD4+joNW3
F62lgRd+hxKSDD0k2TP/hKSBQajFYXUM/MdWUPc0AdDgokA5a1zYSCcWyEfDoRnb
NpsAMBON2WkL/2NBVjCsft+uwqgkI2nU8zhmIUli7kk6B4NioRd0z0YveiOBvVzf
+K2kj5lgxppca+B/e0TZZXcOLqQ/U9DNyZhLQvIgz2+aKSHBPCdYrsFxd1hOPUu2
SRD9CEEFT/xnCUquLa2bK5nSOCQhCKwgPuxg5OS3YZfS/8/fXDMJiwahCZjq10dR
C0sdjK61Ec/K4TB1QT6D7dAiwTiulHg3zMP4ifGTaTZxKZ3FXsPRen38Cx1MCmrD
6mNPPhcrS3nFGSXvRgW2P8rE7htuEUzxUk/P0T6iuQUIcR0IUKfPDf/aW6IwtG5T
jmLlFfpLP0Z4J3iyY7h2904JTBTtov2mGc29AUPamiCvuelx+yQYdSnuchJS4SpF
E0CheVz2UuSdGUbiJDLM43Oj19EsvqoE5mQccCVQ7jUzIEYu6VpHf3V8LCcolVZ4
x1gRkvR3YHd2WhAkhrquzAtMNKPEa6eLkvEWZ6+yq78oBiWFb2JvXb4EFPiX+QYw
eV0HESUZQSdEAqsaitamO0wuKcHc9+PXvFN9JDS+Qlow/D9e+vPrCuKTvhbZ8qDy
FfaFtI08BguFApo794PT9DmQ0s+z259jEyrTA0vySY20yJ/n0oZxmzGEzMcB5ktf
GGC9/U62omoH53CtsjiQvA/2JcL90YwZrPmvVO+nI86eTynktEHe84xvU251Afko
BnYkaT/9Bth+JZ5Pb4sGSQKfrVfGuHq/wIf4clGOII+rGOmx5t63BtwRUAL6+XXm
xvVCIJtrl46vjjBXuJYYYwOww5i1fGdnOgXjtEmMUUwJuYjZYjOFyvpEQmXfvE6A
IxnlZvJwUrV/xScp9rX/7cJS1OO8dr7bQJssu4/PEBsb7rEdhJQFIFddPUdFXXXA
2KZeKwxQb8OErijHxQ0aKAoq7mY32ijFhFUq0dIf+gJl6ipDY13h4R6hKCQx1HFH
PogoSMuPRcjYGsPWWnbLjyaVGjjSifuLR9AaeJKWsgpZNZiFi2Mp02v8yzelz6Y1
DBG/Js+y041pTJ1hIs3zdQx73AZirEa00wQOM7WQ76kIaFk6UufGrBvhJtHYi08s
H6X14d1T8cUmYrv0pGeoD/n0p3zwqhdZjtcsQsHlYn2X0snxm88bDPTuyp8l4tQ5
VHXNVqyJOI0nX45kA1Jr8pv2DvBjy5HnQKTVg+dkc3Mt8guj02Dab2pQlpg2UWYx
sK11mV4fdvyYumXf5NT+ptjGSTCyl42/9wJ5AbxvKUiW6EWUo/uQkPCyp2vg4dcQ
EcSgZGQ1mn4y39ECPwJFqj2xRhIL2VaB8LwQaXSZt1vDXJtXCZfDue5FEfbEQM9L
7KjOVWXlWoVg/31Y0TD1RS4eCe+LFY4c70YI1zdQqn05bX2MTsKQ6xGmVckIRjPm
mGPXuX5MxrI5ar6iaRHWhSGiocHE8DDvDRlASB2YX0CambRSmKjq8QeeXjWfOBlK
PM1hgK3lYeaXkHG/c0FjqfVOlRkKfAlLCMVCoOwjcFKImeC0X1iH25xFJuuPMYHx
OO/WpoG1SQaEHGDL2j244i2qSWrONGczTUz+2z5zWERmSkMEOtcH+8RI2HR/qwZn
Ol5WxspmOAD+bnkXrsuSYyQExQRePOqD4uRiIExA3AT2pLZhUlZY7D38/tbAJDjH
R1aTsiI+ydJJRrL6Sj2h+Pcerm8WmHRKYmEfH1rbQcWMkwBI+eMMG07Vaw5+kR+U
+YQp7TCilDRpjrKsvuEbXEI5MmuAD2uBKtJAZWUP8CQa/9Reb0Let/vwzMXLf439
LTMsN5XfG4Gf7DXjNNRZNK3+TFXH2mN5+moMXSPeakspM1hhCO1UMqbSSwXIcC+q
t8ejFRphf18r//CahqID2XFlzHw45DK5X4A4Jnbbbxu2wsLx8eXZbnpmjEApbLOA
IQdsjyVnQbgsar8zpkmkXa5FNJjeoLQKktdUa7mmScNbTCoY74FwEsxUMkA7nSjm
DJv1dKZqZSDwvwSawDGnO88iu5vzYItrJzc6ZpiOMdxbBWK3QDzmaD6+GQ8h3AY2
RDOBL3acmkVd9IwxupXv0lg0Hy+7fM8rpG7gsTPt4VA+MZcjtOJ/ZjWcKkqsMMm5
cUtUzNjwvpaPPYcpYIIYhhT6C7Ng4re+vfRm28T71Pcl/j0JygYK8mhiP/azfhWW
zuAjRTcOzcy1NI4TmWgxr3uoeBX/q1sBc+fq10iV1znOY7brQqn43O/3VFC2+0Ba
0N8acbAPl8Iu+GlzH7TX7FuNNejLEgxSc6dt7LAxfzMTOx30E1epFgAeMeRa40Pa
2ZlKWzmZoYVF+scSKENwOSSZnjAJBv6F+6YhgC9RF2zxj/xdsJZqHHl+EPVwSGPM
369EieJPJbpC/Jdre8uO234fyehLdCF14e1nwgf/YcKYWUOAQI9TU7brREA6GRtF
gz9swiIA/pi08LD49FZAL3foGOJCQMSipknQwP3a4+4GWeDY5VIAuX7uZPDToj25
0sEuYpC4RzSb8GhJ2ezIJlTL7gWyKzeH2xZpzz7PoJAYTFiCSmD29Mp38W/Tq3Ei
k8aJGmx7WlYF+JGKzXvWWeQGs9tNAeO8NSGjm5lC1uledyIwPKaI/BBGCC4MhCNd
eQhTGIQPGt60iK66dtoIO6VzFxEDWEh+7sqho7pDJM5Yxs3/tGxjTHxKQIZu1gzG
EiCtLroGZ2BF1K9IO9mYUtKO/rhlN/MU+F14GFgiP7rHeYm7F1KM4+OmonabqKUO
Qc03qVHUR1uBg/jPXjc3QK9lX1XPPz17zF2GPW2iRw2nSm7gCAfaGbqpwFaFqLVC
KiWwdJmVACxSlthTzVuWO+t42NmozTnW75dHhHyxbWSUJZL1qm7Xd7MpgLpRf87G
DcUto0SJPpSsz+NpRb7dnv//zxcu09oxppUzDYDOc9RZ1MZao2l61fARHTZWQZ8X
FqqFkvCacpxRU98RmB4DSCAA4taEfp7eKKaCW5wjOR5hmDLdgXrI1amOrGYaHHKV
e2rTMp6aT4l6wQZlorIAcz1ly0TXavd1Hr+IBqYK+v66uarReUeuLUF7dnwTm+u/
xu2cXtaIm4NNBH1JNUIaJ1nNGnoFpanSRgELzv3/9JCVAW3GTR3yKsIYxni835n2
mfqQumXxIJguh7L4T5IHAa+e8kcW9YP2pyEoi3KDdnYxaUflZqymQUw8siJx/mFc
Hw8hbniQPF7P0j0jBvEjxXjLce/hVTZuXYzcvOA4SqnVWxO31ZTSq+zbH3iWJg1P
mFf9U2ihDp1O1K5sMEcP4k/EhAoYuR94FU7KO7mz/rFQc9aZZSCXygr2rmYesde2
I6zwA8fG1CpRzpDTyQYUVq/Zd9Q0uzku5M+CFLOu9RteZYJayZbY5evwa8tuxsHZ
86pe/0VAyqaFhZTI3kO2TnjKK4JTdjBtOpDLEupDdDihySsp18cU0+dXp8Dcb9Ta
/STZXJmTFXFtzdfSvkfX2FS6CGLYCtagVarqmMpw1rBEMp1yPcTyd9i6fZwKMwbZ
T4fvUwgz5ISnoF0HF1RCpKA8KaFvEWOZ037dllSTMaN5kVkjLZt3M6aL97iHAV17
vwhykxHNXH14tKjwjXiV3NtFMR3qvxs/hK1JBnlzX90dh1XvKkKo2xEtbK0222Se
7Cy4ACYvvSWoF8Oq8RFpFj3WI7ogxT4IUox1+UXMKJCVRYsaqcgwe+pbaLldjp5/
K0HoOOePKw0YATNBiFxyj9YCDq+rtEYmVI329r+K4fj4IRmS5R6q7XzxiP6C7JAN
9Or7FdyM4phWbglcUpTs0CXIHZYcmVWBwDukKHNJBDLz+Q1pdP5DPRcq8UPemCtn
CfsefDGJfpjg9UBSTYEmPdCZNOff/V0wsvovWcLY1ka/0TSg5T8hJ0OZjcSDWN6P
B438PlL8JhxP7F3c2XLOAyxVHc+zkQdpm50g4UjBBpx1NoOeBMbYzOwGs7OvOU/l
DQK2VPKfnWIprR5aN7rrhpeb4ZP3P1tIHt2b9KfnMYdaQtDD27Gbxuwvie6qq33f
j1JQNYOaaCadQgJt1b1T000w56YTY1F3rGp9GKoVE45wHFOqrIwFpMEHa4YGEQ08
qHla7Fbxyk3k4tY9+Xz0HF2iXW2IKK91VUU5pyGlzrlt+RD22Sw19EGZCZoJ6oor
l874Mw/Uo5waJWk6plmqgZsvunHQIbb1Hu+LRrJpzFtBx5NZzOerAtgVLugdpmvS
iv5sFd3o2HAxULd5+9lYHjOTkMZLUSkbQK9Z/XvwjtVh27b7KxSOycMD17iBNpy+
2EnjSCFDVDxuPGvO0vHaKzMp1Cr2dOkdPc6qR3Ro/Gd2QV21/srqXxk+k2eqeptA
mDYDnmCDYH822SS3nJyZ6SJ1ohiN8eMyY4/wdr5RQHLjJVvo4fMUIvk+Q5CKioa4
7+U2wTfr786gdWyjDdBOxFFPbbjCU+wIAmTvqJlkDpms84AX/EMPVCu7btjKUp+S
ZKTcpHiInm4chzInlw0cUTwXcyK3T53lH3z1z+9PGIG4vEA1KqjcRsl8M/4pNv26
xrjEnSwPm4SzDJ8WYDXjaGMGbpRBm5GaNJRZdkmUi2QAyHT9HH1SGogNOaoLxQ8+
5w+czfG2w6WTsjjWHQEmFd2ny6pBjYCHMCLG6Msmh7gjCYrXC63TkxW6AjXvuc5Y
5qAjqBctTFPtSTnyXKkHpTFdqsJzyTj9vEN3s+cGBeBaLh1VBYfYZ3vWPlORLlEX
GgnkBYytPrwCwut2VgARYZXY1iC/XPTqbDY56IrQlugv9Mr53NimnJV4cDUqAo2l
ZfoR1/Ja5ggXY7SXcN7jnYc8Lcg75pXis9KqErCxnre+R7fvAckE5kLDRoQxI/yO
gara8wsBZmXpcCMj7AusPEJGe6dBL34Cm3E0UoRG5+Cb5c1LSL5upnqLC5rJYsI3
2l3mNXh3eGIK8TGooElk5Tl5iZPqV6pBFNg6xmzOgB1oqDFGhlTtltfMXIm6U29g
A0+HNtN/7l86wKa/1ydoSKv1cb03ZEOqQVkU6RN3iNTel79h+pcrLl+rtF2fSBKh
FX31kZwCUPe2XeiBaAjZSnuk8HBgOuWjQbM08D2Louh62/CbYtTbME4Xlv1fxscW
K29O3zeBtxQrU8v9KtDN9tDw1kPVGDnsA0Kd6BkOFSW2hu1Uoh2nbeWqMSMuFwj4
QhpML7qzXO5e8SEAua25J8PeKGC+cAbkuIufSSr8xMrYrHKN3XJsmW6B1OSthOEf
wUuRi2TU6KsyugS7kl4UF9MIsqrVvCChoc5gos9BBKDI3kAPNYh5/vJNEsc6axGv
JEQRAwFIeVlRRYQ2EL+pPClbxFe6Xhuz5IpU1zwCKvW0M87WY+kF9JQLxx85/+vj
4Aw20JHEr2dO9iGsUvVsvDsKvxq6gbrFIrW1uj5Sh607JRWbH9ViKvGK0KSIDsWU
QIYqyA+/QGfIhbAVpP+s4/RniWU8z2dlD0KJBdbLll4CWUfTSJF9x7VyqummUCdm
7eBHC2BRPLFAH2hV7eL/GAqaCggEN03ToeMjYRzZKGIPXUFtOiZX0dFqiznw8SxO
XvdnwkUmSMsdvhqfSEv1MqBU+d2AjV+Zwjf83v6NOT+fesd5sacv6JsnqE61vlLc
MW+MniuXu0966WF7aSf5dFSk6Oo51qsORwM1o8sPUpHwnAFbM+K8wBcfQE7rY63/
Pn/CO9tHLVBVBRVp3isN0KQRNZDnjVapm/mRAFcLKKCqm7tpkFlkRMmiyRHS+qUE
+tSiIRYC2SlI65BMHsTRco1EhPKakldwwRdfHeYt2+VbR4+ISjf157Ka4uqxtpd8
5zTJVQ4VYdaT8sJqEvx07GDrw2d1NVdUvEs2OvP7vNy1DdO2VoseDXVfo9GFcjbU
UOqSdtg4ZL2p2XKgzsaZRzUx1yuCi7re4mY509gRa+rWQit1197vHFPO8vTpjdt8
2LIJQ5nKG2bMn18qKXJ12TNVIx5FAfCIACWz3BOAo5RzbmA+HIPRXqyd0DvWM4sk
yq7WPR9c/TB0I+lW6SDguUGgjbIzjFBEBa8D/saYoUsxqpJVx4JZnhNb0tFTXVFH
ybew2TyNbnbvb3tWn4HvBjlJxM2gXWELDQy3uW9WZUO/BOrozbL7YUZvPGRgmdpm
NxRuIrHk/BZKZ77dfsHX5bkKrtUWg+G3qeEO6sWKDF/zk5TnUpvFYmp5j8YglzaR
PO9uYmOOn406fToV8k20tOkdvnseuv5Ckr2dp/X/hyTpzTq6Tf3LxyCHJrJhHk15
675WDeAubi5PqFcsp6j5kyPLOjUxXxeogvn9hbrhD6JUhAbmm3zdJbaXzUvq9ZAg
0GrbI/Jr/d4Zwt3COnG58R4g+L+MIN/s6PZaL+e3DwsOmex5Utyt69vUUBbZ4iI5
1bSCPgBBVFFfGTfnaVHh2CVXs3Ea5ixR2tVBa1PTygbIG1v2I38/PnCArGR4Su23
ulUWPgBoK6KnWolq7eDmwqVe9iQjF/FV/igOtUPvGPexVciAn0e3v/3arGce/DHm
Y3QTlE1J/Wf0waw0zEEh9Yo70xMOckn6ojy0qRki+KL7w7lek0OX7YZBDAwi6W6O
e8tFuGYG/VbAL+9Lu4yncacRgiTG9cjTNMJNCFCpKm1FNH2S1c5dgRXpPauBlawd
Bik24wkT+AEWzUCVUuS+C4DymRCUtKqCC3gFIu3RHYA1rkSxEFjiElaDwI+XJ8Ic
I6rDSFcY5rt0V+sUYDcyR1HCtPvfKnA7K+veKXu0t5qwbHuCew+Tp+MbodB4vRFX
OwwBjRIPjMx6opxVtdIWtaoq7n50NdsDJkNtD/atTpQgT1zWJyl+up2xJcXHK+PF
AE2K5ciZqXVtGVEdTjaWfcNww/N+/JiG8MubcUgy1zQrSbJAtRoON+yxuJURF6De
jCsRL0C/NmEwZSFeE6Ha+ownnigeQxT+EBOqaHB96QEzF8b+SPltMvn/kbqKs1N+
84zaObBkIO2+XzJwOqH1XiWha8g4vlnz7MqEQ4PePlIL3yYEf1R7skRKA6n2jjMu
zwofbJwqRiqmw5nxvyqXpXfbV5+EPbfj6/3mFb35k/EWwHsSlqWOjn1+IatfM5yq
8h4a+mpoJO2uJdBsgy5vuzghmzS5OOI43FnCNOb1GzgOU+e7PBHOpsXNHV8CpwiH
bzfcG+RvYTyL7K01YHHcATcFacuarU/FAXFgSPx/ow6JoN1JEB77NXYthtAowzZp
T968cvIjuhYKoOcce4pOaXUi3Kxb3Yks4AHgpuHZl+yfmZZdr2eS7wJcsTiXbk5f
PQJcvgeUt0VrIUcqtfbk6/uD64lzTuQ21JEqVVdN+E9U1eg0j4apT0kE5OH2nqUq
iyIJYVNI+ne+IbX6iNSu8p6SXJf/zON4UHXLu8whmrfvx1kbo+WsS4rrnSn4kKu9
zM0oZMAO9CYXgnDpMLM/sF/AL3+fN8JbN15fqY2KefprulDu+2cvjt+8XOAsL0fo
uh0B9FkiS7GRl8qczokmPn1/SEzD+5bcLI6HXQ+Zfm2xaLnIpvHeERF0c72eLEvl
9NZ+q9Zsztx0moTCHkBow1sF8SHxySbnYLwr9R+JrcaxtL3b059FtDb7CdOCP4pt
oQlHvjpHfdCsLQDF6s9HqCkiM/OACe5Ge0QMwL6aG+ncp7RyDmcVx9+1Z3An/Tjd
w8fgKTW/kIo9bJ702RQdPF65wIRGdXIV1IiYWMfMvJ5HMEwOuT//CqwqajyRs6pd
1IgXBVJA1+xLfSVX4nB5e4uGQ69XRooPLyaf6W9QV4JyQhzJPyUde9fgsd63H7wZ
sSBAhIt4dJDaAcTzGD9WjMbNBP4nIXvpq6e+jHPKr7rrmQGCiL1GNQu7hBcG1M7I
0NJhUPrOLrU45yOPNA7cYizEHh2xH+dOkT2s+OxOZ1CRXOgzCYFkzyuyjosYHO+j
Iuwp2XOubb6+BM3fvUSDvqvFnOby4lKXWIRhioQaTYfdhJCiy96SNGDxLZRiakrE
/vYbvVU1iOGLXFVlPhX54J24DA/bTBUSyoIysmUS3arH0ugggSQITTNRwAJyEH51
zavmh22D/qEFRhqrn+52VgjVrq/6QKn+ZyjyZ4VAEFxGuAgx1SRUu9Fb0tGnCofN
Kyla89AMtEiZq08NZhjrVq5jT83zfBSA6I0krXveOU9zrktc7l0PdAOYWCRwtRoo
eFL6pvBwZoY0wG7ke/MI2FLWHxalSR0bCBHNJW7u650J4rdem4npzcR93kpIbW0v
wobeOIC8yM8FH/yyx5EyLglJcsgGSUGtPB1P4Ue9PFH69o2524Prg7taPFK+FLCg
+sPhWFkk0/lfjN3F221YnIrthQBQLAH7WkhIBh8fWbr8aurJdIC7/YrAbY7tNqn7
57HFPN/AYsMrXUZ80AQdDCy/gMX6R74Occ/n7+DAgiW8KNMKwFZfxFYa/iyM5r8F
d4mGl/Aez+heLCIEG2Qg089dxnrw7l67Q1lFKSnc8BlDsbFkpLHjVYmx3oElhpPD
BvGAwpn5WZk4VdCZ0poGI9KD3Ja7hyB8u/R56prAVBWhbxV+MoKYTRrAPaU2w50f
79lgBrN2/RFqGXYxs36llU3P3p0T7tbfc/qIXS10H3Nx74df7LOUceX23UL73Cfw
BG+MtQw2/VpHlNBiBy7FcbyYqUYeJmIb23u/hJb0X2DJTeJsUECVDMqkxXWzuZdt
AHa5TCf7a3UDG27bV/MnJxl788+CTI4s+K8q3JZbVBwMAO3mOhIRQLlIQUSMNFNB
C408O/DOup7DiTJAbyctKHXHOTCov7byYNYl7Vh6lnzPbxlgdLL5vbZpbq0HZBLD
5FrYMHNvqjIL7Wbdd0uwX6UoNZLHdErFU6rLyjiLprwlbX67NLJSL0bcvtwFDVyy
mu7QN5rXc5moTsy92pk6ISRhkCRUvIj1epsy9J/m5JUylGvi4F85MgHKGIx/oGcT
ggVashiG8O7+4yqWjNm5QfONarorGgn9aMPZdRRPtf9z+pmHiwvpRQkvQ4lnpnRg
L2idgBKZGH/eQdzBhzGZ4OmxuWnYfPVERWkZwbz/WfRXHdu/RMIIIWPjBrsUNt+C
lP5fPfD/nGPamEg4Lmy9Vo//17VSzO+aWMP21+zok/tMtfHaqgvqC+/WdWIuZcMo
W2SenaikVJqGhh7qbHrv3wJru+/KDuqEqflqFur3SiwdJ3sKKvKje86MrR95qc6n
0OKJq1yEcQFXw7ix5NUhgf6u+lzvMNFVOVlR7zv8U6SENaCnBJNK1IRnll0VuDJC
ynXLPCWCynqv7OaR4ibMRyNmOucRBaMytM+2W6YLsQ5ZBweLmKVDwNJ0FSV0zy0q
8zIa4SAs/Tg8oynj46hGmQDn6gSifNBtzZUvsCkNN/7EH6qAw7yM/G/UvNxjcYLi
ENVNTei0n3MUOCNrkIC0T+ZTkRpRXmvPedUtXi1YRWUdusnrcPn6YQPRym8r+zDl
0+Kg+UkqKogUVzEHV6XQyMUiDrjiGh4tcJ00WG++VU+808hFId0C8AfhL79RpWd8
1blCqBr0Earm8rITq1kM+imRCO37nFAck4FppgBsfbxGfY3HzGormzLJ2cvnlF0M
rvbm2ipXoeBPbrCWgrq3pYDFn8twASeOA3csYStYOATBYv3WTYWD1rsed8Iq9mXd
IDblr3bQXvQ4kfkA+NuHz5RZwH2FOPJBJUjC1/DcLPqVOV0CVJt87Xs+wycDbi05
klCdzZY6JcwsvU2OsoFlQy1b1BcUFR30g5ibPEr/0NIscfpr2pvtL9xvJ8nfcaFM
yNGpR6UlpQyMmbyKldewHkz434/FU5rNW8qzIISIoXP9WTQV7Ppl4p+LO26QLQ0Z
UgGrOHperFCc5p9L78h0dmry8Czs3ajCl1AUTbA1LKpY8shJCc8tYvKv0HFAABZ+
lOePDPi7ifbvLtGnGq8CKfDgQbrqNMxxQg2GUDwfM1Zqk/kZVno6ZrRxBLNMKsyG
e3QZRNLvwcgzbayvd25JcZuaRcA4dIoTZkEIzb4zs60ZLvwazWUZLwM5K5qDLf8o
nySvHZPCxQGVSvPPpUfLqk4mMdT7KmMjW3XNSzMBLQc2L+M2i9tgvvhQsY/zfhfW
o+MlQBhsNk197adhtIXJlWqn3bCCekSl/ZQznUYW5Iu5eTBKYKAdt5+5w3ZBoho4
eEIqQ17CzmxzNSw70trGdWVYOHXkt4rQT0TgL/5apLvZ+wEMUDaiGFZyexdTePg6
LBYjLF6k7B1t2dag8Z9bVNl2tkm15IENzota1Fp7zlp4v7JOmZHFEQg1733UkVMc
QAUBfFCewz3sh4qUXyHE9PuhxjFHIKxDIibBTziI2+BmnBn4+NDPAuDApH70aQRQ
SjkcWH8FD/LyhCsak2InZIiCTTIDJmE+Rp0PHLAxq/y+FZXpiEk3MFTSrvDYbhV0
g5vE/q/SP+4rNd5PvC8KZdIJdpU3WwRw9NEPjcHWn/jue/se6WHNHzjLPPnzlYzr
v1bklz16/a/4UozQWsOtO+gOJmzp6ZI848txyA58szpTL6WCIW7SmLZbJSoShzrf
lS8+QJl3rgK+CaEkN6cL3NOHBhIEI9cqMbjnA/HYIKgUN5dF4OoRvDhjJgZqHg1u
bMAZR6DasyngnsYTRj9Hk2oX+UpznF76OsV6SbqEZGOrtufR6G+j7GVHqDRjAdVX
qrSywhK4CsWyg07ZA2we7jx4RCUw4JeUk9BdLzlWc+DhZ8J+e46VV8PNPi+ZxFzR
nbHTTPMYAlhUSYPYxEISZ4rRfzf9O1J+DalVtClHaJtv1fhWYHFa7at+tzupUBWd
H+KO+755PEwY5bTPjJlLvL0ucPBlfNtUjbxUp54PakvPsVZ7aCia3NEmtHUjknvh
naqhu8ewhFl8eU2P8q02WtK92PL+JaglkLmsqwJCHStBz21djcXZYM2UY3i+2hne
Gy2JEqHHXBx/jVN8iFO1SYJkjKoXGxIXB2jjfVSloj1NNerMQggtg0pfxVCPc5tU
Ve58mRRPiLzpw/mzV9My0X4HrG8TBXhyHIADPM+9PGZpy4tPVf2zKwPl1Fioplas
d9gSi1bKnD8JKGWQ6tr2zC6sMQp+tEFD8gaEmNkNiZIz93cq/15DISaR8COanF3L
XTNSCdTHzqs1zp0GIkDbFe/2mvcALIVN/s21HVwu7M1R6kk0U6cAEV/CGFQ63vZs
qWaBarrm8fincZY0Ha3SETYPOFJCV+oRjWD3mf4XMzKIEOarI1wM3G7HYx7LKs7i
3PxXcKtyFUsFJ0c71Mc0OpB2CdhAHsu+0/cOV0VVZxQAli3z0eAZamH3Alj2NGcg
URWEZq7TRMVjWLqiZj2/lPNbIxwWeSdFymkc9+QIhk/deS9A/UZg/HAoAx++2kMP
TokNv2pyeO5Z/bpQjKbu9Huskd9pXvt/IgfC3NdQCi4g6LYfI9N4vwHJnra31Sx5
jNuLCKgALZ6JeNqvUZdj/GiCIHO0mYXefhqEgxFEi4YskyjmpxGOMfMPLWSOC+JW
q5fuG7k1msx++SahjgjNW+HrBitB61RuHXTSmFcBtFZ1SMULKjqMqTsecCMNktuA
Jf5Ut/SpFQESIP6FFSPurnLLyj2RgSnZN9wa2Dd0GeDhoDAIJmnuhfX54WoAiA5m
AajHtbhjYfS9Uw876O+glIvRWn8IzC2n1bttzo3wKRY18JVfxQiGz+sH4BRKbvNH
nA0fL1IKbAIz8P7CNdSJBiv80zpQaMdBvrBTftWxps4blTib9+pUG891Q+hkO1QV
ytYMvINT19btcUq2/QdmjkSlndiq2+KzpnKSrAWd6enyCqIKWll8rOQV2epHeb8H
t/DMiZc8U3lhhWygK61qta5BvzCwkoSzouqM8hd6WwAGq5zpa9KoxP9Nv5mG3c/L
AWELx6GO1EMN4rlDXDfByIsorAlBJP4udZO3O7k92xzTmTYhMxf2Xhsg7Rjs12A2
ARxE5W+lCHLSt7wemKj2rLE34B3Dx9s7kRrFI7B21cPIK/kCOGYdlkRz6Em/bOT/
ywlpOL3iMpQTHtHYUK9smxUVUw7ScYBKxnhMtSr+dEaFdCcLMBK5iL3EJjbpF5rW
IOeZrmoBR1ki5CZ7MiHOeSBfEF0+SNoEwI8tPBJkBm71Zjpb7v7z2qFgwkG6HoI3
TFiPFepeZ21+pml2WGcTBxSyzmK7MjrJPcB+45XsjBCwTEjReuOCCF9vIeSHrod9
lg3sAjyX+XCYhRALGNXKCMaXgx9tGXZVbul3drztfp9rZo0MUBG7QDEC5w40JxyB
xIo5F5cY3wpriGF/PNkAfmFBeA/RHMX6Hc2ybv67mXjsBp47yT0CHmgyZOpaEtii
ml9YlYcvdF/wxBN/wlvSD/OCbNr8PNlIJZ8iQgaYmZksvz1uHU39U1sEJkTwlzie
1yGahtiTX+i0QGxeyoeuYBhTKxjHuxvAVGYgRvbuAKodGiTRAgzzeAx+bcnn5GgB
dGAaCv1eSx0QpVo7iDsTMrHOIJGtiRFxGPIZjNLDux68rN+uqcnW4GTikiQsfeOz
a+goRr00tBoQ6xkDrLy5ZzOfmb+P67GgCkTmpD8RqkUJrDnmgmuD7XmNz8JwFeAw
y+hWE4sQyCM1mdhGEd5kL5jDXofm+PZ+Z2/sJvOAhLmO7cbFZNzcrw5IQMZLJeuW
ioJ13LPZOaUKD8iimKh0cncR4TUYzuHEq5usWIsJWCbT/9rS4QdLmKmRKOC31Pm1
b8ezBmp49+Y1I5VB5j5iF2j/v8SbX7eywaysgW7NTCfMzj0KgJ/Tijcof2iy7ZEA
h3Ta4AII755rcPc5Y17RcU08WhbKf6yZQNlVXdjNyUP/xqd2iJJK0WexiKGT0jvB
+7/x4mCUOqlO4RznR5pxfqqpEMvsfav8jx2bDenqmpqoXHHdXFxrRIOSIn+m+nZT
PeDHM6NvrMGMnXscv+CvKpFXq8iSLwW7Y4dADfFaYdzB3Rpqn8twFDYbKG2vrFno
sRrMtdCVM50XFEo6+mas4VsVL/wdZAtJW6YZGDpvGlLFjyq8orm6DEuUrGEChNeL
A7CTbQ+lRXjIm/YOjq4J2YGNfw2hL3BJTEAb8bQYiNwoqvsr5ZdK/TonotC/xpCq
EA7XznfH3AeNJPXSoQpVJUJ8iRWT110ObwtvZ5bCGhdujLWNXackew0+J9GOs6+2
BEtBoEp91zeN2ICtg4FPvKTFVGLAGKfXFBmwbooHJIRy/vCwA+XpSuPRt05zYBzs
YPWk9gTNWmLJmCV9JeR9JQ+/9ei3le4KLF2JvSILOR/5tHxkZpOamj1zhogZfWJ1
+H55xFXl6Rwy7bga9ozkn3uX3l7zjaQatkPHqdDnsbzwNI/6feRgITFz5m/AuR2x
NxtlWzEdFx0s4OmLNq3PGcqGlcKabX1Hw2clwW2+ed0lzek2iK5T7HoURcyI2DMy
TqYT9oxhEfNQjM+yJGajadeRh/fqPND9YQWnBY/pxAx44dNvRhfgstO+UFj3xOkk
1fImXlsfxy/RQNGhkH8a9a5Ko5bUBiEsYeJhSkmgVKL0Z2z6Z9i0gB8W+lUFX9ut
Czpip9KBLBXKh5VI+BCXm9cmD0mhcvxVSXGivlOSVaQwf/uJsQ82KGLPDwoKMqBu
A8nGTC5nXsS6smnbcKHiakOnQf7cUG/MPDZfnGfTike+4gwapHAiaVHUIhgxQNBU
rVW+dHYED2rflGc06HreAyP3Cc6DaKku+FTW+5JM839u9gYsk/3zZ56vejuFoy6U
2iiEuWifXIm7Qe4yWoHj79/ZUtMnZa08p+ltFtSehuAt4nyYLlaSu7M4DjY1Czf/
QlCFk8AFVbvQhmSrHcW7eZwfuE3AeGEHkjFvKoBn4Vdt2O2kUyawenTLWMIS9MwI
r29ivRmIeOG2P23Y8kwzNdNPT7DvlNvRI3Vv+wcbbZPwbnpy2Y/uhEjJDgAddtAq
lnLiAinaa/LemtmmySc+j3J1j9kMf+moqqKBF8j5iPiGGOlQpp0dmkzn3T0DW6mU
cB2eiswEG1nRMKc3ZXBunVieBWCBRew02COdIFWGaMP9N0+sRviygUP1xZn/GGd+
27jA00asR4h6pjnkuFUQL8vX2dQgvg1Advs9894KBkvVNh3GtMys3FRQ2dRu2yw8
jDS0mYB9ACo37WPg2vWTZGviJbhT0koK+vY77RxJLnWgrHmu3zbsgDprIyCljDtc
zh7GTK9O9gkkRPsr6FAh4te0YXGvVIL9kwZEX+vrIW8jkulGKKkGJYCl3iZJ7sEv
zmuRC3FTIBqzCfWsc5jmOjKqLwy+nT+//IS9MYnuUgnahhq1TB2LGlwzBXvGEVj6
635l0GZTrMtrLYN2XAKgwQqTw6HR/+0clLM5FZuPCWZa7rK2csffz4enJs9Tlcui
iKioTaWqxU7apgYrM/u6jOs4St2IsSMaC1V9AIzRgRWJkHqyzDKWguYat5HAsMjH
FMS4AXKES6TFJfinXQkvEyDpfsA4axXMwy6MhwUwOPptGLsGU2xnt1ID0htqYXyO
zbCy0Q4QtMh22DAfdsA7FfXSv8toi7Lko4K4TSA62LKiXev1T6D12KIQwrIQDh5b
bi4WI949etrghikHi46KIi57NdEJvAOPMN2sbGWZnwJV2gQ1YPhqE2sKEEsilVNn
mEtf/0eP2LducBufREjewASmKVaEWNh95jJOF6jbBjO8mFturqEfLvT0JaTgC/7q
g+I/RX119ZJwdocKDXaDnPWZGC4niuM2+oxqgYYxsBMU7qysLuFPAJRZpvQohRtH
Cnwafnd8GVSmIWsW1VBt2+o8ay9hcvbwqDJeeYnneFQmnaQC0Hy3Nbz09H/RMWla
toa2vsOmKH35xJrF+HN5/pX0yDp4HhJZ6Ox+aCSmuGqO2xhxrgtdvf0OgnFtQRsu
lEecYyJuNtm+kgcikP80RMd3VLOodQ9lrg3h0ibOl2kbD/oLNZyY89sNn+pqLn4z
yjmpWC9OzQee+FWljotWLPVUrjlIVyXzz8Lkm+q7R3PFGeD5aTLJGLPtpQyEtUvn
zJ80MBZN6wqjGk8JQPKMOORL5jhZH/yEn2wcxkT6W2TEyKo+qSn8QCA8VrKNRk3U
hLhlX0NKIrLb932he5g7/uZL+Vhi4rp+PIoY6OEMwNGvLIaivtOeo6fJhzWvkLp5
TM/khm4fAaoc0r8JHdgOcBDUyg4Js8UIrZbaE10PAH3ABJjfuD907qp3Wa0W4WAB
WUD4POikxrt04B/0QnQLNIISykDNddSFz/Pnc53Hr6UtpMss2FOVmXu3gNmvogYt
GO/DDXkEOfzOhghbGXKq4SBoH/vIHPgntNq3GzSQEaP8mWfYp89RimF+7LnekJg4
OrSdWvIbanq1aWv54rYwq9mYZ7dz14FR3ADa86Uny9C7ROvxA3WK7Z0ykOgFw/dn
20FwSEkhWXM1w8aFvR6fXlERxLIGx2NzYGdcGpmvJ4ReiQhHeExDZeL47Zvakiip
ez45R/JsxUBoJRUlg8PNxX/aX5Ckr2ERlAzO20jRjceOZGQ+pVafL5r4Z0pwxjEC
brzAOx79BmSEiJ9Hac7an9rR22ek5gWBgaUM+4TexJWZ9KSuxK0JrWU8AMwwXy3J
RChhl3kNMwZOYMrfCyqoQhFXzUoSurh5APxfIi2jXHEWKiCQCk0jgjKsk0SLE/wK
vtVSYkoMkN/009QvwSWCK2nCTu8LIqxLWRPUdRS/g3N59bgCTAqGT+hv9neM/Igr
48EhNHCwC3s9EbW/ohu7rEBtTJw6JQpZQLx4/518Avt0nWf+BboiQIlfNtw9TkPK
tWji7f1JR/L0MKiOyTMihNZ4vr+goD+Jrri5zx+9b0RDqQE9UqTO6+GDp5vZtbnS
M7Z2ixVyTtFSwwHz30tFwH3TqhPvNNuPh2QvTDc7vxvK8XWgzhPYyWLBKbcmmez1
iBwdCubYm60xB3QLxFknFKpXXDkB3FVprUZZUt/rAPakdSor2SoHzP5G3NuVVJq5
PZn0xytvezp6gDP/WKboIfSbRu2AoAYjZHBeE77bl4Y0/f2eqEKYmNaMxOMIWwMa
y2xWVSVv9AZudHtDCy1HmYuB43V6dfhWRhlJzSvOn/afPTkAVU0VZjgvPp1riQ9O
DCxKMq4WqjnuP2t2IJ2g2emAPp2cdPYOwjcC2MyB4UiiKehEvlEHhlHPzik3LKWs
J8WPkapk4hlSbmQ/bklln1v6FTdM8LDi1I5padfBLxSB+5M4gWMZNcUHFPuTyZVM
UN8rsy4HY/eMMZYfaZRXXwmgfyl/TllaKns0ucKPN+6XYEBv1GjFSPyQNR7glvqO
HNJmqNAc+sRlrCbR7f7aQaHH4Ykiow03wnCN0dRgRVHMF8Sk5AgjeWQwOwmvC2vR
KCa7wcew9gbQ5VgXzXsTSl8TNEnlsK2whGQx+snuHMnFDBoFbXP3iXd8jfgA3zcM
e5FjAvLckeRTCmuhscxZmmEeX3ce6t6rqvbTzrzDAYUFTgiZMGw0Hi1JDIsgNRO5
Jnxn+7U9LVBbLw7WlWTMgSJxeQwKoLrodWMjdsbS4SBd797UkEq0sTH+um39OIiQ
gW/ltPUNLCPvHwpd1yDwsTitoZuFj8OzstDIvlYK5+gtwmXvtQ4YkgvrIbL9GXwa
7RDYYKzAIcdsDR1Bs5D/CEAiXAJij7QIA2PEG8580iD0OY3K+nq8qqQggbMYgy1E
9w8UnTh+LWrtmN+FcnurpQztBtTCv+5pyL4ACQ9EUePkPiWhiBwsP52YKeXKDz/h
X85fPKbILb9FvbgC399DiwtCBdl+Tq/XQ/FFc7PlUncQQTcMlB6clZXfQcYk8MZe
e0QdSIO27DxNiZPkMyXSU/CqvQ+gpijvUbpVF43tjQ4ZVHDmff+B1QwkDIdoIIOY
Pcvbu0iC1IlQ5HKEzX5W4W54t1B4LKMQI/hp93vjlYHgzs2iAN7Xe1jJD3Bvb2CN
M68SYUjwwLecuVwK4HlZCEjDrhTEbwgYeHWJQ2FDFCo7IohI349gQk+7K8MPqnv8
cERGFhPGzVCVtQ+vtf1gZGbJNBjrtYhrzZ9NJPb1wI2fXYYWi5EednGUcvv6YioQ
NWiW7BXSnDZzmUl7g5tm8q5/H1ePisl6tEJ3I9c4JtNERS328h0aRP9EzKHTRTuN
2AfKbOAJhZ0OxTtC0XeCxv/X5gshimBvRxo2kAJ18SgsyYZuMTTE/0aWwU5ECG/Y
OxZo0Y2EJl9EA6c2+S25EPN6S4tUstR892HAKPazCO2OqHn+Y13PqSQWyS814MNb
V0ntoGZjmFZyLl//DeMqFtcmwBe6wc3/QTYoOu/orToMp0dKiPn5TBJYZNKd8nDb
6gCcVjcBrorFxBzsZYEL8O1d2oQad8N1d7Z8QNrl7j5QdV+/5I9rd43C5WZhghAG
S8Cuga5wMcG+nwnFhWiNm8IM44bCNIGfnCPNptNKfe56nxNSM63Uw16a+X4sL2Mz
ewopPbG3Lpo7Hnrr77JCx3uPzU0Nf3AK/oMYf4fIiQFa2quD0/LmrfXBDATe5AlG
zwN8dQzfXjYRJNBHCjaEl3w2oCqqoySg0KxIp7r1eEKjueKREWEG/m8oyeG0cCU6
4b+7yZ0fJ2iFHK8A2JqSMxZyFJ904gR3agUUfSZk9k/YtQFGkE9RJAXxrqUQra3A
xd2oO9wZBxkC+1zWADFnZyBQ4dFArk0RVGv6aHAmakcOy8NH+scedWdiG9DN2lEc
U8mElrUNosceSJ7xgpXwLJuNJTl1GJEe2FrORM7N8RKonU54CmkJ2bkJwwuUNEUI
8rnAMdqbVi9xWKGa5u3LUSlZjFph88zzfqDWBDV/jE4VB+a3IvUa0R3dCcM4WhdK
if7NNqY0DTz0cMMstKlByL6UijrtbqzKDB0xFsw9j88MGsB0ymwBL8GI9qWCc8Cx
L8YgoPJNC3EKAF//8+KaZ/QpIhb7nJJSdsWixxJ4jxIIri9nPVcojtYnHbBaw7FO
80M5cyKzItnKG7TOK5kCjueNnJb6wmRwjT3Xj/S3iZVSIDA8Fnsp88/Ihh1VawEB
BKF+h8UUl6I57kdIqTXtp/CvXpZH2vd0z7+fkHGV4Atx1T1mXrI0762QgrNLOXQG
gkmlq5/tmER8oaUhprbu8nDqWURYPh9shlHdb0O68Mjuy7cJ10Kh+LbFpzrxCsDO
KDIBcIFHiAxEUHnAs8FEtoHDYl6VlOlArosg17kUhp5JolEjeSSQX78VJ7zbXK10
UaaawcZUVfQdz41Lw0RIvNMh3TUMvtk6Bz8CsBo4BVs0XPBd9cp6462JZ/UE2n8N
RxenQvC50u45SpWK8e4N4G5kgeoTwqPQJ40UktOQG2jk4A0oUPuLG0rStbZFokmS
nMSgUzkReTbl1u1/vl/iOiqE3NRjlcrfcVgwTDyEz/Hvjao7P9J3xDO4GikXl4IH
uXND0vvy7iFkwNZllgbmo7R/++JZ2fbBfFR6Hl7wQ4wkEtcsjOpHjRYzB7Do33TF
3elAeRhYHqRMwSD9dUcYd+2QNW+7znGedGtb95HZDk5FoiOlpNlaluJcCdgxIndn
k3H2/eVHmev1ATSy0DYtzIExDEVK5qDYGgE8hrQRCtA/OkTYGBBoVmT12W7OK7l5
c+Tymwzj7aOaPT79AhglXFH1+A8ZbNwvXdwrqsZ3usqc52332IKr3sigvo5iYtWA
/MUtaqjSJV1M5ljfVxTJiVrPfM4gmFolqUuyMHI0UNRyBSJLV5SNlXk6UNTPHySf
NL6Gl2b8pav9ufXuKZ6PP5568v/8cpwCE5ybr1m+4bkAIOYsQ/2IBlZy8r6gaHXA
9eBdJmepUXi15/Wrt+c432wQ1P9uUxPxIA7BD7D93wA0RFDg7q3pypa9gWVa1n/Y
qXM/d78ubzfZ/orFdXzOEE40TapGmB4RmH9nAYuC+juLqGLac5RWe6nE4W6SI7E+
MM9i2jvKyX7Az6+jUzbY33qyHFU2DPHOFo19SIRl0VwWTd2xf9+xuWFRZ4hmmyNz
Sw/C+KW8M8IFdwraEnUpMq4gxL+DZrprWV2jUswdAwd4SBtEIOQt3vv20jRNocgl
FBHtD+X7WzBssA0QQ7um8pCcar5RocGun66qXeFGQCegOkm7iIUPWPqvfhBz0iPs
hAUUrOktOSXGiRyn5kfOECFAp+VmCHpKELNHFwzwajnf2u5xIBdULHA3lBFQmESM
qfDQUP2crMQ+Cvyd6Gr8hQAWqllk2zPMSRtut+YEvj3Vdu8L6JVqZCh2zHjBcmo2
S6FYBKzXFL8FJtzEHhPGi63QkrXAhzpJmr0OgJe0jh+zdXotuUMBpddwulGYHnem
AqiIe6t1BwqBfxn1PoyIvR1R018kgg05QQqaVPK092PA6wbM1/KREAJbXalTDB+Q
9U4Fus3uys6JzU62N8ZR7CkylPbIoGdiWDhthgCd04/0CNYvpAIDAj/L7UZiOlBj
yLJpX1TQpc2pfdHeHFOw4dJm6c3x0dqwX05YscOgr0ESSFf3EjmBUcV7UOT33WZr
KFkfsKotXcyJsLkYODmHGqAO+WZ9zKvP4gID2ls4GEdlTtyD8vQc0XtYICERf4pC
oY4GXldL2M7KH8Nr+Apvp8N+EJWAdfKQMHDMCmC1/uviqA87dxVydoTzaAMf4BzI
pZHMfdXiD8+TWYPhSszqSfwzsx+xlEmYBP58CB8hFvQ0oRLF7pEI/n4iOtjAf7rm
QosxwHRA7qM/IB5IMzkXXJlif0ToyAcyUrZlQX/dfBXJ/3pdP4BfZu3h+3fC+0FR
ZC7pYqUIVn4qptn+R1ESqp3gNUuQ5LYBmbmpoER/RxevBMM8SRemyAR8yYt09CdN
owsP7RWLpQWlynN+9Uhk5HZSecjJRmxRuooov4sYcmpumvbQllsW/DIvGxVfHgSv
dsc/nVvKOnTRKA1gca+R1urLW3ZHL9c4LzOwubWntZPeclOtKv3vT8Tm++cLh0K5
MvOpzbKeiQktWeLWvxUY5EGtpJc89njPia5bNFUWZfx4jpE6mH7y40q6Q3F4Uqa9
f7Fz4Nsoy7YSYe+zaftz1cMm+fsh9smlY7ywC51Q4kL5ZstQKHUxBCaIwaZ6nfDN
XQTZTuziR1MoIYiu0sE+XcnZDDfOH67rJu691t+hqgIr8/LN5POOUnH3YoTwrnfX
j7+7TVbWYPYZWGkXK2vN6jSnzJdVf3zgz+p4Rg+E2loW5fwewfwuONhTO7KyWc0E
T7+z1izsFM6M+CEwC4p7lfklNcoevrVLnn0R2cgMXuLpEQQRC+tAstAVNK76ceq3
3lMB9+/Z9661AMKJQuehiFgOnD74tqhxvJKhoWtaYRMpxktUiTn9aCv451T6PV27
tsqmDNBhEqKMkqIMjCGZhvtFZW4T2/uCCsGycmOoo6fme03Ne/X+IrbDX6OV2G0x
R2iO/n0foLdJkKRenKDVHstzgtmsHxs2kCWTTXCBCrGKNnM6ZQVi2K6Op0vt+uAx
npA5OP71C5D2g/NpRjp1CdOyQhwzcq4127kFQxjUGh0q5Z/PT3j2hRMVcjpHDk6P
mu9JCfaPO31/Uh+UfuUI8yLY0Z2g7TGGEZEPVMCqc1KW08YgHuE4JKs0PAxA2pMU
gdBDbOkSxkelu1aqroSQOq39qD6Fzf33r1n6MhTdK5FTGXBK9ToF49Zq/2aHbsXm
5CkxmZYR6ifIWNBH1jOTv4SsEHgDirqMwimDsdmzpAeJMCNwcycYYds4GUv+pZzI
TMCuwmzAvehw/6w2eLdor3FrG1hoWp5Uq9ASVTW/c8IEIRXzl7CYPjbLoWpcjmYY
GDY03Ek0UGN8jNMkWVVD0vlih13vplG9JU1c8Y3U+/XianjJEY90rmuSVicSkDSm
nUfVew9hoDOOEjDkEnu/ba9IVryGVt653+npeQm9MOwNHJcH0FiEo6T/14E+/4hv
6EpuhAzWW47k20STGObERzmCF46RpMT+XRFWDvr87/We+AnZ7kmh9BE60HoA7tKr
RwJ89mvBfRH64VHgjo+Oj0RBBGOBP4n1Owzaub90N+QviUrWPF5oe1GtyZwRNxeo
TYyC24SFok0kMNdKgC1TD0ihDX41sKz7/w8iJ76TU8v1iSISrDAn3rxdGti0Xp6/
xP03p/VUdsZxtEgdYRpjYfXoYB5ZWkKJlLPo/HBaTDW1Om5MtuSZKFyWESqwwRvS
hHCQntcpn6M5LQt+xkkl6dVwy4N7ZmoihAmrhb/icEDwydV+SWIi1SDxIK9tj9qu
schoarXycG8gBRt1uyUcoAXB83h40fzODfA4dLkMaP4ST7ovBFHFrqJFMUu1SM2j
jkYDgyYfCsyyeZ6nLe2D1Zf1gZaNcjxlrhJApahsIic9f+q4zq58sglSq088Ijzs
IPGPoyJfLQ7kHaRr+dc/MoNq/k5pk8UAtq1W86XAtsLSsHpLWK58AwKNDJKO3txX
80SDm++vdYy9OLnV1Kj9sqelV21DVI/GL3PRFOmmQdptGUm3ty7U2gPATorr8+qx
SFSyptfsjRU5HjmkLlvzQl8knoY+Zob9bIzNi5e5+U7eIR3ci8mNWONLldmSyuIv
bpSWG/jVZ4orDCFRWFa/3dX+ziqq02gica49LRAhVjX1rxXBzGXbNsyynO+iOmk2
dMJ11mVFbVt1ICHP+uTvKvtPgZi+vDULzma+NLwSSRQQk/SNfWYIw37jf05L8KLu
DK3rKbGb6ReQ70/rTMYdejYmlOPPbWqJv4YhBAwdB88BNT3aJ+FE3utqW21kQGai
B9lNoIxK+UKkHFy9HSQvEH3a/+2u4MrKzIrDTT7rrnZe8GkogW/LhPo2Vi1KVw8d
9fl0ojDBdYV5H1DdJIE4YLwV4o/4QzxjnI8SJ/AJKKgEt2++2UvMxpIZ6+HJLKLM
y58+cMnAztW4bmGPrmiX8blbZ4bTBxomZ2o00BbD4NKt1E/ICcfkI4n46F2Da47S
qeeopn0O9YPgChUrWRXMz1+3KkSZJueZBXAn/QBXKp4G33pPisxVjv1tJuy781rc
OVmFdPRviC2KbHUbHoOXSx1y+O+ti99Z1WooYbpn3tf59xW5p2mUv8Al6llvGC8q
j/YR0Ro+4RDdhCf2sa7sCG6nULpdCxp8lwZV4ALamHoX3tOTOa0BOolhOelcITVs
dupfaKwTziR81o0gFmKj/aMydaaXLEaqu+pUR1XhomScs0eCCSR67pWHTogaM4e0
DmalgHXZw4TojZWzvCcpcH+9CTNZcXqGGMhJ8YZGZGInYIxouEUX5BrvR1Iapaoh
1sRkXCdU4K+F4YxkODhJrRTmWqyfFj0nLNpM146I18FEkURRNfyESfWJJT3wgGQ/
2G3WXA7ne24er7CSBul3uEQL1kwnQTIuKPNUKbS0Zj5v9522Oos8J/eHPJ51Cj54
J13/V6puUQkuANaIRvoNYvuR1ZF/dS+y6IdKGQNEKTGKapXfS6Hrjqaa8wjdydcx
b2/K6597nKjb9kBSZO2xKFjD505ONoaYIlPAsHJ/qfZidHWGj+Z+A75Q78fqHvx/
nZ1C4cq6xTPZUar0sQuKdULBtepu1HVAOj3b4N6pz4N/uFttxCI1jzmsj+Os78wn
8O8z3+tnL0And89zZnB7pA7PHD5ey+v++lMPpv9kXCKAlh2AJ0xiJFLdLuUHoFCd
VLFwIc8R35UOWZnf6aCyA6wGiuYzbkoRE9HtokyBYUawb4E/eqojDyLG3DIbkfOE
BXzpFpeBF2aymRffqTfGfg+3F6Nef/AF8ywI7uPxVOovPtrBk1qJVHIvx8andNZN
AraPF02Q+Ate5bEHF46hw4ptFUnxIL8pKlNOVmg9SaZCA166lEbQlIQsd8pX7Fw4
j8G3Fur4B9iKkBzYGm1kH3OfMDeDNU/q3SulVFUJm6dfrna+t6ZaSWYYgwH1FXlK
NUkDq/N7K2flrK+ZPSa9MBdhMF4U0wjyoEUjIjapjfM5F5VO5ORUHhAO7cCIlMrT
8sp5WgiKjt9laLit4GeiIwyHOF4RRpLFU1DYMT90avjHsmpiu3hAzt7LomBSaB04
8EOZ6+OkwQnwmU+cuZOMzTWwU0IFpIGbdnMEwUiewzawd2j9Sox4L+byaWE4RYeo
m4EmZ7LntPYnSfvNvZVEfyu9rM9IQJEF6PpwKGucrRoDywBgFgViEl6g6JnmRJju
vIZB2JF4h9D8ve6KhrTqGu9XiokjQ79gSZla2tjSJ47BUWWppI2pRi2Uw7uGXJy9
UjxOXbxJAvjCDFwNiSsb3ZoW8ADC5xnulRkER1fR3Xk+Sa0dEHVAUxOJ8OVT02m9
3Z/dFTDUpk2SdDZkb1flIHtHYVJi7xrDWymWq97JURmPlYD6CaCYLVwvTMI5RHW4
kNw/7d+0J7kzQTdBo/RF3XOxcSGhWWcyzKFtr9b7kq2rtSZ4/vsv9ZzkzTdoxz2l
/KsvUgkDjI/SRYZvK5OHur9v47rT4Q8TRoDIFetJjMRB8e7D6MQkKxU6jaBYDdpb
PcxVRa9Di81b9CS23lL5XQfO2++BwS0Q6T5s7xffHAnA4FSEF+uwboJ2MxObq0u0
xtp3QRrwa0tkDnPyTgW0bxj+Z1zMbz6AwZX/8fEwgaQws4ZmGvF2Yl8O7EW4kzR5
1zDxLmhZPpGarJhOrQiqr32UW6Qjy29+j4kX7jOykVYUsCDGiSsVb85mal6Fbdfz
rAnRlu4mbzYtz1W5vpy2J6nUyyf2DUm/RV8rD4RM+a7/wWjV8HTzeD9W/jJcq/Yk
wFDMEgi/NwjASUhp0EHV+QXNLVrtMrJGwSEUG6hb5ET1/nenJWkAbPsWx4IlcAhP
tzurih60axWQWZLzlZYAw56OkhgpKtuZIOTSvQEd3tc6Lkp2KFinjy4PRRCnDO04
nbm7sj4DFB8ogNyyM49mU6kQsgv2v+jPaq1yvhdAnnRCWoeKS7poXQ/OZuUmnDMD
P67M/jsHr0+Jy5KWCRjZfqblSFWx+98eYl3Yr368wD2+0HEPh89VV4UrLl43BjCO
phoHsGWo5ZwoWElok2ZfxCpaDWhz6u/56/AymlFlM28xkG05MO5yMD50uQlw/gtC
tCNClzoGAliVQshURwF8AyRYjgsLDsWINq9hm2NlauDhssbOpI2I4gMgW5hnFU6/
QAv0+9Y5gJtVrByQjNWp+sbpE0n86BpRvOecfp2mnqEKxvwubNETK9M7DfCOruK3
gtmDxVDwngSb7eH8tkDV5yzi4umFvAe+OpCrb/w/pFliQcmTKcyP0xfdIlXnyVIo
htuyATa+FsfSukZ01stHAho68Rs3Xj4rbVi02gMJPxgevwQtrn9H471zPWrhZZ63
Da+lgUKC1EMBTdtEZg0fIKDiiHO2G2rv5ZzC5U387tbUJBkfY3j5lx5QjMzMBIZP
nySlLz2jpXy6/00JiXyn1rYTFllokbHUln26e4yykpmCeNan4eLPnr9lIxCzB6Ip
mUNHo6rStyj9Xjj3VFr6EHG1RymDBewFSyDAUwgD/cN0k80mioS2iLAxqpQPmuwG
wYLfixawjmBgntxHkicYRhJen52SIKhHMVsUexi4ku2OZHQEmeIHOrJf7jKKjdGJ
/969Px7aS6LRfdqzhOim9cFQiO+vbJSMFhX/IL+U4+QJlkHm3XK5hyAtIXWT4+I9
LUzPFUo2X11Z5F86Ijs67lAlehtkn03yWpNxtO080tio+CyLp1mDl35AZIj+/0B/
vBleH2NeEWdiNANiVxPMjgQ0vLAnX40Khwi/aeoTAKC6/WigweX7/jPIrfN+XtQT
TSHpSpwWnt1WKmBpaS8lEKHZeGLqF8AwqTbeC6b8CtB0cnvhso7Snflh3DAbzAuy
sicZGuzaDp2bkc7wMuX59WbNgoBkzzfUCqzLTMS4/bO18QMSsSpZiALwzKUXbHfO
ewMyEeI2k6S9U53kJumoOrG9nvpCGPHnoklEO+Nc7mWtoxufb3CNSdN0gK+6Iki2
8rFUCjFyOFyc5GY1rqxgkPDKxzAWwkTZFBRhxoj7oabfkdstw8/kwG2l0BxIiSII
OXckBBdwyskdQZYLTju5f7IWTvZz4UxZaKiBM+Xwk2q9IP5SLaA6ZJ6DTgB/ZlSS
I+MLXFAbecDyIAQ1IUR8wfeGEVSwewDJvSLwZNUtfZZALF0YyL/b+nlALIAhIx7N
/WYBZZfkofNDZwVSuyRKIgy45qJupfDOFFx3nAjUX9lXSDYZ6kRwq9vdKOvb3gY3
yrOwNVTmG1xP8p9i1Lm/6Kzc5p1z9ssJbcwc+6jiARvyJf+FSYy3R01mK6Imgrl+
NtWpLSgbf0NV2hj0MsQinmhOgCKLK7fH/tTT106FKddQRES0jq58BqQ8KVasonso
ZyB21LYQjM/uMylJBzQVOJUrMwzos6RDiK9wbi5vPIhDFvtgwsa2SW8FRAloOJVP
kb13lEdVpLwbdkORMJCVdcdr0bn3Y0BAqBUA/Cyo+wyAQd04ZSDgbCXwXLu93Fk0
KL482SVRiDBPF7eaFR1yAbJxTIVbP2J8QCL6QahSYwI7VuP/EFACEQNYmrOxh1KP
FbtWpwHPfktwJymjbPe9wUQXV4yrhuJu6wB7NF7qz2b+R9KJDMQtjkggrhie0SqY
WtoznoFMeZHf+hlrwH8kTjqQfXRz5AfgX3n8m9T0IV97rXwKh3NenCk0BP6ePTGy
dS7rpUqSOw7icBaYd0d0JuPQRWfLyupW04C69fjWaqBy9K63tZ6b6yFiUXaaaAMY
1XUTQshIAJjliH1NjgBet1aPSM5W6C2YJADlERADBhqn4io3mkQXMZ4qllRw840N
dGvg8RvJbhXMzZOp4m+t5ZBngUSN6VT/onddAUXofh62XTeDFbXjcohydEdyj61r
x9m3I5xK1pGuv1Gjcmee6W04sDGRWBQW+kGUhEWjNhm6WDPNAx1zpSzWF67rwikp
DiyxAClrSw53ZRo4nu34LD4lpIiN2K2Y3/g7SnNhJ7+PKiQG9jWg4mLbuz0HZItd
DY9r/r6Zts1JM8fBF70ILGNL/XqCu+O1jVRR38ziCNlxEqMsCMuBygCABB2BSFhr
Q2i7jPAi10d56MzPoQCNP2oUydKxoC3oke7uFIJPHszq6eybRRE3kD0MQeDD93du
iooFgDVyO8vTQPjtbbbC2g2+8E5uG3sjMdyHSsGbmpQgnGI4FdzQOtnPNaMdziWg
L6NKGxVhfvFn4RHf+nYTzohKc2dM6BI7l5X+DeXGBsrd3EjR/aOOjLpVYB2j7Aq3
TRGQOOelAH1HaIeVrFzGbzJAGsI8f5eq2GycadIhPMl4GDeeqi8nVbzt+vfNun1k
aWuBlabAbzQ+6al+W6x16kvoQ27VG9z5xCddj7wFykDxRJ23pZayUxNaFP18N5gM
6x8c1jUmoFG3mVzD6wAv+P33ASmveFWZ9A4At0+4bkzXteyEkZ9zpfQVGUzAeIfy
H2lgY/EC2LTM10aWYTM7VxSfirLSzmBl6233AA+JdhdKIIb4PnEWZy1wB2G9AX8A
OaTpEcsNzw1jyxJVftYl96z2dElh5TqXrVZo22gxq/g5+L0JjeJkyxwBRnkGTgh6
gkWmlAzNBEMkv1y4hZa/fMRffCPdiNUOie+C1Pkkgq3LwplOQ17Q3htSclBiTr48
BoEFepXJ3NNgh/GD94C4zx40N73kAiv33tLoIH11dVHi4ztvoHufr2qsq3rb20Xj
EFXjADaQ+p9j5FljYeZKWRwTsVMQtV3cE5zPznpPv46bVFnD7bN+Pprl1zbTWzkk
hare/sCQTXqhoJmWgQUTOkPAvc15NOpkAw0BcLH9rAEnk7yPeGwwIFMzlFRLIpC5
A2quEzrMBt9ILwo/9O2y1xcWDDcBirUkDVouY02WmiFvGQY1sVMccYTwVrC4NCMj
vcH5anl3eG9j7ILh2PniEyO4zOYwtg3tZ9M1WfRWnF3M+KeO6lOGrUihyGzkBqOU
WA5vmrcz+HPCY41TvOo+TZ8MrxHfbnuq4tX4uE22Hrisu4OpImBKkukdYITTa/ti
4gJOiwPxWhTSOtu8iP7hBPZQAvVmXLBVZU25LNiZ3ZmDJriFDVQWzclEB3bZ6bTi
c6uv5fUmTROCJFGn04BX0W6IJ2mzu93aCPhBi6++MgbK8B8BGEXzAFFliRgKc2Vg
/ARjboEXasJxOKr0KQoCZpPZB3Eg4naWlQ33g5/YgTWQw3auCcUR1Rar8FNSNr7F
ipGFpJUkUBjYFJUjEwuIP1+3M3eNfU9hATXtaXoy+axipA5RgTtBacbXjuD8N8c4
q5Q78J2tbOxfPL75yYHrNSJ3fPbh8mkk6P7BjHjcbmr7GA49jhNZUkuwhgDXaYgq
grB083jKisW9rxFiT7mbJeZ0Xt5tCqyFKVP2SYmMYTytgLz+wP8QfSkfZUc8jBdE
rWs69Vn+oKE3iU4Q4i1f6LXgdjF8dy5NigJKWvWcAeDBwVyzJfM9sX5U+yNGfYRG
3SwlFsbVTfTpfeHVWmjKO5YBA3VL9JW50Tv6uUVxzjpbbiHgNtzdVKfZTT6ZSGDt
1tRS4PszGiSZpdNHptcX6OTDEILged75oyyDLT5TNUKTuw0CVKjlngtuqBw5fEiT
NGiueqbWVKyiZUoGI3ydZV5Cuxxf6G7ztnRcOwH5SW7r9J+QK3n515NN/y83a7tL
nVgb/9A1R6z8rfMTtWfE84/A8bjL+eG2ShCpBzVT13zyJ+8PN4brmkn49RLfx/2m
SV+LAxKqw+qnXyv53DDmvOdO9p4h6w9wU9Ri6+IUzQTJY2GW5vN4XXdnD05L5BLI
+zTZ7ke/aq+260NnvPFLucWZjD2u1ulu49ficJyDZ5+NHcu7x5eNXafZqAuGy4hH
O9HiTeZrhHnk5aHUfwQMUmIUyb0UP1c3JKsx3kypqW4ENHIhBtibfHWzTiLnwAUL
mmdh+gS9bpkQHyzEPSJ9SxKkFIsz16aaWjkownYtuehI8tJ1Y8gEFb5Ot7ze+x7q
7xI1XSo00fHq7je2TwsFH60/gCWR/nsTPYqX7SZOvNm1SSujkQS3DUhAc53ZVY4F
MEtn5syjS1Rqd6QPbcaMuYiSlCsDhV98h/BdPB5VQRQKvF+RIyymz+76y1HogmMI
DOtInW1NVUkKGKVysL5pQXZEKSJAM8+RdX6HRnEDFnux33VWRY5sL4Uxrp7ZV1eh
OviAqnDWNQ0yPCYyboN1vz3PcUg0cTNlPYvYOTLZz0e5XcNjzP/Ek3TbhbZJRaCD
uXBKFKKasU1fx35PkBDOnjLUcFPuewPF/UiVL9ibH0C7SOeWLezvetpH/1v/l6of
xBtLBRTfcftqC1Pr4NW0OWuMXyBpgTg1BGFSf5kuq03M3BXh4M73iSXETDTMoCvi
GSjkO4kB6MaQvYDhl3HUWPRzvOrguHqK00Uj10nMbhtB7reC4NkidkBpbhpThuQa
o3G4FA199yf/e/eiDR8R09kv+yfXf8ghG1dUZdfGRO3nN2809PqaRbDlcO9wtpDc
RhXDeTcnv+RIRD96I0CZowNxfe5y6HZn6su7GvJyRP6YLllpGJBJ/BgSuHVBoHl1
OD3Bz4dd7J+QlGm2ixvmha/aRIMIO9v3WupxXsDScBD4O64FeSvasDrLIIuKH+nA
h4aMWPyrc3as1ohYhnvWOQyI7Gkmc32L8Iycl5EeOn/kmfsD7B4yelxHjdoSDWUV
0MIjpZGEAr3Xlkd5UynUA957kXOztMXvyMQ8zr4kkRSkHZn4W3YPpPrGuNhMjuzK
E9VL2aS7WNFBdru6hIbFdDIomP1q5V8SiJvng41O6SnbDWVd6IU0z/HIaLQvf8zb
UdQm7jmi5/bCOcD8YBI+p2DM77SVKy/fXohI6NVhzansTPOqdSk5gsLG05abhBWY
sGyVSy7HaL9j0+OIG2AshJPSUsHpMQFe2vXATc5frSEV8IG6V+cyuzyYiXtOBZet
45n51RxJ9HPXc3cMiNpAhqn4CF7KWb/IjUhG7RVZLhQ4JYhjVi9OpWUjq4IXW114
OytO5h4jLbkcmvNLXGaZAI/PayANZ/wSBTFpYZBfrfZ+3MWl5u/UmEb32TXTwerq
hHFr1RzuaK9EUC67eoUtjPkzxteWUGSnBrXr101IHc2SgkZcYZHisoN2PafH/wDq
OK4oZPXx7emx0mZBLfNlozswX6JkZz1UU1eaMi+zV3UR1D+gztFKqlLlwK+ZyYJ4
fXiR0rklvQGcdnx2WV64+3A8ALUGgIuiIdwpyhPvtJo3HwQm3alN0GNQsxgRqmj6
Ignj/jcB9TRuJUWYrZhPGGtTce+t4oeaGvCoc9H9jLDxOsNimeOtNSFExP/T2RM3
xLXdMhdkLZLqKDM6mXO9dmznHa3kjKBBxu8V9GY8RbxR/bnrKzhsUWIE94ZVJCJd
xcI6BhCNKdQuDjTmA+EdVZ7SZC0cSQpN5lOSRZj/LlMZTLpJsnSyS4UOOkk2H9Pr
e1Aw/XqDvlolkDzG0z7YZnpS0l5aW6npNt0iBaprmCxQjeCWcVW9SjDrJnY+/G3f
iIjxXkJh1uNWDaek5ahpTTziPppoEbfyL4SipRvMgJYyLr++7pCe+cnRzP/ISu4F
MKkPQIB/OdiyARwrOJFx/QXX6yCZ9Q5NfACif3THDM7K0tViN+Cgo/zqLlOLWif2
Wo3RDFzgrLOA0xTjLa+EETHY68f11LyaD40pKlQlBwzLEk+Hn7MTBEAC7FRZI8kp
kDUJa2b+cA0fbT1AOMx0FAOJLU4EYnVVpfc8wVCaKLatDgH8BVcjBqh2WSZmHX+Z
DKZ5sb3zyHMXJ1J+lEvWvkI9+Angeii7iG29dVYlAs//xWteZrndrEAtdpxHo2mj
BCxOpjSOPml9zjHS+T4WjJ6eUZjgGM5uSAJp2KomHjDuuG/twFWFst8SZLBe7ZvO
hYNZXXWt/rF8xk/o2DdqPp7py42iVOxB30Q9iJWIwx0XNmYLZPM9G6DEhis6KGF2
LaOmLyM1Ve9iWLctR24uGsEJR+XSgjihEsFy/pZ788QkB1mLDk1+DWBgmUaB8/Jt
CkibN5d7HBAg64RxOs8tLdRbOj6uda3RakB0oG6at7KKanglUuWqP+0WGNH1200p
ADoxu89vXcukCh/pE153jyWz3klwEjJfZCwb4U0c3glYY4lKpxf0QU/qGCdOCXPJ
xg/g3RlWlDCtpjW1hYjkHEUKhd2pnxK78KI7DlCIGJnVqN2RJ6GCxQS2phIOSDrs
hNLN42lcuQuwY1MQ7Fx9Vjqeq6vr4qeGXuWt2pU8FBc78SpwCbXTW4D/rFp+c2P8
E3G8WO62mJ2MYQ2yyyqU6SBbPqwQyQZNsloUXgN99coOQSBMWdXB08F5nxP0fV4+
UkeTt/jWDt+tR8sGrGajlzNM4UpS5CXArVJgHuFjpIuquWRrbnnRCVTlJUddgpzk
g0OViCEPnu1AqCMQdb9QqM7Ez649S7a7nCuTKYgWH2TRyx+XfmQniL6zbwkoiIw9
KZOkbtMsSIQR7E4yH02wFlZoiHWwA0MZWrW99LHq8c7Kqvhfm8T+EQh8z103eH15
Xpv9ZcRhSV2Bxuu10cl/KleoE30LjMb23csokszVV+xQhkGRayO0Sg4ZDLmy5MEA
HmpqBcOd6J8R2uCUJyTlkmNIeRz4L+GeKXQKxd3DB0C1qmgP49TeOsRf9Blc5LzR
pJqM3Gy0ZKbGleGTwcoqaMq4a9F0v6ijS7B8p+M4xOjP1agSIE+RVrlD1xGIdg81
zjV1seH+lRpmF2yqKCBsdafn+h+6UuI9O3J3Nd04VYtIrqoJekTULL365yqLEkPj
G+w+ChppvJ2VfZyZpgd0xZJwMjwNtQD4JUS/8WQNm1Ksj8xmtK6SbdwI3sGOuk9g
2Vmtimi/ncaceksGgRyW4D/7aTZair7ieub8EVFB4+joxBKXjdd0kr+eSNC13crW
7lz806AIt728S2HIQXOrFhwVjW260jlojSZI/sqJinuPa6uxaJJkS7A4XJ1ruT6i
NZ3ARAKnp6bLerqhZlZK7L3fum5EIqa8XxEfx3nPAg9iUNe/tXgkN6yCNsbXQKfB
rOhCFM/yhsi+V4HeXXLcQq2pDBYWaG4F1cqcgpIpELXF/vc0WAWD2EjPraF/CrZ1
EhCsMgy+wjF3ixIywlNYOigFsZG+encfhD9SgLS0O4nnBpwGElGx+V9rnhYO3M8R
WIwb4QGCZsLihV4/8n6n7jQq5I/2LtE3Lej4NkYMV0WC9GWTGf3QIXi05v/Jz8Za
WBq5bXeQHGCDgG0Uo4KlpKjI5a7iZzOa7k5Rq0d6Ld+cagiBhOEj/x9kLN0qpZmr
m4GoWzFXAcOb2ob8rjxMyD5fsFs3ybwpVgrUPZYjrQxUw7T7F/C+MUjLps6INpVD
XADIEBm16ltKVe3MVqEr+8au/p1bCJhSEEdSk9NLSXbtGtK8nEr+KWIy6+OlSMc1
aY329a6nMZY6AZX34ght+h4VwousMF8sPV9gKCqnlmIDA8+B5j5mNbyU/SEYzImv
hUChPAmn3TGXYABpyh3VlbfPUAP0ogLZdNbFETaayY8ytcKIZY6ghpmT3gzUcZAi
x7sLxx34qiLLBA3zW/h6qWvtJYkLuS3+yA6yyTiOtUec0Bym0XXkDjCnBsVi9eX1
Lv90L5yFZZDqDvKGxL2eduqSo8zJGmbHWKmP3/yypYZ9MX6Hfyr/klWXSDTlU/FS
oVw/Lni826MgdAQgC3l4MSXGGDIe6DUdVdnlI7go6wskCj03JAtX7Rp4kLnBLFeU
OvQClecrZAXGvZ4ODH1XzHYfOLVvJNQ6He4EmNWL++0x9TBhE6ruf2waHR0jRQb0
6gt6ZuOvbjzB2udTu9X/pAicBnFFRAAbUDTvCgrVhcmPKkUecyuXrxKOFZ58ZOKs
7nZXsMuBMsTzQ1F+KIScU7rwnw5J1I92P9GYDb1efpQfNRmtG++MRey7ZzEcAEwx
AnlSsoTQcmpfNkhq8GNfXsdE7jjInejXLt3G6qNragNHfJjGWsWAsdD/5AxV7tSr
U+SqG1p4GDQ02NisgDVL3mTzADA3NU8WIwBI9lLgoHoCfopIJU6cmYPeZDx7Q286
gV5nA/YvINqD7tgq1rUGUlAq7DKSK1+CMVX8zkSjsvZXu5HIkJYDfMeGyNtoKTMB
64ggXoq99QKTUbRYNW4HO6LVcGkGrnlQmVYHBqkS7n53SEbKiBDqOBY9qryIt3HP
uDT8zaRsV+zf20faw3NtsAH/75sUHZ5aordqXTJgawHWJLSNtFmgDZzVVY8nzE+K
ywEU3kBriiTqzes04xbySPC/E4uDyI/WQxiN/rvJ91tBzmf3coaOjh0RTUTEYo7/
AZtNc87kNW/gytr+4Y39DZszf0eYEfXWn2XlpPBM64GiyF3NjETjM/T49jcnc6V0
nkJLyrhcQ7hR1QXjNhjvh52LlXKa+Eu9CP1umt/eZRQajnOLQHzaqfqjMScQAwa/
W1YnFp8i+jqq8rZtojzPfr+VQ9gm1jm435p28XJZBkcALMwy18eIIdiQsU6Nhq0p
1dDCFRuOWPvNkmsMddY0a/3Ug/8jX/WwKZ/N1vf4Qf5DmXmdcIabdiKtPpwO/tAr
TNTvZcJbXuZTsdCtW4eanlVzocUXE9p/wg+X4CfVUxefYO5Ct1uq2gvt2QYymYxo
BvwOrVt3wwN4yaA76lKDrP2rTuTB/HPgE3nQdwhag73CIhZRyyDJ17L3GkCrkG1O
cue+Efz2F5LISpG+PiZgicUCQPC0ZORmHhGffhchnoOiFcSl2BBkHJ4QZgPfqGEG
vhyFGKBQ0hSooFgOqmHGC0tamYct1G8X23gE+LbE/VSmVCJvQvVs2G7c2gfmc4qX
ymTgcIiY7YscUP2WIldi8A7CtpVT6p4uZrx19HJ/GhzZzjxPEQDs7q4Yql7Fb4Ag
/u3XDiFui5kn0nrXQ6JbLAIqHFupqHg+SwnhSNY9o0DhCYL7bUPmPF7P1f4GSORZ
tX25KDhQkBhNull39lS7kfXL1blf5FFzZ/OU3VR6AhUlDSt/Pba4GTYHXRv5n6id
CS+64dK8wBH19pmvqpzy71GEoIC7aTjZjt5olr6B01KysYVcDHtSoObDxnoIoMuI
v3LWFwbDOhluYHwDKgKPcfmMPiS2IFIiYWnLr30jdkxJIFVpdQZdLIxV5z5svfPH
plNx7f57OtThodVeBg9/3Xtmm1ypffjISjpHfYaFCvAxrK9qmT9r6T+aeHUrWSU9
QU4LPlZrbMVtxIe1YIkrpwGIVZ1Ktp/P11hflS5ZWwdoTBFijwh0QmRsCcUCJEnk
593rCJm0pP4DsE6jIHGHP2ISVZ8hGm+55Pudsf8MGeNDoJeNBIQSyo8rb04MJk6Y
6wQGQyE525biqNKqv3Yrnnwj+C/9g/Wz0ZuKq+K1XjyXphCeULsNIyyfH1utIyKH
OmcfAKsyvqojgvaNivSdSHS/e7E5b5gioaPu+6zjVEqztDpSL/V0yBO7ndFukwil
XTXkzijB6MuijKmAtBn2WcqSvjEHKccEybn7p1zFmkMz37kZLMyUnDifcyxFibFQ
lBmyn2kmCkfE29/4mSzMZsWrWBs8l4/b5kyJ4X8bCO6YSeX4ZgU8Q5wg4nybBgMC
+dd89SX9jClVUr7/2wevHxU42VxAIu8POJ+K97ohZgIhpgVM3jTzlyqkxUF0X6iO
fz/yC5RwRy0EqIuZOKakq33ahAIWIL4MDKwtauK8kWTEdUpcEvud9FM4dA9m2dKj
2GRqvrBCjA8yDQFIWc3B9AiOjlyA8VDV1d7Oxt1nmyr4ofUPYiM/e6CjYyTzqact
Yj8sZdL1OUFg4U2ScYmD5dhBtfIfZqlBoWXh+OH6J/u9h00s7Ke/cYBMrGBGnknB
CJ/ptwAcan8rXrASLlwoIn5B3lsTc1OQXNzckY2Jh8pUvg2x1s1M61BtNmtS6lne
GSQjaoZBqa52oF4DjFEkEDqbBfecMZZ26XzEJgh4LV5Sq56naLXa2OFHS4d9FeHf
8uSj8nB6ALgHdf2/D/swIJpcP57aIW3uKVPWV9waIMXt8lit9t+HhfKuRteH3mSI
4oOFoRUiQuHHEK2xPBeo5b6LI2FFU7ZUUkvM9754vDX6W87GDdSPEX5n+b/9yQ5i
UoZnoTZRAGiaT9rsKxTaI5oJp8B3lOgqXN9hY34r96kK8l6GyyW8dFlo4pMe072f
4LjC/o6cvDsy2jyBCka8vTYizSTznfULDUHjX0N6G1U8B3NsDj7lUA9EgpoJX4D4
x5fCn2llZ+cxCSnYipihaDrL8hZrvL78l06XxdHdUEgbYskVp4xW4fqRR9gfJHaq
msgpuJo+evfB2pQhcVJLD/oCZ53BI3n0RW/d1zdKUFOjPMEX3Sfu4QCb6UOr+QX2
6HiCcPd46cGC+Xocsec2wHzv/AaAiXjxHJKcXfh6aASIW/KLinxqdZPP9/Aow6IY
HFO/YkqEA6H913A6nu2QdbZ7nUvED0FhB2FbG7Z4W23b0gf7LN45kIBrv0p85bDA
nL8dhDLlcCPYLClI2rWW9JV7m4jfBJQ7OjaYMMTyErNHxqEOi9X1A6Jiu5a7B6fw
XGneqm+TUovtTMVmm+zRenZX0cE5Va1Yv9tfq4lCi9CTle4gnN2b2Sj6FrTq11JH
K+oSW2LsiNKj9YptNNcAdYy4xfdhjSLgEgZI6gjFBwIW86azgEse5Eq+H5snQf+S
jYogHdotmONNwdpKachP16dTYSOuQEhK23XhtvGVGmCusDhX2g4f5b95VWtzHQ5S
j9B8czDxLyOBC6XFBWFPYcnYaIYojvlKlvQH/l3lIHnMg6IZzyxDV/aKcqxYv0UB
lemHNaFvVaJ6a1CcJP6gDOWVjcYFUjhS5LCTbcDx2fTGDJFBKYGwSIkiOsGwA31w
1umAUv/SPYgFRGFD/CTdm1s5/YEUJUgILJ+f4xx/gnZW8It5vcpaLhnKSXjstrvC
pm7x2QheQSMKKCKK7QynBPm3vphaIGCJrLYyxhvYXb5ubPG8DoF/Xz8jLxcsenNu
N7NOLqQZlZTkYT13GCHEoUs552yQ75bW5YXYglCSG1ap9Lc5c+h9iJck5IKSVxG1
psz1+Ccrhrm2D4wlGXoPP0BQ5Wmk6LymY6nXLcclBiS/a4iNQWpr6utK5kTtGkd5
x8VTE97Rg23MxjflutsHw8q0d2LodYuF7Jl7+AjGWOWDo0q+hLNvTOq2/JgnfV97
gvRQlBS2BeAGdlw6r+u6uu3G4KdIxmXv/RuYcUWahPvAcoRppAe49g0becTBPl2G
Ll6/uRBfYx5y1NBLSNKWE5GwwYQbjCvxW+wqaXhvZD3oCE3SEpszI89G1FUdJ0B/
iL0aSQuhijMQ4qxtFMZuEWAZLNhY6nXchbtNGOJUSbVJNnGl/A3/mDecwnkTp8X6
2+W+7c0XDW+djZp7XGXCbu1vej5TrDfGWndRHJL0pQ+lDJX6Fobz9kT63B1A6elz
oxc7OyZrUiPnGzqQ68AZH6YEhraMpKohAAxoyLE1kxtnXZb9h9roh1vIRaYzV6qz
zI1S0ITmZTRP8i/+WJRqtBWBkzcaSL5CgtnR2kD7BYyJAOhzg3vq+O1mBnx0eKGc
Fl/FNIUQcmG4kvxXbeqyfFaYdKECrIcUxU2R3KwoeDv82Sp+XdMyqEwUqewiU7LN
RU7Lb1T3kutH9BogShPjMnnVq62V/G/o7/nwmZirg/e9L1S0u5sKDsrhDuoUOMi5
avKeWwO/hYSTjelAZX4wY4WWzckYKF4QVgsXzx2bgNIuO0ewyYvpb8oxDd3TkLo/
MMzDbf1e1gfMtcc8m7rJ9oTTKqYOqLU86Cbn2zK8x5wYPXpfbjOYyJ45cfvXOYMK
mrMuJOfL1Z36ysMtqagtAIjPAvOBpECyKjm/EwLgKZFDwviPPpYrAPrf74XxMKP2
NGl0e1UhntuO02/3d/xUbGjbFs9IBLei91posx3B3B/7ycJt7nx+Hbvy4s9zW6nP
0geqgQ53k+MMlsh3Xttgo1XlUMsgwwo/x+7XspdEgmU6jex2QGGQp4v8ZXiM5OlG
IdqOZRi4jSa5T67lM6i3kAyALBRHLwAOXm/LvUvYLl7qXK1IqE4eyZqCBt+6UVLQ
qhuGGlauPJW93G8IwPr26EKPQw+OC6k/X5qWEdJdRVu91pPtp7NmigK8EIQeX6hM
Nn6GMhQbLXth7fcASFhU/o9m2unVKb6DkJySW/sQFUCIo2464zB1AQITB3rZ954M
I3aPQG88XJ/GVT/iDFY+P6AAqBdxMm2ru1QAVnDS52Eds4lR6kPEZkINUzh4lMjj
hfN0LA/A8OXvfMO4DJtqpSje6ZKMIhJK5dAME1gh8b7suVVgs8H5wJp0z0f9gofV
aFfDFg7qCpSXUIdeuEApw3KWDLSIrs57Z5cb4MKIA75U9ZFklpsItDz0ic5FUnON
axzGTbPbw0jOZKJupFLL9a424zrKjvTbf/y0xIzRJMEtfY5l+2XUdobchF3/+WIT
JiyIG1IbmpQVtWL7RO4eEMnEwyQSCmU2KMubQ0JbLEbFxJ45GQ2WIcPkVhHj3fMa
E9X1bSYM/d4pBj3UN7Qgpl/GEKVDipDGEFEtPPV7snZ/crBOKZGfkdIVgLFdfGNr
QmW5NRwMFyS226v4tF9G8QqqOUSAwEzvLQR5qhX+l6DVaMC9C2YrSo0bLAxkw964
wdnXQyojP6qkCB6+KPhQt2RPkXCbk1w4Xvl/7dS4xrh2C7JTJuwCFrgZ7b0pg0eX
o7Cvi+VGsNIns5vq7c4DDp4lsANg+nuvT6sMyw16pPGrR+HpLtBF7jicpI1L0+Ds
dY0nwD+Q4g2kmiYSS1YS46hwKipl8mJL48U4tiEBWqJas8KX/XYb3a2Sgz/5Eff1
OAEJEkhElvBMpkO/RPzc19tVzp68GJrf63O0E7ypdyRL3Iob9VtdOKgAchF/iXXU
HvpwaAURPFCDk+71yyMLi17GrXwSKLMvQebldQTRBkVMtMGCk//DjM+juos9SQdY
3MfJPxudRhdpXVGLmxT1Cb0LB2AffIvRg42MBsufGwRp723+sLtIpJvOhjeoMr+C
1j2iqM98wWkiLVKra9SxjDe+N3vuiXuxrr2RLyHV/zTj7XF2MGsHvHjFmKb3hpB4
1R3N4HUdHPH1rx7xQr1RnaTptWWFhNb2C2Ld107AALnZPPoH5p0mmKskODHkuN3X
ZKaMBFpajuEBFfcyM2deAcsNMrM81QyUDgOn4i4MClJwZ165inBEIzZ6v2/yquC4
vCEbk5lmgXU7AuQw1G+xkOU8zeqf0FMHKM9go5vyozC3tSa/rrtbMkQuzI71ybR9
X8kcnpLJB+09kxVGASzcZfbxnvBFfrcYZm3eSVwOxDlYq+29IpXg8dTJ2RwQ1/Q4
8ioKvAW5jAPFf+6IPj4mPtitvtEwk7E1qs+CT0PHS+n5Ipg6pQ8DdSKOAHYQtRud
KGcSJK6ZLSugjwV7w7y1KmtDnuHJeGmUIBcHgRWDMv3rQ2vZVkV+Y5pGQOBCV7Ez
s5//1aYKGNVRogTOm7MPfCBIrFVj2BPFq9ZeUOqg0LnYA6bLFzEfHbwemRBpBjbi
cJ5QfnITIuItBTWcvaX8G1Nrz1EtVWAKeakMY9HAk3HQwP03HzsDUylbIArelCEz
7QxkwTL3ibzaUmbZvvoT3+/9Gs0iSwYbRw5qKpFPspHwbVtN4aETThRU6ELUQcd8
A8S0nvhs/2cEg6xRMp9EYRvwLi2mdzMP1UPzQgNOHBiqEjYMg2ZbI6fBjcR508RT
h1qh34QUJTqsy26AC4RpPyogvj1cMIHmOhegNCdPxqPKmTP+a2nezGAxMCEE16Mk
PThZikCeqwG8Petfb9TotjWuuJCXL8vn6Wll4wGZJSUvIDUsNWCOUZKoh33vtz/U
Z5pW+P7hkiIhpqp0XzsRy++5EQPqmburwZUvG0Oof3RSW2ai6oJu598evRM1d5re
pcwWyfEqOA6Rlxi2SbPoYBIWVTA3A14WRsJLQJPGToqyl2KvH0St8VLRoSv0Li+m
jSw44jCGfTvmU7n4NN1dhINyMdBHU3onBqZPz4e/gZfbq1Y3dnx534VkWO3oxWlX
Nl0INohJXK+zQj/AMxzCTxapcnZLQrz1vzD3fKmHAfsaknkrgevi/Fwjg8qhyIWm
pky+VarmjbuN/nQZTMhuUsJBy4ucwkJ9BynZ29/JbrHrc9z+LffUQNbjj1SxZP63
Vwc6uf5ikOE5Bwzi0ES5we0oBIqKoHGx4UnYtmqWRjJ/G2TJW96VpEQsJdyXOf0s
DatU49gJNWidMwGqQMN5nfnj92Hw3Fi2IpCjvLl+VtJweVGKXxzKZpCSAgA04xZG
fngWUskgP8ZHIGSFuniDWS7KlWR4FdRWC5c7ZHYdvMTNQAPBIqUVHtcWhcJwrzIq
hxV1ZNx0hdz2nMcMSRXpzLvbcWFyaJxFyPh180ZhP0M5JPnBSOLm/bxN86TiTQ9X
FwJSirkAV22HcfgdFWbxftZERIa/fFKlVKYOdfODO8EYZ+1ClzDbhRhNi2fbMV0W
x2X+eL2TtjOtI3jEgc/b6cITxwki40Zziu0nlbsT3z+oQkb4QhZ7U5fxHWRz019T
2z/ktI784jkXfBTZEbRWAA0TPJXp5JL8SIfSBGS3AYUVLFb08PgiWebyJ7MYwCUJ
ooUITINrp34nkLFTlC+gzEvZuJElY+HWbvOUqhHgu4WZzde93SDakA9OpfwPmpdP
LVUrjZ8I3/qTb9qbFU9qL8EqvKPgOsNNFOoPctFnHSKoiSKcl0Lt66uIjR5twCAW
vBg+xGkZUevcrkoMNkpv6IgtKFWy5FVrE6j2NO6EMV2mQlSaTVnCmYqeMviomBrs
8WZfn+dnwJU2uTbWcWcidjblB5UhOac5kumTpNSAn8unNNor/n3hlTtmCvvWYwBS
ZIzF/0/pr0kjrjlOsVrHH1HSNe6WWlmT7IbbTBYAVH2ei4vPCrtXq6IyJ+kMMYlb
C+XOmupk/dZk64XAept3UuDJpF9SCmUVXwXGCIYAK2858ZOHKzFbuSmVXtUP7quG
pgKlj7h53cNigCkz9RIFpvhSS0hslHg2Z/1Z8pkddBoGDToGCBJCQv834m2C+XnP
YMRc2BsHM3QltBIeQdQ5mXK436NafrcNudY1zcQ+NFC/9fpMX6KdoKogkASfyI6L
S2XEMhahy8w5wf1QpiZdH53UGgqS5efnPsvwI1u3+4uBQKxs9D/ze6TibN2hNsLU
5vPhp6G5nOztmqE1VPN37mDHMrYYhTJEXxKMiA/6aEqUoA3uJuo3/FXvGbb4VXM/
7Aat5NfropJs39Q91Zl8H9tR5VuDrMesWprxF97ZqadF+eSYRJSvfHxs3YZA2wGR
ydUUfJA0MnF6jJJpkrsc0M1FZ0+ARPsdf4hQ0e9StxC0yDZm0g9GRG58cyRTqBf9
XwPFzshGxePAqA6hrmnNIBcunwbx9lSrPv+JBmMOEE4Wb+BQgk0T2ZMRfP2TdkB2
9EnazEN6JKJkf+x3a/MuJUxg8a5mqdajIyPjOwLKVXvqYn4j9fhSQCHi4T8ML2ew
1YdezVbYjS5H3mmFMccql9K8M5lSWf5s0oe7rX5yd+cAFUe9QI9zVyWsVYB4lylm
o2gfK+VIH2yi1++VI1aGXzEizcBSVWA6UAzvVRUC3SS8fYC23PxCeVICCpZomN9Q
CdpueZO2eQ4tvJxP6hMkpGGOXp5DmWf81jKCW/sCz86nIGN41C+JWIPE/Mk/BXGi
FGuph7UxNelnhNIEzNUWe4t+Zdrfra31AHTIyAxvbhpcqvi9boW7inj1Lp9IyNjD
V+St+RBI/O7s1kJYuMyUAOAC/GvXuSbSicRl4b5FLkuZQjmXRdgKkoN53YYihyXw
ET5GdIkDHehyTFh0hb94Efnq0SUDxXZXLPBWku37QBIT5TgSak5nYWNF7hQuqwiD
CE7SolMWBOMvxycIGcqxwotZ8T3onvafM8qVvTSusV3Ur4NUimkZv2xxVTCuIYLK
CXtMJpJ9gFfg9KwCDJs99TGubXd0Ij0mLxwWUNBuBP7YnfOHhglO1iTPyQJ2SnYl
L8vLQXMlxxMRX2TNKH0rIxwa+WgutV61OwvItMsw6qpv3BrqnveUZTxdPDpfppW/
8hN/zEE9RgF4OlgiRg/VPYoqTSDS+LpbiPGppBay2ugKaHbisVl2gyofp3E5VZy2
vvuYMLLq2rXZ/e8NNdT2qfwXTuxWd87++NbsWKP7ujOVN9dFkCddvru0QwtD3Ncl
xZaqvYJVZ1Tx0xTVRuiKzqXLrcvBGjLbnIkjkcNk46DITK9tUQrXofetiPS9KAxX
1XUY2SNVAVXE9HR8gGr+6IlfHpIZDxcpWDuX8XmBmfwzB3sd0Fxj7GTTvEkGLXAO
j9jcKbrsRhYliYn4Yc59/CB+d7LdeaTjCvrLkMenQtje0Sk18bX5ZIp/xrnUwxo4
6yRnmSCoOCYbSRCUeuy7dFdzXAPwIL/HpR5gBC+nC1JMXugKJ6L/iGC0RlrCVEZo
cVAKS/YCLBr4Y80sMUnXP8NQQqr6cK/qdgTjqeUIDZz/g1ejxePWxotbz3nrVxKZ
RgT0c3lW1u/mEiQsFt23/mfhFLbzHWlkkn0osXw1CHHMFXRuHFzPc0LFB4shCw5U
oUfQenCLY6QNVZNdhoxuGwztiOXtBHVVziJzovZCyXzCWYaaBYSlKGIPkD2Xwv3m
CfWsZF4B3yAjq8ElrmWiUFuSe8zATAvt6m76+vrOHkLjRO4lM1Pge4eWyHPno3sB
rOeZz+MtBdwcmnFKMbkcYELehdDu8zh9cfr99N7kCDn3MZRl+40LbU0zvMV6zAK/
YAxTxQGkSiPqVMn6WXALC0TXHXkrFBBtLiJHxW9tooP/4KvRDsZNlIKCZH4SrVNI
SPMmUUthbq+S3kf6GKpMuK+xWPyE0ao9yEKh956zDEZ8d7z4AQ1zN5bcl2nbyOEN
IaLTYhcH8wwyoVKf+tpQrvfQeN8nAQ0ohIbsGvcApd/BhelJLFmRhfoAUKCQldCH
UtQpUi5RFhDI9x7yduiBycLmpMWsFiPeHPmvP4MIOhUBXYFUsfbpzbhZPJ9wmf+o
XK2wZm7vPxubDEDITE2BcSMdJnkZ6X/Z82p0fU5xxHxNtnSFqJuk5QqOkEvAXg5l
hcGKsj4CPX13ucfHpP2VqcJb+lSvnfAF9nVIJR1VxkxjPnBcuuQnqsAsrYfgE1CH
ikJeur+wfc25PKQvKJrQ1I6QFy2mxiP68aZw99NTAQYDejbrSo9LzyYaC+NQY78c
LLR0Zof/CgVHRPxb2VQXIW2WaSl+PgeYX4gN4Y9hL4cw5EiBaL7zV/F05J0qCfSo
Zw3C3AiuEARLxjdgfIppNHbLbpV9wLVwImKoi2cUuu2I95MygjoqrrYFf3GlGWVx
ATsn3VOne/61DfENu3OZRojlg5B2GcCF4688VP9bggRNjhPrTGxQt20jomrmebFo
6QcW+xdlarOYknv4B5/zJYQPN3dyb7zM0DerlmY/OPJVuOx2EircegD7D76t7KBk
AgZrpKLhIuVU+FW7/EwrzjaN+zKZwmq8j78K3ICfZTEJjJ9NDFg3scr9Kzr8dZvT
n5LoIc829ca45/haopAw43prwjLi/1Uv+Ow3GSYenVzBjExAx47ks/1D09/b/7u1
9gR8WEP2oZ3FwHrwpgD3G+TCLhu2sg3qtMDyiWoBJ55WcBeH/la7thS8rQIyKrxh
TGwwdiV4U2WAMLcAQjR6dC7kXakxs4X7OZHRm0cAgEwmtSkEmA4YCuGbLD/HKqTe
q69PPf3mqbiVocy7oPj+f5xRBKayVTRZkcLBXNzJn+V1tHBGbQCOuskTDKfyyPAU
ZaqdRdn/jL4CPnIFbi+4Jxss9ksYZbficocmyEZVAaB1UzJpbSAq5XD94NgcBcQ0
tfkAPrTjWkN62WhuhTEXgekATaGIp2oYteu8uC6ltHJ6qNZF9bmWEmX0JwG9V8W6
wyP/E2iAQrb4+ZCI9HqC3V+0mhxNMSI546vlx1Ob8LdfgaNXYmUlsd4a2W7WPuOQ
91of1D4ElUeaV/bRk7zuvUji7l2osA+mSLae5cfCYlgiVgU3K8EV/UtU+445mSDV
K38kaLy30nPJWcIMMx9qakVdylsyuaWmV604PsOA1V4GBNVvvkN+FU/5XPHlkamy
3NT1aVoGCr68ZKONdJlYke5EoU/J2BKN/X6vqNLa1cMmj2/crswO9pwCSQdzJ355
DLab36cZ0m8f+S9vzdXfDfqmz1W7/E4Db6iJQQlOpnHKcUEbNO3umMxFoyzW4w4e
d8bugdLuB1fCrSzKDUnA8cTYoVqEvYMbleHNQTP+y8TQBVlUBJg5PMbwgP4tpZSG
y0YFK4qvcOOWyAGfdwhgXu4tgwMOG6iBv+9EkeamJnTj2NRNy1GFFW+5EC5uJ10p
0eUR60ogPw7PMSjm34ewU+wEMtTjD9Z3ujMx0/QYmfp/sV1ZFZ07zRIEeDXG15SC
OS9+MSaa1UMfNx1CTQ6u1JYopay+N6KIGfG/SpdtKA8/wlhDwvB8FLUP/uSD2vgi
z92ZbxxBvKtltS0v0wUso/rKGgRw+5WuowxO9lUFXzvpuIx8Iq+XHVqUkhDo7Ueq
z8z/DK3+qPHyCAzWHZ8RCCai9Qj205gNrsCDEZJeCv3jMiZsTHYZDgikWupNaBmZ
b2vb1OvdSl4dFeNvnkUBcRV2XnB15J3UjpJv4DymB82IGwpzu0OV1pD7r0bVl3WH
F9uKv7yCr/L3L9hVsRa3tg1aUPrOKcwn7STW8Sm8fDUQz2/Wnx6Kaq/C+x2fqCE0
36mBYPjLF9iRUELk4pZZ8Icb+j5/vckMOqblmW9RJBAjHS8Q16HyBt9nJhgMNlma
WsulRwIU5vJ8tJ2QJW81wZ5JhhXKby1AIrxMtK5Z/l9RSktnHnbTdQEfO9eaCA3W
xIgU5Pg0s7uL0iA2dE1j22Vdi8IC8iysf9FBexjQGP8uD1bKUmkbjGM54j1P/psq
Yhzcr1i0iCzdS9rT+n6cIKK+Z8/HNnwo7Wv7J5jYZ4Z0O/yf2rILxBYgPWUxvps6
uQTSyTN7Nv/7VuOaUUch/ml+/B8816J58tqEuQ9+1t2opbL6HbEN8ZmfG8EnpK7w
2rQSXshPIjEWnAxOZUzyAb4LbaMJekCUDpXOMnixKm159VXfYEJxdM/18/KTvGFb
wGYMoWw6UvKim81l6zjAvS+muFoohDopluuEM+hZRlzje9+AqPDg7ggfd2FrYQkE
u5biblaxo5WLuS2DEuO7anz+DMEQCk1dn4V0nzUL/eTLTcNsAIwrtrtkrFg72dS4
7PyE5oXFtCIvl+ZlhhFNovrtNIBbVioqLS9iWr5mN81OYSXvfGpQINP7Zgi7ACsK
Qzj8pUP++gdJjlQHYR66WzEdTCoq3hEaATxvqm/xua3mOTh+Njp0vMBgrn713XX1
tzr2wptOSQkgJJlVbwsle81vFBQ9Lmvzg2mu6EZl+Zvjvh5f9uWTk40Krl6mSFH7
qy1hyaVGaa6kJl17kUeP40D0LxS1Dst0d3byAhYOh4ChWIXFjWoIvJZqxKAunbn0
/9GXQpTp5aKUdReER6qjzCmF9jZPV76q9LQJmuV/T4hmO5otB7QCCIzA3vkZtDA2
s236tzRC8iSBMMjAjCwNVcz0WlWDgBxS/qOMBWCWgBJ658ZZYjVbaAbgapULcAG+
wNdAZFGZtRL9Y7J5EXpBx2b9Mm/HLMUP+0bDzTbWq/HJmPzw2zVTkzkKvvoadun0
GnQY0VvxoJeN1GjAGaErmeB2VcTEPw0gWMRGn+tU7jh1o1OFVZ7XAMeGXvG24Vhs
sbUNG5Bp2sDqO3ip+PaUrb0cWvVZ3z3/cBo7Gxq2U+QlekpIxb1LiHWMfLRNAxvb
P9US/tbEfcO4d/CbgSn08wTA0EXz9Ef78w86eylpyqJ3/tKygB8yuT8g/JBmKgQg
czdCtKVud5IB0vNy3xK9wvJ5FAA1yIe4NQNjJbdkboLFeO4Tz6lEBLW00WoDIbvy
RyuljDzURMug3CtJeEG2EDvxmFkeBTCFxZ7Nh4gLPyTuOvMlGZ30rFurEi9qmxur
nzrFw1duPN4Krt2n3ILu1KvtWarSvbn4jZ1xrZXYsMIDhxF02OlJhKMA6ato6kPi
/EmfxSX4pPRg4KtbgI0vyWM4+DJC4otB6+1Oyhqgpw7YDAZ/95LdvypmpZbakIwI
MaV0AaTW1EUKDOaOrks2AHo+PwjwpLyWehBIArr2l6hVrEZhprqvoh6Ma65AKtNL
MBK/qcYVxyPm6VksgFy2boeJr7xQKwOoyMaJ1+GPquFaY1ogsGzdfRUZ2AozEMi2
ljkodrMedjTrV9kouBmvPfsWRGhy1ExpR7sRAzMTdV4LqEwRQxoSAKlH9X7AK8tD
qwJcu/ypK7AGjjRlhrvVumH+oFS6tzyXqDhZ9I5k8dBdPd6cOaB+X6hJ98QlRmn+
cg2IVZ/GZb8/0lIHwHasWdOIJL5VE6KcQCFpoGdwmRAQjFWpvp82Bgdft+gv8wJQ
CizwJPkwKV6/hnAnoZlrYK6vCfyVuhojHnA/EzKgQI7Zc8bCS3acBjSC8EWx9B0F
Fzox+tf15b0t5HUgrr4VJKyXnWY0phpddWdKgeTHS1byv0YCIpSX4p8rC5q6xalK
6ngtpCg3liugHDApn+FLyMVRpkoxyJhoQZQ+/iCVG0g+KJIVF8hAOeQoWO92hAXL
MGWtVXogTDvPOUwqUCNaKFo9sDDZGxmBJpdgfpTJ625FL3FzO37vOpQZO0yR+Be/
+6E1BheNUmE2Pz90kPfK9a/Dw36IsPWBv/dSxzVwq+i5JQBjqlAAEeCi4a5cEoda
Go5dVVI3C5fid8v9Wpv3LZERrcV/aLDEMCsr5UNnFCvPbK7thtFh/Hl1cfhWnC29
k2ubMPB0mxyWMh5jgC6uDXlM9fsN4k1YnATo47cUWPkIy1utiOXuB22zaoxTlxJn
6FnVTrXUZXHElb5DPnLzrahN23RIYIZo1KhFKthqHM9yMh0iTsLX4D4EAuziqxSz
D+Y6nsF1SdtLTdNPGpZE8fsaeVKBmMXWza8sPbgVfGNy0lj897/92GYSD6TMC7hE
nz7N7aJ1ByjY76nBW+jM2fVl3xBootfO8X3GIQ9YiljgdN4d3tBq9ZX75z8hKli5
MVOmgDoH3irnPj2vRG9Y+VzgXpE84Jw0WuFMRfuIq1Q6j9CfyoBsTSJy1fjuN/pK
wVnqXczei1KH+/+Nf3JUg6/QZLFZnaygjsiQFJB5Jc9fRbm5g9HX8+pDBT/oNdmc
M05ndluGxNxBx1q1VSdXLVzTmmQGWLkBtG28Nc1ygMEL5MkoRJ/nay3+yMH0tkU9
Vpmj1Lms48GaOrGvl0BRJofgN/UoP4uXyCHCdsQk1VljoB3MpIG1n0gjmS8MAw/J
tP40JXrx3R1WWGXev5TZyxDUZjndjGSC515fTCsX3BbT35Gd5IiKPEkWgz8Xx9aw
GSok1JA9c/8HddQH8aZBtkiRv9ObhEbiYh43v3Eptfwv8PitpqzX0noqrFr4eEcn
w7YU2z/YLZSH+SYgQJOq7ur7rz9vCNyttKXcDKVROyhbN3lmRMrjQpdD0luj/vmI
U3HCZwNTxYYy1Gk8dtTGDnidYok6L+0XdWKtcAJHCFyBhKoGcZZErhBziJbYI93c
egtWSE70guyzQpatkv8VZu8aqIFevqcNW/xbg6F0++y5rIiUm5pC7Vd+lzcO9qLC
14uYI1EMC7+mnJxzPcGGh2ocXlp9tZifUenVjDSQ9dVT1MsILVJwyWFOUsoyAfrH
L6/9NxfYpO8huRmzqEmXyprXdegi7p41lDcHYpstISLyahpr1J9gpQJ1Uv488Nt7
+e9+IEXmJ/jftRspACNW5P09J3SCV6a9bXie+j9vg4Rw3C05c9gXe4rM7qLWDzU0
fpycQkfYtf0gmWkah58aMLk49BAd5eLypo/9pgYkugwWnVPQy9bHS8bCoxnhG67Y
gB0nuwbpqU/yam22FRCIX9CClG/6zN44TFyEvP0/gO2Z6lUf3vAGX61eK7XF2AEH
Muancw6hF7mScpa5lfPMvE3cHaqGCNZidHe8DWl2IX9BtiyxD5wqzpgVcS+t8lmR
4aJDTfv7MkO70WZvAYYU9A==
`pragma protect end_protected
