// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sXFtPllPykywO0C7mH9jhwwWwMsIAAviD77BrfTcYkJorj8NC6Lh2dQi+Y4Gzn+B
V/JQ3WB9e/WhG7uhJ04aQHB2FSb+jLvBJOJ7+o64JT8NFCSrYUD3xGVdVuKFldqo
7YoxCqxUjLsHwURBBOoccXea7kaqBVOxAzR/M6mV6k8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2304)
WtYn50zI774hWRrxb8gEPhOgj9k9k83q++ZGgWnVl8K+OlCUySpB7MzsGQeRuok9
T6OVAC0hLbRzZQWxwUzVWGqSbuJJp9LJ1MWdkNYuiYRp/OuUaSmCuLRkj0PGdUfC
AJNQJam5kNjWvmZQjsN0OvgPU9bZRwMx1/KDx2x+irZO/8se6u+zAWtc9TsZN5xY
AMPcn0EVNGx0MiKE4WBX9EPyzAat63pJVmwbmBJK/Q8odOUOpmGbsLTS6S19q0lq
VlwAdOVXbyoEN5KrplX98tUQyHSUP8PSopNoA+YIlJn4se0iEJo9+cIPE+BUigmv
0tyQwR1tBQNkRhbxl17kT0EeCRmW+zI4x/+0FLenw2SnMmn0yW0Bpr/bqgaUNizI
3xlM3eGcquSyzrmvudip7calGk59kjl/k+/yTwAZ71uR8cSKyKjV9z+Iwa/7m7yE
6KuPfAxG6+8ZQD/gmmNgCpcDOt07EBAiwdMrhC/iTl6TXO0Eh4LLcZlcc/NKdQVp
H7BrKfGOaNSOPLKBWJvOS3NVMmsa2ZrKTv6TAUj3AGb8lA3RIlAYJQ5KBun9rtkj
NBqap/HJFGu0MoqExrezRF4w7NRHqa3WEbfHzwjBPKlvGSnPIXg+AQxg8qn9l2o+
K0hFRDDHnn/T29PQKY1dHpyB4mpNM8cdZoZJbqQ7lzcvWM396rBJshIf3SHvGZ6L
dsg/Zao/52uVU1s4Gzg3r4Uu3Ieg/dlk4WFMLaL9nPZeizIk1Weo9rCPtp4zMtrC
jN+0AKX7E68QLiaOshOGbfgzPpeWV5XVmVdUpcDoyMF4QgYPR09ZpGIa2LbwrfJs
5XHF9FVHiyMWCHDuat9pMErHlP0+qlbBZ7Bg7NIEHR25DyR4JrIBvMcrgVRSDEiz
QL7Xc+LWERoTuZH1B5opVzvWwK0gLtyEIHKCTDINPggWua7OK5heAbbVTpTRAiMX
hpAiucEEM7VC45ZSCZ7RXL4SjNgSelJOnfX9jrCX9zHoVJB1DhqvVrDL85hQ7Kus
Ub7TCsTNtmdEXLlbm/mI+u8Mdre8np/Y/+sDemaz9gXCF+x9kRzULw6VZ8p/+9i6
aP7eP5wNZu6NWy3QZqkXdeTG6WbegvTvow2CMK4LhAR5En6zqGk94+C3jrgfTtnT
fhqlLq6kTJMFTCO9lFVkPt5zkJUAxOMa2kqvZ4az31KK3pZDLf4jgSH+nvYCMhD5
cASp8eSVCqpb0L1zxWaLOz695dKLpMex/CS4PNV3PrYI4QxVxGAhXlV5SiRbIuek
t3+ezf3vITDm5PuXSWcvvhTGbKGXRtFnMnAbbMwF4BYdj3DoKYZh4qlZYZ2TrQ7P
hdx0Wxv94ipfmykrJegpfRC60bLavu2JBxxVGxcwsqfbK+asXM3DsGQtYIjzwXQT
eb5UreZue7ZAiReugQSGAhBbUbglcNxUQcu/1HgLCP8jKQ2gyEbofPi7VSoCteLa
wF7qVhqls346kZ2cfdcuYqFRtGFHA9i5DIjU0BhfD2J4r3l7nZTDB1pz/6XUUtbQ
jRMrlEtrlU9qXjQD/UdZXwVzQQMJ9dkmX0lez22mMcSXjzzMwm5WU26LllVzbaIW
p4oM5MEC1Q9qeDhkzuZYRLNJ4P693pwvlwfoIdlJIC1+Hh0U5gOctZbEdytr1KNA
vACNnaiwiFuMMpXiK17sNxCVWsu8OY/chNckxV4NevGG5bT4tz9JggFI/ymJFWEZ
TM8QS9MC5HYSl6qYqx7TdavYU7hRE7a1UsEw5dmzmTxxNx/U18B+5n+IYoQZslFY
Q8/8DQY/TBAdw37yMeOwnqcxR5cDUSpa7mIiVlaOIH8kQFSsTt6cGttgGjM652hl
2Gq98oAadTGey9yLfRyORIsQKcGcvFTAWi4adHCHFUAV6OaxJiKMexxWij2v/nhN
u445exDYhF2HU4EisW0pSTDxqXNpyviX2Xteoe993NJkZu56DpKm+JVGsAJvfcab
+mOkiFtz9VlvFpIs1MhH+ie2c8jTfEjkjm3RDJLohJWvk6TIqim68LxuuuNItDWe
W2VNVZJ5PpMxjmz00g2yfxkby5o1QHVQkv9i4c5vs1F4C3U033mOUSGqEp6Kc9YW
giTOexf/2/H4AzLA2BmlW8l5sW5SwVTE3Yz7qDGBU/lmTtG4mrAtm8N6Xf+R4ytw
Mq0HEYAPrKmRnZUnTcy+vjzIC8NxHJGvRixdGMwK6T6zPAqsjIERA3z9JeiHlPuH
VcvaUSp/6PAynIdMZ2nOxyC00wUBxsM2N3PvfYE0Q2MeuwnJYVlpRirm6BtD80pL
WDuZOToySCfmAyvPKiJTTp8AMjJcIzPo3yFukbi0a1xdtz8/EfaWrHFo1gnIyn9L
IygA2tVEBuu/CAiXk/8guHW/+aEtQtf4ONzu79SqcRj2Jw4emeiq3ZiZn3FQ00if
r6GZFqwOSJ24g2aica/tB2O8lQkTL/m7FH4V0AdtblXY8vKPeDI6I+DJpbKtz3H5
ttuVbv869mGVN1lSBXhz3l2O3uLsbRDVL/TQz6ZvMJBLrHZ3r//hGeZUpIz2P1sZ
oGv6nEtZJi3XLXyPrD7q74XWku/wVzyUgMAR1G4+oUv32zRnqOPQJO8b6DbGiEYq
qsll+p4aYHruw/ey7BosyjygAiG/pewOib2aHrEm35xVF0SKYjX+9Z7go1PYnsYO
OcO+OPGpGT4nTgYsldWHunj7NuG5uxrKkd3u9pPpau3ToEVv1r2Zk70ELiUjH54W
dEpYPUC46+4Fh80Pdx2Kj0sdH6jY/04MqhRRIylV8TSLl26i6OFIybKvRdat/0uZ
pow//wGM/kLSGMiSua6O8ROAyFZfvvqzvvYe135Ps7Q/MF6HIlsUzQIW/96wV5ox
urymgRTeiP1+IYnH3QYe6Z2wobgN9Zs1+m5YCVioEV0oapa3XaWQrRxe3t8ZKXfN
H2JmhafrvtIDK+M51QarpI5FAqgyFnOADIrnZvgnhcxFQ3HLCN9ddVPTyNwwnFoY
t9OxOZDhWVMd6oesb75n/LL8Uqip0X4EMsfFoD+bnH2aUbWBzTA32g8iYwYTalbC
`pragma protect end_protected
