// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dh8izP02RssyPiD2ZO+umAni837tQP7LTZuuzs5M71tO7LVUw5cBdzEEf5RfvfQs
i2atLNuf/KSm1RAO/mr34z71ptVHbmeJwEYp9MfH0Cjj3+ZZmimXGgrJuku+o/7W
/BxcdsT51Zc/X8b9Ls4Z3HbY/dVB2vwhJVxkqE/kY/c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9632)
7gVMrVWABkLOQl7Pe5J2bGKc+lufHBq01VEnsSMUREkrqixVj2Yz9y3JKONfy8OZ
IiWvJr45zvxUD+KXULIKL4OSFgwVOCyg74JJfT37WOO6cvamk+P3NBWw/wsCvVLB
9aKb9H3szHB33cU3CasB3L4d3PNOC0iLbPCLQUVe3O5VsvvHE76zTItQFb1I7Mt7
qJtPhYIZB3tUE6SYe8yOpnAh89ziZWXmq/3KpYBRQhRriFwL5STOugV0OBbvnYu6
5ycIvBwnjzVwV/r5rIqbKEAyY08scDh3GhCCovQ9SZLq1t5vNaswC4aHsw84xbF9
IGgwRK07vDFDnJrQFUlILqZHrlZkHnCV3oWo/skpp3lX2Sa0Y7HoxqVzxeEsxKJ4
eda9bvxjwhvCGsjZfQEcwGNG2+ouT4r811D7D8p9WMzfEPDAgNw2cMZ9kKk+qsXv
wEwb/FbO5KO6ImMqLU54SpMLWOUZoS5VMV1aCLoixsGUdshJ+xqwZOm+80A3GSj1
M9IU7HiLWgWK66fZMAawiEeu/asKiKV7cIgR1qMtQ1xvWO9E+5JZYxpOwGm9cekM
v2ALuaGr59DwOjIAfmvT0sDtEtKtU4Wbto6lJDp9KrpCAjePAHuiYzDuQoZf+9+3
NxBhxYjGzn26TuV9SuDCgN7yzqIXXWlx+t3imqJnpU+fLaDYmh/48zgREUn89r8y
W8Koi+a2yzLnmesbIfE0DmX9zfndPitOXRkNQv1JlW/BA9NboZFO99aYR+Nuafmt
tgsRMIdVj3M4c7asWC9//oTkGlFv1DcKJicOf9xdGz9uh+mqth8wVAY1gMmgwoSR
q4cZzImeq+2LJQR1Go0IeKiwKFPbqBsbY+UKcsI/+B8llol61dIMoiSK5LeU56s2
ramGfrH71/TzBYBcK4h332WoAY2h0rzc3Vn9aE+UL1tfOXTxYyE4IYhaPihfGw25
btNlDS2H3PBnATk4kC6FEcEWtxWnjU4/MINK0IR0v8mibRtuhW5WNetm4mZM3uNG
Jf0npGC8TB9YK97CQztrvNXT/2Ddz4xjLpth2LtSyV6qceP04SLt1/UUglOCQ5XD
Kmedjsn8Crk6Gx/JucDg6qhRNUOYYcJIh8imweOnY8yZhmIzw/QUK2MpRarnwnPY
9Y+iLgVD0bNqS55X0DZcW/KgpgKzeixklkLeEPWGysbd+cP4TNQbejLflbReIU3e
zeqZgLJV7YPgG3anKnzmtKwSr8mUEim4poZX7joE5P2sytLgGULvdL/eYHu5jEQq
mBq46uuMQpO8Cm9JfdEGGLiZHqq2S16SBmeF6GVWIISG71aDLhLF1zge/WIHz2GC
EnF9i+clcC9ipNyZOaR/mzNAOC1t/+4TPEtgo1YBPr1HUkzshSoSDCog8Di2DJ8z
JKER7g0Vr8NqutnYx10CqPXhJwIz4dowt8xwH23inJXbMVdh0yDx1Hr7DV4qzEqO
ls6jMZeiNqqPXPM/kRVnRcrmRV8HJ69VNpHZlwsCM392qYUsZqW6Da82j0lSNpf+
iEiS5LebDszOBS0jlsQjyyi7BvT95QnX5aB8KMxraVBpfLmi+q+M0bFf0fLDG9Ep
txfC5JKw03CZG229vNj3UfVHSlCSMMP5MtvCT5xmI5XFK3n2dk3RYkuDK198y7G3
j4gVkY2M+mKznWwcS2HVx5nF72cjB4RbYqmlMaRZnHpcGh3iyqSeYUtSXtu5157K
/8VeNKK/CjKBeoQZBNbwn9hG4sJI7T9D2tI/ZnekjF9hY9e+2MagCcNNgQBM+tdU
zLtdqIvbsWSDO3hhj6v82P+xf9KErIZReelQxvaFYmB5F6002ZwcKb1AXnxZpgTn
reX9E3iy9E9bhfNg9VgEzi0qV7A2CACmSwijxph8WQ6oXZFZ4/FZmxRkmJh/yllB
t+nTnL5xSusmq05Ivpecd93snE4MxNRR7zP68lpqyX9WwR4W4k12DOJGnKble4wU
Y3vQXAcjrYAvM4EqWsN0IBSP/Pm/3gDS3k/ZVBjwU9PEJIAXajvE0CQJZk+dp76a
8lOrROR7+3vHCp+8yi/LiX3As6uf9kgsiXKRqkntPU7RgoNg9wsGPHtdeg8QRQWW
wG4wguz933/5A0jF4Riu4zQlYSmpwOOf1EpFTfpizGp3rLJI6MDUX2XJKQ2i5lIP
DsKTuVIqqypR5V47ZWXeX+xUfyy64vpMotTFQYF7SM6pJZ0woMvmUTfEdn5JYoTa
B1lwnkoTp1I232E6d0zlxFqNVCFDknIf2TRN2sNvX9AK3nLgd6rXfU3WQg0OhSBR
f1LugGIuu29fEQMrBN5V4FfjXhs/mKsuhypu7h2m6hccph3GdQ+w2E7wa+dd8zte
vnVRHYzZknbgsy01y5kp9wkwyM3LAefRZzjgNpjvAg8YrOKx+HdMw08b7dlVSp44
8pnfvbLjiXBXFP4/BZ75WIgUeLaTKhLnprA0tD5ymieXmETZKmaqKkYiBHvlPD7x
tVKmV/CJZY9c3Bg+zV8D0Xznm3UwZfUCmtrLLSd61bh7p73sU3MBHQevbbBK5gqm
U2bsJMnk944u1Zhay8vRjoLVLLk8gkovAUzJKmgDTsxJkCSD2LHH8Unc5DxtoNKo
enAm1f8lNdtDZUkRbd1PBVse/GQV3jGYES4xKyZ0Hov2vwpTqMF6IfAFGdCnYTFs
/eI5CEkOrmapvQw3vC9sFZxddQ/dL200oyzNB/a4EqUnIm0hezKLy15Xt+RbxOh3
hlyEvZZdwmm0KX0g4Mdhf31S9VJ9J3JRw3rjb4NPi2Hy5k98ocZ7dQE6wsHy44YE
Ba340vh4SkpqauzF/b3Twb4ydTcTjD5M6VEn3SSHwT5kFmJp4+dsNmAavF1v9a1Y
XHkx7//MU64Rj54I1+9hTA/85uqwtr/d8Srp0cGdbbPQhUEwcvBDe0Bhjkl0q9g1
LbyX3wLvlczBVs/yZs49DD8jKYbN1sHnWagQQ/grtXuHcOWFbEtcRgwCCCg06UUZ
rWgBKl1XWHK1yL8u8uh9jyzjTf+ifKyMTskHNnL18xxglLc0VJ0EYXklJD3TmSq6
H+77uX2kaWIIfiWXCyzihH1wDFSxv/cADL8qTDrEmEKSmZOMLIlBMzjx21ggD/xE
oouiM57Bsqk9SM5bewsytL3OxY96DuT7ovqmX9vKYcKLMgumcGFCvv5qPupYF/Rl
Pt9siXnnJV12Ap5MT4GqvbkL1ymUnGLpyPdk2+OnljASYjOgFuCG6qw3imICcZ2D
dmkR92K+Ix4r9EcBY7InWzLASe02IhgJhuSBi7YykSm+RNMnUVjm++nws9lb2n88
18Kg5pLAgXnk9wvzMkGyB0ybtI17rUq8YM9ks7V/j6WMveg5CQKVDesL0d3NZHA2
kYzBe27Di068iKiv8XikvDnGmLgwtHaeFlDH/XdsrI0QH/dp7ZJDNGTCFw1xcftg
gHmvMwMqHzq0AyA/7aQJjEU1hPg8drGFOIT1RvProziH4EC+21cspa+Rf15YWcu+
U9wnMXcasG8yt9lOkkKEC/+ydG1H+JwX//UZvWeUgIqCtsatmyqZUP6SMVD7ILHW
M2aJxQkX+9iB+Gythivn/gQ0ZUuk7dXyQCmF7gsfhM8fYdPf57nwp1d1PVpYFAUA
CvyOv7iY4Mn8Uvy3f3QqtGbvK4oD8feah1+8ejlHsCQ7M3AP8qPznPZBawLZ6TRG
2a/YIuO48vdHN2kpZ9LO3bc1cIfwa0QZtpmLamxonjshC7Os6/NXK2L/AwoW7kG3
Tez61bK16zO8iqnggbwoMcdv7/CMPMDlANhsOXYCPppdz2RA+DiN3kueu5Mb5OQt
2q25FydCO5mYSqHDm4VgQf18bfu3Ah85Q1uuK6W0SX7PUbs5ucJlZ1krTf3sAKC3
lHUHzVhB1BoAj5RD5vbBoKpuem8NRe1HG2kzBW+blElvrb7MZ9We4rceNPqUC+HQ
R5OkZG79unrWMR0sL2ibldWKvrJ+wZHGT3u9rwU3t9MHgxmHY/JWVkWP/dStfuZP
bswYonPjb+vw8+bYIw8lKpBXW3I7uEkjHFtKfA+pWvzt+6y3sG3agPz2Cqym+1Bp
9IAtJ4x3r0G5rj616aoaktJfeIM8NsmsqlW9Wio3b4y5DGdz8yUOsTgRQ6HDiWeu
PCYVjnxrCVmOAbh+LZt7M7tT65JWA9ooJyo+ig7Cywga5e7FSpOPWCIklp12mTGk
NQ/cDWPGUrI0/9hAPRQQeRDACAmxiOSXp7FQjIFo0PJatmowSRPBSmtxSmR/lvfL
FY22aEjPmGs6DmubR8+c3nUPoZWHqJGb89w3byG5/dZJhTViyDjz1zVAc0Wg5ijB
dQfkr1r7FaId+yPyaNWAr+jajalSHAETVRUtC4qEsu8c5vsi1y7bWoYe4TCAcRpa
CAFU/v/dsykEOBqBJfc8ib4Z0BmkJLlhxVSX+WF5IGF5TiuOuAXtKrambJkdUUiB
0SS+fREHlDLZhklVwuYgO4vMUCpyppmf73dl2sRl9M+jIGEmpWG/3kifuQCTXXHE
h1wcqi3XclIUskl1PJUQ2z3oqk4yIg9MgFop4zTc4Ngq1ukjcXk2wBcAzQp1BBZf
FOtnYpEqOUBaknid/xCw4rO4Aeff+/5cG1PLHV0WohXxfMd8cucOlk5k9Weqk1/r
qVHiOjQuyCaieIFRHyj7td5RcY3uGsoItGDReEx6PZ66VzcbCpM/4plvRB7BDucF
MLMiwDK1OBYAST1xRYewZn3hePV49coGy4UX1mZzi+JFNcd8lQFlsn/zWLlNkYGW
IvsaNu3va4YyM9/U/F2bzR27HAaVwxDVUE1I1/iKBHJh15vAD+hnvaS6dZGfM0qY
ijskXKc6+Hl3eN9CiKQvlEvOJCkLOn57P1K9SUIRm1GngcSL3ojbC65kFLJte1qM
8sxxJK37GsLomCjr9vBKqBu+LF4yDiI2QQSdpYiDlzQqJ75rA9Ef9KstAmna+cXV
KEGOuDQNegPpP5T78sLPo57sOtHxBM1ekvdw905rden3tPITLrxSKNYJpcmjwfp3
AdWALUPhPL4z4eC06WoKxRoHXtsT4jgGz/JU1eXR53cYUCiB5GnO6ApwU3Mi7MMW
gzGzOJpjnxOL1lgsTYZn5QCNNsYsRJUSN1Z4HRho0Pb6kFR5WKC2cLrHCCdL1mNJ
hpTE7nJA7foCQYR6PQlwPz7rNftkHfKuTEfmTYmh5fGSJjrArBjHVsFAf5cB6thf
DXyPrrN2ze6VMtSD3SOa863oEQb0j/T980D3tHSLBSvLwHQHuUCJFZo45G3ZV8lG
ny6KAUZUQ2QUsKSFhyDQeAaz0tKw9itEbiiC9mzxjRrEM6NGXAGPt0Zg4PJ0tsPj
SoMTqT0uavzUjoC+U0dLfWY6A4phcMid7pbCbyRyAjTwxS4QWKLe5629VXGb3bsV
EZ17BFcr/ir7qbmIviVrc082gpMItjf7TkQ4a2KJCu3McEUcAs0A6YSwhy8IbjlV
NcsYi9+twmxjooPlG0ZhgFb/uHzsUDtDTmexsUGa+OwmkuaGmMGPhSFhGI1shN8I
IVUPS4xZDaxtOhdidhlgSfR3mA959z/mghIqLrGWMhlwvS9TB4xtF6Ym2Iqzurx/
Le836ZjgWcVSwS152lseZ+8hJ6yF6LDnOjXWrgoLO5s5ULEzm8gYGyuQnxuCGviR
huLHxE6SVeouKSCXM53H0IJWJf1OSvDmOfFTTvZLnAwM6wLygcQCD1uNcHm64PPg
XAQNrLS090YX9X/f41JTF0HpJIPD5WtEAvTA2im31rdc+wQkh0zCKnDtkbdVv3CJ
9540gmbg0n1wz3n0SkVxrZhA/kR2lwv0FekkdL1rCtT0pICBISOeN5+Y75qZ27KW
q/DbntHYsd9kgiFuZX586S6EwIcyZGd/mXIYDz7BX4aIqdbrpNoOrWYyApOCWz5k
J5lM4FLqhd4DPfDEu0YVGnDztMi3nAfBM/AVRAY5UyzvIrg2MxN2yI1hwWLKf/3L
5jCAcQIZhTacYALqCQIrXT0JHGXP/RJyUfV9XGYz2eXEdUyLMg80/EvRdrOy9yPb
nRpn+CA1VmGEkDLdO6XnOwDTlLvpqQqfbpPqiLSBFh3Myx1Wix9r+oQUVOIxhKPK
+iaDJe6UvCcDXjw1v59tsj5of6nYcaXQXi6dDvL6GPY9qrJuHITbeQHcm9kFgoWQ
rf3/Op9+lo3HHoTD3uWDLj9ZuG6u+HzRJiR+oXmRe6Ie3sJscfyLWjYma/gxfw6A
nBEqOgSWPHrnOz9gxf2rYBURX51PjTAqfzuul+CJGmbMJGXhkqNvONxT+CKiow7J
qCbfN4tLty+7PZx4ZifalPzV7wqhehlFoMwreFqXnWkZHQHs/OgX2V46MHTY4SnS
Y06K33Ev1ty6EuihMvp1tdL+ruQiHjtWt/Zbug6ioFX6EI63BlEu9Gm/uNElC7ZY
1vozIEIZ4x0ANn7HMChY1KqnzxheMh9+ovDQvRGtjKpu0fh3WhGe3ZeVYycEGebY
jQIUkeWSUMSLDLACeVOxwXLWaeMvyTWTNaDJcIzBQ2BFxHqEHSxAY3h/9TEMFcte
+H02C2Li4GcvKW/uZchOE2aAu2Ml5kppPesIzmUiF6BUTpeivEmj26HD+yx5w6v1
S9yFMtGlC9b9FXCi4rFMwaWWSfdWcKT8zkl3SR+yzchLhiRPeAHchV5SzkljeO1Q
FKqmE2HSBesnj/Vt2P/84dSG4TN7u2t1F80jG0KZL0R4inR0CnmdCf+wm2r2XxuQ
WlR3nh5LqTvzye8fEVlubiujJVePLdDS5+lPVGkwRw2TDK+Jpmnz/fRbxX+3IHQx
smPONyVSbDCwTeeWdi3GFlGpaonJGdpBtQWCIadlxyExSRyqcqI/XuXf8tdvxPo6
d6M0lBRYdaEpQr8GoasjpiSJblTqd2up6w0gjBRkMK3X9f2wvNumfOTQJhNmUW93
qKqZ4wX0RQX9ro4mjIbKduTl367527Dtb8zL3hpj+kmjsieRuarCXEU9urFa0zLI
bsF9fS39Nr+ZwBrii6MVCf+GkV2BOE+oNCKgKrRA2XRj7Vr8qU+WqCzS8eMg5D0N
5J1bGK9IQfAN7uK9gzWeM/q+Xj6irT6KUwSBxbCWy4iSu/X/QtsG/RU49l1HDHxB
cjt+gge2Y0Quy5x6hVFJX/doVSAMIDQOJj74oxmwxsYewdHQOnVQksfVGPPjn0Nd
2/NY+vCiAxKFxKt0ERQv3fiXhqavWYPgdl1ZhF/GsMlna4hUZmkyffuEZMhuVL6Z
SWtrHZuwkY9UAkKml5QenCg60r3JH/Ji07FIWGzHTEceIDPidiG6a9D0z4t84UQ+
b7c0gDOyc0vWPMyz6AURIWWjCYbvCAGUMVxSKjad/VPBqgqemGnwyEhGLC5Welzp
i4Os5weUSoDb1vTCMZM4HKlS488WyYvAqKHVh4bWQ5pEhJ/mlwEjWiSiGypSRwRj
llDXM3d9CBifezb0WaPZd4HAqSQQJBoCBMCW6N1TXmhgzRXK5O24B0ro0PAwyiaF
WONER9q7Z2ddD7HwSCc4iL101VXxl8PwgNIl5Wz606CosHP5sHdbgt6wi5OC0R8O
fIuFIdr1OlanBG4/5ykOOdLYiYFSiO3QsgPKdZiTMESeBWnFmLjtZFMORjgpmb3m
+7NMp8ci9eO/Ak1y/xjyUTAogEEA7XNt7OWbFVXV/hhI8HUl529/rQqZmAXPCTGL
FpSXy0lL8+s07xL48IJIP4f4n97fUMoZGyNDWrflRT9zJNRg9ZffB5XVnIPs9OMe
FYty2DeDUDqBuse1ZIzmoDGbKWVFXOyXs9QZBfniktCvPSolegpLHn3XiYYO48zZ
eBB+DVQW9eFpjLqBbhgm3kJxIHc6cjjJeLz8gHFnQ8/TZ9N8pk/t3QIpXVvxB5Di
6es4ii5uUI0op9ukMr7/qn2byqVh8o56dRs4KIMdX4McDXXRvh5oO0El38C3FJn3
KwvHwZictcruCAEFxTMK6KID5gQ03ErOY7qLzXwRgaa/r2kv5RCUAvE37fX1OiFm
rzOxqkxCoj+lTqIC/YKJx9Z0vRciz4ZSAbdlhvlOFvEX74DKErc1RRYCFRCQUj5E
x13fcsH8nogOstallS9QZA9NugDpoj/peW2/4vJT/OFAOYjlgtGe8RCnt2xy3y5y
VXkpxFOrGgKQgktrS3qpvCCFKkWNVLtQfWHzbqw5dhgujKXGWmfhdJLP8GFrOnba
MZ/emuua3XFIpqqvH3OVz5KvMp96NlIDh9oZsGR9QfGMgW0a1bMQeQXUjhVwR3dy
aA2hgbJ8djZV+WOQF+H4Yma/EwlgiI/0vHGitkDfpn4h4lv+0xkLP4hWZ3Vc3Cx4
gHFJAUFBtmvo+bvEAnRV9Zz4UPEcS9wpvrgTRc+Z6MphENgVuSEI3524LUXBYoI1
XociKUC4/NNl+yMA10jr5vydIyzX2cl3V5W0k2nAK5CDPk9uX5NC0yChwyOzHHom
ssZPxcZg0GgbZqYWCqyjcKQwtHWU/FhveenfWEu7CtdrYQE/o8yOGAiVMZFq8DON
fHRr49z5XQ8T4T0J2zlIMKDllGOhWs46MKjKBH1OXGQVJXhnQ93LCdmd6KqfwEmt
i6ddvd5cHbAMSvQeLYxcI9lRfUDA6FlR+iRfSd6Kb+0KF3+/iKeDBDV3Fp/ClmUT
WguJckYDoBcgXJfBFFJDYx3ZZzxYXRTF/cZfoFg3OG4qX5HCa4L9tysrei2gEwoM
B4lu3an1sol5AbNmvC0CAXPtZ70sxy+g013uhQwyvicP4KRk4sqOyHK6G4/b5YRC
/EeqKMEoiTZQPN5yzVhzyZDKYNS9kA7gkCDek5ZJHYHO1DkZdGJaGGxY0/eVWZ7Q
TVUTBNqjNtRVW1scOQHkLluXA6Q+Y8U0yUKmdeicAsdWTZ36Eu1GBAZaW9OtT583
8tNn9lPeJvFHdvOqeaM9OThCLwW0zzj3c+6GEFOBcc74Avwo72mIIkD/IsVSfrq2
CFuhY/K0rbCr68DawdFFWthMgbpPxv0+SHFf407s5NSqm+nRT6ttVbG9b7QN0bld
TA1b/BJNgX26IVGj2RUO/K2vv1PvDFv7/0RgpMzn8gXAsyIDaXjb4E3LjHpHZjaA
uDLv+5r4ua7ULT5/hLEklzzb2zzR7R7g6tgOX4GErg71DonNbXj6E1m8PBDODCYY
1koNT7behbS1UfKDJHD9bgH/abbkeCBVA8sJDo47C7IEHG6Y1xi+ffUVaA/j3CL8
0Cq5ndRSc6RJisNxBwc5XA/6ySVUiIO/wOEdc3SR6uF8XOxVrsAgUIQxDpzxFuBW
vyVMJCmP3VqQJfoHZc1Edm+IasFByX2+CO4iDXTLoCvlY6+hl4zzVzSaHGcu7nOk
sHRcfWbx0vjW87c1oIeHy7uTH8rGA3Ch155fATdC+NoXZNQoWD4AwZ4VQ9OP5rss
dGaZMwXgOGiVZ6wH77UDbplZtZbetcQP5KHv26+bxSTr//KQ019bSIoOnjAgEiSE
qMi4t/YF052u+Wz7Yo4qthPZ//5HgNTuJ+/vxY2Z5dNUJH+Ig6EVEiO2/qruvogh
GY/JBigAPnlIaduXrTLfBHQ7iFNyJyYvsbY1pnrXrP0zg/lqZFd2ZE9FqMARGa63
sVhnbYAY2Bn/v87pxfDMTBu/m4lm8d60PwVE3JZ5GXynKOA5M53Kqkw+IzpK645K
uO6LQK2kc4mRNmr20JCI6W25mlEswUSNpY5HXW/k1joCOuJY5lIx0VTcI4o74hxM
5GE97hYQfeJ1M96Tin/ZUbzEIWQGYS8Wx/V7tWOU3x37b+IzmbdBWzv3bu4t2kym
W9yVGXdnfDOI8c73htdd6C87VceHVEVIxvkceLgXu75JCU9T/60u44+WT9dJhk57
dRRQqQQUEnQQL8jr9wXHLphTPnd1CTsKDOY7RTdpJF0iNYfaHw38TMYbwASOsa1J
aQYBxhCPrGJ4ghV1LYV8enz14PXNeF2rZomxP1P4zF2LJmJdu3AgdIMZzHMhaPVK
f6jDmBzrrxvfjPDMq5j+a7HUT3+ghVF40hp09wSyZlcCYshccei/l2jhpgCkPzeS
cp1ovVB/fc6Rgc/AHgUbqrLREVIZLaYOwe4gWn3SII21p8lGvxeuZqOXpruhdRpx
EXdNDCdc0mscQrGDL1Omke1kWsmUbbnrhVOKV8McB8Puakh+K6dA80Pfzt0mMT95
0lzzn0cxsNePlWuqGRP0V87/Rd6ZV76z+zYkBOwNr3JZlRh/41Ksu1l1yvlVmZgR
IIN0aXQlz0xG2wXSh/A2oVMTM1hW2eRTjvX9JjkJtj04iCz385heFowkjMyJPYhK
bOsRsS9jnO5L2/MLrzg+W1NJQ96QVP8ZRe5yWWOQIiJlPT+vYVcqH+FWB6EwG8Hk
gBeCVPp7F49kuDKApZpYObnFJujyrenaZx8oZNiR6SNDkn2j37SoAEaqZvxxDzuk
Ube9ITCHUfhcQ7CN5z1J0ZHxr4/lYwSAfa8yNFppVM1m9xSz3LyLGUGJM5qMwL+p
w7X0hd3B7t30CHlJzES6EmmMFU3uga7WG83MADVo6aGxHX8fDd08bEVjF2lapGch
/seYQ44QLx7hzFpocYrTS6USGRCz2W56fMHjoprnDAV6mHNwE9F1Hh7bHY8BjdoG
wI8V5jwMJt8VTFj8XIGEOaiyfgVezq7FV7VgezHpnZqn9wizmPmkieNjxFQKHz29
mPoi8d/5eWZ7kcr+d8eLQkxZuy1UFuejrfRZN5DCrnzoBqNq4wGapih0/zIe+jpc
7je6U2s6IcbxEaQaY3bdXsNkxTdk7lrFPY1972CE2gge/KEqPmmP655embvXT2LK
9vPjEp6WSB/Z84I8ErnQPcjk+k6MVjlVk/rxKSV7NXHluJmT3UuRo7cy6zJLZdWZ
pFmcaKk9iLARnoVYCppShCpo46av/geAVQ5l2/4eyxhATXyV8jhWM7rk6viBP75G
8HFhly0wQgkTZ4kJLHvY6Xihu03GaKLGopiuNuVOopQvsm/AdpQ3Z41eH8NHE7H0
bupeSN+WcUyQQRduRONHuDkZaDBvdHd35ngjtv41AE0URjo996Ms4HuW7bptuyrA
xl92vnxIZT5KaRjZ7sg5TGbVQCo6LycuyJawzycBZlrNPo1+FuNVBW4OOwm2w0NP
yRsjRPro6WNYLFZt4v0ybJ4wyNOXZIbCImw4Ct78PLF+FHsVSRfHZuHqq2GGXJnB
rxe85GvuuPeTiLDiwAfXTtyddTTNnIBYUgFcoEmnplhdiXWwZrDwsEXEVImGouju
HolXQaatDyzRWMZPFj+nulv9gQZiCQwHLDUce9XeZNcqVA3dFhxAyBWp6h+M/ipx
uw/7g6q+QwA955tj9aOEPwNed5gS3KSMbl48ObY7BYJBItdCsFBJ963RvtMEQbXv
KrHya5RaiAkjHdg2p+BkyknS/QJI9RTKx4oHRj5Nt8hpwhqVA/MbKRO3puGBUBoR
Q5qm6Mf6VIrdSQoCJ6BWj87SnqatBBg/yd7uMfKS36Cvg0MO1xNxImDgKMGwLENY
F5Xssckc7DMkw1OBOii0eq0eNYTnK/QPJGNn7MQw1PWkdhJTWfpdSqh8Hg17Vm0Q
zTHywEHv0yHtTWqV8mS7ibUmvoHtcBaGXiG9/w0fJsaZABhh5JY+RiloCE08Hn3F
idfxrugbB+gtXXc0fhUwxA7KG1ALdTsamwRsW2z1Zg9ln6PihlxU+1vpifW4lkw/
5FfPHn/FT6twM6b88NcPvy5qZZ229ol5BkncOWuNTun30QE4UQVF11he69eddqPL
9t0MjelW1aVmuSYUcGQrNqN8sXZe+TUl/rMOdq+a4PgSqc22njMYGtUOLF1uz7rc
glBvyUJ1nZhhqbkrqFdDM+UZvWXj4bwDCfyNuQ1ir5JB9CpbmngKQ84eO/jiAP69
OSTa84TenptRMenDNkAsUdMX5DqwEGl3P4Ms61wNKuFmLz7r3+dW/WCVy+O5wZUh
geHkHhPb1en20XiiGVKui6LurHxM38dOasNq1upITA0Us7qAoiuea8ldSzARPQR2
3+YT1a4r3WCZVOfuEsnom5Qrq00CjlzJfUICtq5Xe+8T0XrkhwxjQs6pAluMmYI0
bmR/GKC4FTikFGFZlauWhmb4oE7Mm/p012wwvoosJegaveZaJaIw0GFixFljxbQ7
254tc/fSZm4B6GhyvI9zYpgQqDuadlvTVhnmsgfoQSnr9Y4oRMVm0Z2bQdU7HRrF
QphAUpjsO8KUvwtkJyxaYVQhqXCvgmagFKE8SxV/J2lRiJctYYyZyavrELJhZmTQ
G1cFCfZ1tclwReN+R4nycRsgcHaCPaM/D4mS/81kI4vrT9Ge+hHvYXZqow0Bl9Sl
8lKUVe6fw38Yz3R41EM4cR3TDxhg/jfbOwR0zoY/C1Ip4ioDLGZi4Tf0ekNxWRh6
NUzSpP2rL3t3KkJWI58bA46oV6TQRNK1KOmApscMk4yJafkxdKveDorXGQ8rLTwk
4coBPmpts423Te3zIPxiUZ1xMS3mmZx4EkFwHeJrnyEB9gW09DUpFGfMxnratdL5
0fgj2zeSZ7hBfYByM9aV43TuXYt/u5FZAbiHpd8Z1DE0cRJOa2ZYEjTqZTgue6ON
vyRbsGI2sdVpOfs89e7MFGh5jgPhssMlDpDTkNgQvzgjUqZln6bpB6KrikRlYHCO
3vipA0oHerhrdRsRddxK82RlW/rWrai98UHlLreemFVPHgyRv2Zvwg000CIPFmZW
A3+zQ+wIaI65c4smrCEElS+2lwdNxFuG1CKtCYuwdiQ=
`pragma protect end_protected
