// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oMjvFJNhnMn7cVseDmrR332LsEGZiY5fSysVUz86VJfVufWi7VKNRp9llGrsyAai
EWOrAMdTu0KwmI5GBXle3MASK/RNNRQt0s0ZtZG4pfELj/vY1xdlt8x0G5ENh0Xu
KhqLgNG0ywdrJr2iwpUdNQL77X0qO+KegMYkPKTlECc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27600)
NJh2/1FldN8YnLEhhPJb1l5LOFnbfmw1wvsQ06ArBlf9bMh16af/Iw5/ozJxqr3t
RldywUGrbn+IZgD4R+sdvBdH6IxVvQ+TtouAYi0T3ZH8ZFMWNZiSwyONvJ6xwkOa
SW/Vw6S4aeQEkcLfr33HyYHVKpaIPcbJNGoUkBne2ZdbHr0Lmt5ZlYWwLGszoWoD
VPY1oFDHqzJ+DGTH41W7i/BNMf0WFD70+1aZax9zHg/c0lcwJIPBHwcIahcnU8HC
OQnOVFI93nXNxwitZxOlEviEhayBhLClZZvIwapaloEpIOc1wTBZFAMvFoUT2/fl
n0BzcsfdRier4JRDEt0hsWNuPk7BMoZtE9Lvs1Y31DUDug51iA4+Ww0kiV7f67JB
PcWoU/nfZdFYi/V6MLPaLilJukysfrH4AGZLu6nfQWS3ytnNg0uu9PmI1SKPliBk
u+8L8jzMOt4L+HD+t2Fu69+F2AUIOxWM+UjLQcIawZ61k5D9Gu17EygvJl3fNdjE
Dl4UMkBNUlvCXM0Xp0bq3RMWOwT/6rvWFosiP17q9Uz47Fp2jXIQIbmtS/wY7cvV
182SYOkd4t6Jd1hOdzQpE0ZeHGJRvNT//1MVsKG46CKClXMtXvtXAo4SRZljDH5K
alUzoVmOVonYW/2Gp0sZU5eT/o4jbYmA0V52nlzDA/brDiH2jQ8piXRlnTJCR4Z3
dP3afh6v8xn8qIazNqR2vxw+LaXF5W4DxcASm8bdSMHSq5tG4TSFW9o54am6jHq8
j+ufx7esGpw9VgU5BscShaw2QGswLGXRUigxQSbwT2SNM3sTLTky2vaUSZTW8roP
IossIRGN040meXAbiI4qX1YhHbnx3pf7G6fit8W8GoqjkHUBt8Ug9N6vn+KQ2DFV
g+gfyHvgZqxEj3oueKOoq041++n6E07Eerzgspd3k8ViAvG/RKY+l1KcedGQWkVH
cEx/RVNo5TKHm5tV8hS0xuqUNX87Y+JVTCwXhiSFETqXfyyADzrqqsSeW9SWim33
xKl610bunric3fm25r3OGsiUpMmcRCg9NrewY0NMdAk55xcCAK6EjOcTGuAXVZGM
qXIH+wjhqmJgccKlDLeZ60Vhr51649tJzOJ2VyADnuCeM7BlV+yBAwfO2ABhI1Qp
bhMsWmlyEpSu6Oio1/5GMRQQeoiLADj+tFWfY7HCgodHs24aJPCfm2W3NcUVlaVO
NynvZ9Nn5HxVTFGrA2TWuCQgrserX3dkeJwy9nJJ7jKAUX0uremKjzizkZStgDmw
bWR5nE4SeAKgzOkAFQqHI4+DPklN/lhGI21rkjqB07cojozee4j2b9rjDRNwYniy
SIb5KXyMpPdUKI98N6Tu3Tv/CxSp9nEM8NOdpDYACnF8OgSlvgUjm3nXdt4LmrJr
DAPAhD/LmuTHWrcaUfFTnOEVVbsaHmGCCFGS+CMSHEGfHvcX6rr2bOx3ECKFlQ15
zY8cPhpCLV0kDWHYk75wowU/Pca+/Lcm3tk3QqYz/vjff6tRIMamsjKQSly47MYz
GRSmOKFKDD2oX7JkT4apv9plcbg8JUlNiBAQ61KJP8HOBK+dMiJysxYMPz3kNzmk
1NXUiaxY+WpDMVxhVltfzFn1CsHZ3VDgAem0F9RIVO6pIYM35C7NafpdZp549jLB
Q/2Sv4mbWI29E+IzpTdQf0ynD+m+Bwwh3xgzEPOG4mh58/YDrnhYeZPc+BuqsqsW
ki4++mxobeXccquhSbPZ3GuYVsymw6GbzcrIB3YDJb3+A5QO1HfhYkgoziYISn0P
cau899R8TEpqfg9HFTAZoHE/V5ER1GQiTu/XeYWuG5W0eNv4D8gfZAbBDiZSkivZ
NhB4ogbmN2lsuY175rJtrz7FlorlXWN/kooruYKFhIxXeId+cByVguUKIIlwhUFd
7L39Lld3POZnPrqcO8/GVT1dVjIMVWBTtukY6Wkgl1nmvr42SYUwyyWEvekU5e8y
805f336/QHuS1qO4kKYl3Q+zX40RxqpY6KmnT3xhNN22XDXdbDFFNEFn6boZx9R8
a0Egjk2Ye8OEVBmGoPY9WB8ElO4n3rwv6u0YIn8RwsOWx8tGacMoMCVFPKPyKtyk
JpkxxF/wPkd0+7Waw3ccOQ3kCMM7fxd57xXpFquzZKLgCtJc8Gpiq+0ZXRYNGBzA
d5FZ9LdYO+bawFLQs1EqLu/gJlilvF8hyXspAFH1ct45lLirC2JHWRLdYGEmNIVn
R8yUMzZCoxbguBi6Qh77uxfJQ7TwmWSCFuHlzl/6IsvOO+pqn6H0cNpQn8Kz+SHh
Wm/P8DL5O1ygM38anfs/B90SlkvBw6oqkTLRPbScLt7JzfkpBnkmeZ47ZkzrI5La
kpPfaNzpEQcV5uPNN2FpH3Z5eAh0sUyjZ9sBjuRlbQLa20LZaSNYUMfVebghko9n
6s4j8svbqS9wdcEKBiBFJj4+xv5JNfJitScvizPwOjXBiN7zbiqnzQ+sSwT4TVKQ
BekRQABppdUfYD9ZlYZp04QGG3LCNK73ExzL7PrE2uROi2QsrcgB7i7KmEaabRGG
uXLjSK3f6Ri/gFWYh9ZfkRMluXDPX6qwBw8Xs+gJ5S2CPsrUklziX2SJ9Nds8njq
MPm3Vmx+1ZbQ8SQ9J37hRP7/3jTGRR69NMQGuRbjEcJTuBh+O/XO8plLvBnJUx59
BgGBd9TIB6NFNCmgwCcklXWn9Uzy7PhXne61hBbwIZdWnGJsyZEYQaM2KkewiYeC
GP7rHzxXoRCnhEKsZsbyGFWFTepb7mHuKgh1+6wUcLHf+Q+/ijhkARNbqYCEnU5Y
oe2m+iYI1yeBCc7kTK596SJ4ONm55y52rBDSL4Yetql0k0dJ/P1uwPXBWSu3yWrL
G+wgp9Fes13LSWan8gwjzV3lbv+mSUFIGBnNIr3t5+XkuXTrB3bgnoJMgfA6XL5v
1+0kEcMJCBN4yK6nixgotDYlcyxwtIxvlLzfzl90wRBzmxN7lEfCOLKqfKeUV/PH
cRIa1vjGb1MB6C8DkwNkEQaY7MbOlD53dhXYu3rsPJgg/tfpduX67bZP4qy0jRVk
iK0pBknuWgkxY7s3ph96L0pbORHx8dzAahqBOrF5OXDkDXGGDgVCI147+7eP/6Us
rvTh8szmVxsKvrV513dKDZD7eOJ4eIkjPRKrxzctgu85hNi7o71Q6w+j1wPT7HuC
Ru+fQOr/KylSwrQ+94dRJz6PD36PG5EOlVovQ/tDzrktcK3YMZSy9wvlkZBWuFG1
q7/UhAbTViQsnPkcOysIpqbpLCKxsvXvYNg5S6B8GF/R+zMvE6y3t14+wMWCtWC7
M5yzcxNjBDjHUp/cxmfS1Qr4SOhLc2hlxIzYlCchyEpz+nBWHhf+XtW5pqn3vg2p
kZjXRoEPxwr4TuRhy4NvcS/ytNNSnnyRMUw40/LF7NvyDr6BSqOC/5IVt3p2Xaut
FfT9d3yneTZf8PaP0Q2+UriVRBRQvnmgae7bqPmSUpcjAGrSgoX5vCKOYD/CR+pm
flJSuIAvTDKtS3xOup+VTW9ACn9XgXOPFo4YkPZDKUFih90BTmSA3/zaVPQwTa6G
TQ4nZDKgdElmEDRYPch+2EXwRNtRpCU8sGCAkjIvm3+FjkVQuA4RpIkMnVGwxRKR
vz+9NQf5t2D2QXA4kRxYWKKuSs1rJjVpoQPN98iAZxkH9g26Srde+ISxhkgtMSl9
uZBqo9cDsMNoyHy9lJ+l1UtbUqHzfITgs5lgZfg2EpbfktljtAGNzHAhftVZ5ZFs
5FK3OfooNND2zGVxxekvrUTiZdc7+tCKEmCjmB3PYFQVq/BgcbGkPeWmmPisXjvS
vRzGDzNwQZJrd/uN3KQbprfscxqnBfd8VuWWLesDC0dj08VctmP+wLeQTt8wj2Ah
StOAG9ZNgGK5yUi+MbpC0bViCk/tQXt7ghBkbUP49A29vIIcqeHNUEjrtoKQKWRh
6IT+tylvNHEvuofTjNpgXySVuJdSsnMNxdJsbBzzeK9AzmXv55BJemWQdI7NXa46
5ASjKnP4YmNM2bdaWUPqFn2HbjuDIGGq+f0gw32x1CkqvGrh0j4JX8HSbUjkz98r
mq8B9Yw6xkYkXJgdO2jR+uNyGyWX03PE/PrXGAu62g5L78PkFgjq/lPDBkzN9BLs
OLx1T7ODlAxWXRA3dNgInu3OFMvNFEj0frXD/9b0Zfu1tCoXSdEDmWJL2lwxM4rb
EKM6/6njeA98meEo51Lnp/xZPsnEIasnE0i/q/WkZxWqFe9ntpz/8Y44+XoH+ghL
3Cg9YGQYBoHfvsUUdvt/c49ABtE0i94dvEHKMwSHSeTfQpA2UUZAHeP7zr4guBVI
afSWCBW/3k1O3MJ2wbECP+xLXOrA+NFY5QoKvgW9mAY9Z7xQbhDhY3f7DmmBCcJO
sX733xQvyxoZvdZpECqQaoogV0LljdFf3gR2BaxPaw3pu2xeG7G4yGKNih6PotMe
551uUdcat3OBkEE3+v7y8j4SGRUyJEYwlPdUX/ytN5gCrqn3sN7Zm9KdV4SXgY7d
EitjFOVINvkebfhE5NoA0OELw5TNbM7SFlnYcRwAdYjMT+VJ8x2kmicX06kZ6sOm
qgT2vbmT/gM3KIA0eTn3QsIK10zKEbzY4wEg1UaO7N5zawGmvaOXyce5GsmJjZ60
5AXy7G9zIrQUP5WGyWoGzdpqxsrryaM9n/Bm2zS7Q719l8uaFjxLhga2wp2bBhoV
fZawCDIs5tqIJfz7AFjPWqfisPdXHTO5Km3m5dPO4Vb3d4DOJXQm8e+jrbRIH+YY
dNkgHS8Q+1m/ulIpQfh+5ibcKkeELUedP2BxyATVpmA2AIlw7OEMOJOVWAxHjk02
kzNVBpKlGU2l4X/mAGZf6cZ8M3bBOs3OJR/HaOQ7JShrktCeK5+tmwpg+tTKZn+b
Fm6dNaIxPg0cTGfNBhZR/v7pdHnjzOvAIOKwueOJBas/D89BlKUrNovKSmzfCkXY
TELI/NgTy9x0slWTycCcaVTWkc3tWD4e/8LPJ9HehzL93plGuRE45zVLziCyGyPU
mfS33qQEf45wuK4tgG1HmY+GmfecUsBk5LH3M7gd5gCImGpf54lGIt4Zpu3TCbxc
vItrsCphcbISyetQvojM7J3SyKJmuIy9y+JsD0n0JPxMbzeabh8QXUKeOba6Qw+e
ob5NzGyTw0xY68q3388OJ61igo5vyidTSdXYO5bdBBMSPK+4QJJ0SsDwsda9fetT
aBJnYRlZtDWEc4556jTFkhRaW5PGrijV0qOBrmRCuxPrYEY/qd3wXBpM9jcwe9rG
u/xnVmY+23tAJ0pDxrOuV///vksk6WXJP8PJgA/GmkMjUQosE5yaNOwW0jHKEKVZ
0zJ5DTRhp0MDQ9AwSoGld0tUnMR5tTvK9oNscwfaXtwfBmfrzQnfUYNrAHJd5bfH
hjoKJfEusgbqDzdbn5/vUk1mkEB1nYZczd5+cN1phNaUTAEEGqYqYNLS1OqjNiLM
YzIOt1b/3MaPPGGEbrQ2HH/fzVWUuECska2FYrgNPpXpcoT5aj1VvV8l7JIs6SZP
KBIP58s0JmuTBsKI8HNMu5hmQBPGOuhmhye8bfYRNiVsENeRaapfSPO0JcsB3W5p
6I5JS6p2mRL1hSz9uunOz6LaAV98qHOs9PuvUTOFvPI/EKd1Gi9Le/4O30161WXl
v0DZKxGavhB2wpAxJLtsbXJYJjc2bILrPROZ8/1c9+3VRAz7c4QFpLzdZwtRFnXP
UslTFpVYNns8V7xLk2mnRsGca1tXi2DMro1xB0daiic5fk0zGmHhoeaJQeRu48bf
g95/zZC+7L1bz1YSo2P2VL9+VWtYb38HIxi2Yodt31sMCCl4rwtOC+c06EbjUc51
ImfKQs5NzEXKXcNjYJrvr4gLrbE8RHCrdlbPvRD42vjvSZpIrRGzfkEL7MM3mipG
XRqVNZLmHqWIt8oYM3f8hm4Izi8zvzn2OxLvr/IUJlc/QdpQiOxWm6Cs5lyYdLjd
9P0BNjo5ajaqWXfbpgnUfoFn/mtfxEFefgIZ+DvKPu/wAcXMcldJ6psltqN94cCn
M9Univ4PgiDND2Urcu798owSb2SfDbPO3wa82arK73b85QrPwBg3/Cwf+xtJboDX
WcztADxBFUpzHgH++uIAYWW5sRSMGHUDsMQ/U5oN+5vLrZdPfRMs2/KC9Fsq/oBg
ekdW6s1ikMyKyMiIObIROi//JCUDChUoig+2h1iGfL29gveOBycGARkfHCLaQrEy
+50i/XE+S9wli8SQeh/Wrn0hylry7TkU45FTb/tGwUyqVM79s7rjHlxo8bL9jIXv
sKVO9vizAJEqlKRpYyBmZQySWIRgo2H560REcYRiNJED19KlMEh0SVrnwpYUAC5T
4NR7Wxuo1xD8PjmThNMGhY15HEUMcxA32AmvABDkjXgsScGwlKIp7/Vaqd0JeyGq
QCHuWZ6v3nAZ+3mi6n/N4dIa5MCMKP5DRNHIt8duHA4Y5HV5iT3dTGq7l/Y0DG9I
QQ9WWWN1LUG40FB+NJzo7/Q2EXgkz2hpzaO0XevAza3A2Q3xTdoGok0WO696VzhD
G/e4GWU4dxBfmxHX0H/FMoGi2ggUhahiWPJSuCLV8lqQIdq6PCnyUkKPeih9MzfL
UFNTch+hD7Fybbw9SC2AKaxzniT19URxiADvAk5xzRTrokh30olyKu5yWEZRP/mx
29/Au6Jby+ySJHwAmNIEfbOktgCa/8WWVdSypteKx9xLIbpeUCmT4W7RgG0Ewt2v
ZX0GmLSYZWDs3pIylmkn4eNWkHDiASXu4POXC+xP2PC8mU3bSRLSzUkt7UH9/yPw
Edgct+mJcaVnuUth8m55MFtUEyXZ8s2K8LUEqb3oiMP03t9k6nq0PQwjbikideEN
5ofgw+JjteYM29eghTj6ToeukVtIOJsOWprEMsN9m+ynupkCgsfLFvzuXQ1iyaY+
Oxmpben7lLjdRCjFfqRKJc81E9cURff1rk56IICvNd5jocNm0DV10MiSPS+6pUq7
2HIcKy1Ef7+PFc1k4RzbBnFPZgY4S9LCQMjL4vfmCNQc45/rk2JyTln9zyZiT/ET
eCCJ5CsWffMUu16zV5x/pg2CMarnEOKX41eM+WxgRYHxnOWInVl2Bg4i2dJ442aV
fwR7g7nODQr+OihziT69BVUJE3tA2SkxqXtY/Z7xlpgl+sk79v+LLk3ImkoZRdw6
VP6wT6BW+kT3KIdVZn8kM/hrZHQW+bXpPXZH4/edAh51TmLvPhzUa1PWw9w5159p
IqQ6lUV6ixXyrydH1tqntef2ZeEebn8rpATDRUY6gmZbVs0XXVEVbRVW4WJSakFQ
5FDvOXTsgM+plV95BEss+2kdZSADigp6IPqkZ6vMTkY1TCAtihRMzT1XVVC+dhcT
a7Rhq8jn0HN4/gTvu5ANn/B2v+b5Nng+5R8QSX8SDfXCGlSkKNDrnvhlv6o8Hs6C
RB/6RJUodWxOdDaxTWhl1fPXZH5T21NAs77BZhCkmfzShluGZVmZDk1fzFwYEYlH
iA01vSP9tqUbF6qHuhqAUK5GAhEnrx2nGdvdrQUiGrOjJYm+kymn7m3VME5fm4tB
P/rB48jdhq0jTG5KSQLpk6BVL7q6Y7ybOhC2zE92BMNZcSzGEWfmhdl41PKD5M0M
sOaITVVx1uVQPUT9RsF+wjmm7T3GhOSa34IKbvufO0oZnDRwXPeTe3R8XU0NahvM
e9M2rAnySQQS5Z6r2azLh/IqkWoj7QTjk5aJsQy98MV7UZCJweef7S6b8BkG+8D/
aRjRROhdjVdNKlwyS4SxUDCCOuUrcmxXZ539uiw+/WpJHC07XVRBmgSgnK2t/46z
WPaSfpV70ddqDuQOzme7oIzsLbP2gOkJ8gZahJHSr1+KtNvyWDxZ4mysv5vWDSRo
wjRpuOazUDyK88XjvEZ/RfuZlmkS4N30JSSlDxSUHhVFnqpi1ie/83wIHGZgYoVO
VEUsDEm/h/3TrPFmNgBnv74VFJENZbhyv8xQ5Php8lfhZPW6Pq8FaCG/mpje5CC9
6MyjX4G8m/xPRaBC7yGcVihFv9pnHwWbjK/k6ETKOjc01Xi/Okg3CZNQem40wX91
jdzwqUhGN0Br5TMa3n953Gan3461GeeIxD8hNNMSEXGxPIayyDlQxLWsMmb9yxo5
MQjDZUC83lYlZ+Cf5VoSUONpbM1hoQrgf4e73QsrgPwvIwelcOHXs/cBSw74SqUI
ui5fuC+RnNwQ8oHP+2S5OEslATpDTuwk2q4Ga8UoSdAWoQnTMykQ5N7EX1ISHaef
ezsw5sXRnc/Z1UkY+A+yJIU5A3/WHTTBSRmxDsu9WaTsWeeaMe/xHSIKMQqPezGf
oFAZa1LOZKUwdXTLNKzVzfSHVnVY/ljh5M0BZ+3g5LxEJIKOClcG+G2fr92HlfNO
SckolC66HQl2rjjPjAwd8g5+GQRXH5pQ67rP+NMTE1afOf/f+Ga8C20TTQy74Z7t
XGPhXejyLbR6O5eUmkQ/URqaE+gog+p3DKw8lta6rWBNL5eC0Fdy0t5CxzyWk+we
RIq4ATff6YqzenodndnScUaP+An6sv1QRoJpI5/akVdJFkCgN9ujB/fpMs6DtZL1
/OLQYH01bCkpJvsegksntxxfmoqCDHrj6+Qj2QiL28DxPhzauQrxaO9ZnyCOFupm
QvG8bIXAFTK13fClbY7EctJNXuqpq/senU0UkLegGh9QeVm6q1hJ58qgz3XnDz+K
Y6QtTnL+rzsQrMEERPkfeOYDXhgrlrasnBxva9Bp31gYPGvmZRxD2zcl5XUt4IEG
GEPethxZJ8hgr29YqAQRS59px+c7HyxHHgT2EzIb+tryVdGNfHzp+a2rDf5mCM9J
i/fCL/tkdlMh7Pon4t4NcTnBgl3Ra5xjojxBMA83P7YVFKyzv0CUNq9YwALQQA97
a35uPGPBRbg6ihevtw1pW1FZo3MSswfv8cpV5vYRH7D2U7SGX6A/yvX+VcEI8/sS
Kr4fq0K3n+zjAfnLT9rMjUC7IjlzEBmULmJAqJYI2UEGdH6Z7Foq8bko81DEBewM
+vY3gOHBZeYeFWlG3DWV3ar3LlM4s+fpBtryw0Vg768UlFX5ej/v+C5eXLZgedxk
ga71hL6nPhBg8yJV9cRsRao9BvtU220e9HyQi4ur11RYWxKsSPWm2AbkuyF+1kmR
Wla9qUZaNtrh/+0O0rJpUwitGJ/WC+I2Ii/ZoR/+igm6pe9Ty24KZp3V4s5/8i5f
vx8pyUw3auVNqmzVufmJREBlM1Gpv0a9mNZQqXNIeG28bbLNCFWCm64La1mLhS2z
UibBmvoJudFC0YcQ9QP6/1hhMsGm4GlFJjArn7y6rMWxx2qB/kL8mGlzHADj9M9p
1ID6bhqtUHNpeLEJ7DbUuf7+9Dkv2VKsDvh6w7wFkbuXp9lTX8YAv/CbUQ9gM5Kp
W3sUq8v3Ri3lXd7eGTEg9wepP8WCZMmWdtIXgTgybRDdMpDnfroBFoOZf1s08YDt
cB4fcQnoy/1EKxMWj2xy3iRdYJJm3aeFiawjZ6BAUVtPu/9yRb7jPlnFMHUSSXCn
vPJGE+0fBQIo/FVEg81jFFsihhR4oYzW2lVkS2wGNbxYOFHGdzNc6BYK+RMjjJij
IfGtQ1w+EyoW1bfCE9emuvd8JldFOiDpmbPzTCZaEfHMj1HCUZhHGYonpI0Klfc9
/wWUTTUsKIq+yX9fj2VhdOuSqF2pFk6EGuOhGBWKwFv+umusDaXH6+5YH7vI82JM
GW4TO4QKp4lqi7DekKhQcgSVxGVkknTH65EeUgPClVa58827sfrgRMQscd70ANDb
u6F7JCYsyp8peYXr7lTzY+FdZ1Q8+rfXFzERp81OoU8SS9r3lAwCjc4vzfJOsSBq
wfDKRDTbWmmzJ7PfGJeSDBAgHs3TMBVpaukDELN3RQNPIHPlN9UFW8/K5KSk13oE
LYUt9MfiDhlzXACu4y4mWWYO4DJbg4t8ZmqgWC+dcrKaHpmccg48LGEWZ1+mco4z
OOTalaZlhSy4fluwWz2vVre51JovbIsM0sWVPOJMw5EJjy7Zv6DsflmOT9jj2xQR
lLSgdxBs0YOhU1lWiPBu4PidPXaGBCqv1SuH9aB3Fgj065WiPRsPhiOoz/0tqfgr
OwX6Gsh7dSdmuMHnHqbOW/mwng4AyhLQJqLixg5wcPS0+T0TgzmGSxhjQk4fvnOf
d/EZ90PXnVzffYx4E6/5ZEVJsKbmIQod7HfkygrMDKsGS0quw+mTdf7czwUHqrQZ
b8AsE8+VngrFL/MU5xAaePsDzsdwLzv/ZiF+in2izg+ecGD26a3bV2Praq9r4ScT
Gm8O+um/EggxH0olU72PLR9QUv5ZTcWp1ihtGnqnFZ2OGlFstkiJWx2pIUbDP7TW
/DBXcEXbSt/YWEpzjYwSKI3aGPUNkApeT+1mJPgOkytWoH3E30ggmtKqFcfbhTW7
h/tpZANR8me+oc5aFiHoXIbM3MiO/SQeB+bcP8YQGWUoKoGkwd+HM/+N7x6/P3CV
85dOA8WpMK7emwgsHIyO6TUHaR9vSN5lBisrkaJTU9QgqmAK19hXFG2215OuNkK1
xsTQQ3Yj/356lLgo76zsHWaTeqgAaS3PeHA7kctSpJuQ7cRPHSVYx0U4IGfmCdy/
v4OyPhrDDV6iBB9aMrCAdD6nxRWuSG6siNYBedLBTDv+eNhRRqqC7YcisfFBIH1m
MOx1bGudwAHogAeIzwIQJ9vHR4UDHut6ngXeD3xUgKMEtPVQmPWE4UX5OYCVejTZ
YqubkoAMdWIdkKZnPQAZTbC6vw0LzLHD3571DbCU2rflb5M9RAu4hnv6nBWdBOQ6
DrnSCyiMybpB5sWO+4sAcyRo0oAErNiToZmSwNDKJ/wG+61DJrLwDhjFHzCeGzC4
mf+p0MZwBil6wq/hF2jbrrhssef70aZ+kMrlP7xHvLRBfF7wXnwPKCRaXl5yYYDu
cBLCaJBXPY0xfnxaZ1tMC6dJI5qCPLhIcpVQkhdMWsXX1hWvHKlyXXyoZ4HTG5sD
J1vWa3t80i/Vq38MlkUidDYqxFY/BvVKlSGD+fJbgXlQR+sAwVW1oAJBJEjTqvCo
QxqohJ3LEsrZ2m88T9VpwCL2FUbcfdwDmn+VXUL8NFyFvFO4hv1hLLqAOY2Jd0q5
rVQkjwVvTsnuEMRZXkfeEmQ5coDfx7cZCYExm6TT04MHz+UdWe4Sv5N8j8SQANFK
9eR6dXMNhof5HAClNog/qt/I6hOmaCvkltiOTxyI/s9ZlWkPE2Bil987YPF75WVc
AhIC4sA2gdw3lYcyDV/CFYiZjdYG+q93ftQY46z6HAOiMK+DytDXufm7GZVPf5JN
y4xB1U+ZLlas+3NPFDObkBp20DqDHwkCSNTHavbVtl/oXP7wUEAPGYYHxcu9mzIy
UVGl93iS3EczGBTMl+bbbRYU6jpYoPWA4GUZ9IZw3VLxM8RPSsl2nBV6KB3mFqqK
HXmpMJmhBzd+nM4QOWT70mEHV+EjXU69rmksUX7mVyVxv+6HpqGuyi8Zxz5kjYLW
nSyitOW3aGpwNFJxa+EC6M698irsjA+1snblB1aMdYSkA5GYUbqn6Ar6T3YGW/O9
TWfMpTN/zCXtO+4TmnJM7Y0CMwguNXoHSzv2h+zOLhHyR3XvM+7ba5piFOpasFVi
ijjiMelZE4xFLNkCpPA4RjSKsEAqApLPDzGziwC3apGwHHAiKE6mCNB5jZOMTCLG
lHR/IiiHperj1g/Tlv2Zy793RrH5ptfH8tbuOxLokAZeq8pcV84IsnzxghFHoiF1
4y1PkDEzv26avZvAgERDAjThJUTbdqAksYb2gIvYUNgveoc9HllVXIkdma5tmYzX
VP4HLyG/hynjQnhYIhHG0t9R/s0Aw0byS7E+xKvCa3k1Qt4iElakbZlTZy2adYMC
WfFllhBS45VHCOUvNcWFzhIY0BI0nu4ZRQVG/1IfJh1Do1jQeUNv3lRJlrD9kXWy
o1WgFNqzoBCtr7y6mlxXoqidQUYbTaXGkWupVuOEly1jsUenWCHu+U2UbT4YmKxt
TfMmOt0BNhKayFJTX8DqeWkk5zv5L7BQJW1AJWud/hCPuSzqoqLYMFRuHtfoh1MF
oUtLVoiwvwsVnhs89goB82elDESEEec/ppn1cAQYFeyugLwbzaXyVHjr9cC2mFSx
k7ZYaqsyHPS0ujcUTaCwk+RCiY73qXkmiH07hsDR1gKJdQOVE9PocBawNngO4xOD
55qjCw57xEXAH85m+WBpy9AGHdhZFJZ8r7cBtp8QTwFRTTJbC81jcbE8aaliUIYA
QH223McSG2/HEEH+ZKuud0NPvvdBhdKTFxEjYCu4Gz0MJiMKkeG3imxLQTuxZp1s
m7qG0jRWq/lvVv3R3fLMMyPbzP+7LXUuSOfYv1UpFKalEg9eOq39WX66H2qUSC9D
XaLW1lNLh8pI4FHA2jddetfAptra17zuA2u5K8I5wGqwD5f7kUaohd5HrlYpo5ht
/+iORnA3MJZ2cFm1b/oPU4VfQiCC5ADiKN9+J66QNvROklzcRifkQDiKg5TjjEX/
fPH4Kt9xhn2cWNzr5+c0sEex3TyKu8VBh4GLyNBho2m3eefPMyVbiuaXdTUFg5/y
UJ306O2OVYFWLUNCjMi670k/4IRvoiwpQwuY1iCrRGdPCmBBP1HLAPlIEKs5JFGF
1WnkfzO0R0dyZibAgB/DXvjwy7pyjLqJ1jFi5StGEx0b/J8G2NKLRaVkOlYuoSoS
BrqbCQHRmTBvvolf3uKjzcfdDx2VX+mVFtbUyjWU/GzvVPLowyYFMhUE8AK1Uwsy
Luav5QgBdH7gO5Dc9C1c9U94vlPsM5iyhkswpgANadpiuzglHXx0/u7lfadii+ly
i9Xy9JwRtkPJn8Nk9DwUQdtbv5eJuvLa0DniDq6P2lTw4RS2YL0I3qB7QwBjnvki
xMULr6ckqUOdgkSlCyIUeaOGD6hV0jL3GiiV2mHH0ml4dAEFAt8uA+arVTb5yHFI
355QOdLYQZ4BfMSJdzSof6d77C1RXU9kYEVVlGzjf7dQtlnLBo9I/cmUwbyVQ3Up
bmtbjATXwhaUG2Ro0gZgYZZ47tYoNT9Lmw98Cb1TTRHG4R3O9KYDyyMbF6JjQ3ov
c5ujQqz5g/kBlrM8MSMQJzMyb7pm0CqyTnRC/2Xt6ibkmMlSOYRPNyyROGZ5YpwY
aPcoQPZu9eqCDfVVz8nQFtXbwFTafHUzWixeh5AVIGcVJaTw+8olA/sDANgRx8cT
MTwBJuqzS+XQjWHyJKG1GqJZHcHgmFdf9Wpw2ot2xbUVI0oG5P4CnhfVMN2+snka
+UdHV2D/AlQzu1Gw+zw/mp7XDDQyMriHj1F+8d3zZoG6sRCtk9Gh2kJEF4FUw15O
2eu3ARgyhNOAUMNHcj5WsswWzVFo5AvULCzcnCqflBs9GIm+73Z8/jVuqecWesO6
Hl4xBQa2Tl3V7cgoCjfctmW+bBopuMFSkTOEQqxc90DKAN7bO1mDXyC3DazocSgI
kEy2VhQ/iC/kzhPBIiGVMSn7ZYWqPbpoZSMHJUTmwCJsvtn1fIZlFMCyxBM3Q73J
XEFv87J6Wbahvt+ZX1pFjvJCHNwI6eh3Pxp6+dCmaUCwGxmhk1kgzsBgKG35BZhh
X2EAfhDpO2+C5O0WSCLiAPEbTuqjrNnygtk9UXqwFUbrTA564tWSiWGyugzCCbiT
WoY/PX/Gn4NkrAmmfg7EjZrz0CYIx5c9+iNiStBU/itXACtzUruAX28VquowpPBs
qmq9X0gjrVDI3mCk7T9QVzNv7v60feLA65OSf9FfZ3MiTNm9tj4+/8S5WJDAYCSY
SL7Mli0n9tF6sEv8iEZ1RI8BfTSuynWG9Jel75slJCfM56NyTgs5BcuJ9bzpZLcI
xeOIl22QLsluNAxVLIi7yk2JSElZFjYY5U8ixZwb4732HH6nLIBxqEbFj/HCLkqJ
H/0ZlRS5m6uQdPlaZrx2gcjjGBDZ00Y/Tz5XV5W/tBN/tX0vlUZ7qlB6agLSkk5v
pgVY++Dpsa7L/XJCcTx65qKxXRiQEmNQ9L1cg7UL0KHE/dCHfKXi/6nYgbtchZP5
5rrPGHqt/CICJZwwXneZJTCbbUiyWjANkBbE8XRGmlI3WPQ5dXFIL4bBQ3Gcx1xd
gnC0oGnHieeRu1GfZhEVQti5YS6mNGMBdhyHJSynS566s8GUMj4BNNG/99vh223v
4jrLD5AiRuKBsMFSN/5vIjThZxuDKXaSLNwOXr4FIYx39LtqMyK88lSr7F+k+1B8
VEvmGe29DaUpZpDDGftxUzPaxZrhaLLTuUlfMtd1616PsKfVo2Ai6qVHjbIKLAB+
X+AXhcioDiDvDqH8gj1w26PnyTKRy5Nc3HhM14+q68a2Tkj7t6cTe9Vr2EhnkbYL
oIi1/3sKvnOS4M0rgOfd5WNjnnm84ScI69yD66qRHxWiJzO0h0ZXDJbTvL0CCm1K
oFY6gGfCBcqLQsQ8dlzd/rs4LSzEVzm79cLxihpyAUkhXokaq+ZyZA2gnFRpR0kl
2BceDqWRDZ92vG374QhmfxmSWwsEoPRokQTOc6SQ42HKwe1nhzKjGD/xZcxpsjpc
iPOBgGQef5KBvyLUssFNntcZY8rLJP4U5Un7ToLHBI+37KT5y9jlBzbNsMqOVOoM
RXjH8qPgCoL+GqVj4Lyo/V8aneDbr7lRg+S7EhUOJqkSr1F81Q5LQiQsPLPiEghG
QAlqTQ3WQ69+v6PvjmMjRRAbyUqsXS00EoU5IAbSsKjYYf+KkuWXcWmLOG7Xd/Vr
Bgo9qQJLVPZYWgf15n0PaNmDTyOdfJ693MTiT5HQ3mkYrnaZt1Rkfgo4prc7KU1i
ZU3QFBqP0KiM+N2FEFe1JVxm/+1kRBsYFaBUFIc9zPw6GArgsoolWtebHSjb1xS3
ir+5jKw3lLIbWZFmEKcyQumCRaBP9rsws3tqOkEEpibs4JGyolW6aRWzA21rVuJa
MF2nFDfcmlRgf5W2gUy8SlBxXXz/JLdr9I1j+IRCKBEH9q4s/Lvu+iCkI4ltZPcr
RNor+wJVa+o6UU96ho8OkGqVRoXX0Bh3hmXqVrZBhq1Yln5Gc7EAgLACxCMbjbPO
vrJ8/F9QG/30MxM57PNQ5GLWrYbcAoSnUgsoV1drCcf8XyLU3qFJonoNThpiULnJ
pRsv6AaritD5y+nMAWaW91ggghsM53UFgR5qpD6xKEaEJ/KgKEg20xE0qXIF5rnT
imchEShFPgikUzhQX47eNvOARSl97IDwLI1bKRLYaWtHQlOly9tKYMJKwvTcLOD3
XZM/dlxpTSElAUy4b0dypSTPP7Ogd9u7rAdNX1AHe19jWB3/na3NGGLOp0F48IEF
eXopK3FQ6uvKpfVmO4mdLfXRwXBFbuffekA572PXY5eMTPtu6ELKfud8/WSaDNj9
W1DkotTnCtEaB2savFb5FppyTyExF8RmRIE3wXWEjY4rsDETKI1am+8pq+evT5zj
QjEWTiwDbuBCkDLRV9dQCTXepmHa6pwny/gGy8/kgKc+6uKNrYgL7dQD6gMftfHy
mCd/HWbvLoUnVgNIcwi04ZGD4qhBQbsetS3ig3cEY6oujhiFM4towYfBWVPDy4to
u2J2sjj6dGiKglKggHJ/N6493j6hyOCdb5WiDWyzs2gfTbVK6FX1+QKlRoPeId8V
nQWUlnIkV2Mv7uzZNHjMQrAUUHwTpNd3vWwNUx3AFuSCACJJCUbyU9adulYlIrgR
cBUmro8k1WCjiGxQHlh6yp6AwaWgYsQTKFs3gq6c9EKqAHYx4FG/EWCI455V6NRo
K2Df47gqZteicKMvLYWAtUvy4JZwBtGugJlBvknafw4FUemWAwWrTInuX4UyWXEb
5Iu1GLj1mruPxUaWs+q4G8gScqxjVJZBES2GcXhYpnuQF8xHnEeWyB4kfVJak1ka
OnAVKMjtUsgHsw6CswVSJ0OTIxdD878t5lKx2Uc28VwiR/uTy8dGZGPfs4cN8JFh
9rjpcwoQ3dPF/kdOauddqXIMWL/3rV3vfn+NISfelLP6ZYy52sxqByHHCdhiYt+3
UGGPIOOTe8rMAUGzHduA3sKxrhTSx1gMTwcxwFzq4qUTtE4thjlZfDL1v3f2nz3O
jXT2gT2o8DGmIuIZdAqt7NiHoda9xUIqehCfki9i7Yg5a6DkcVLBIrVrZBV9tRt0
y8c9z89AVkJGl8HMSlsrYfI90OoSJiMHQfvT//5wpgmTJ5sR7KkKad3NIfWPu0hc
yWNKLYwE2zwZAGhjWAXGm7b7i73zfan2XkXCbAkct6MksHy4esWFKdhyvKsRmRuJ
nRfbuvYwM6/UmraEYd/SFzCRYN0TwpRvLJu4Oo9/QicogiXgSVEb1b5KJonvLpDs
TNWKuknL4fDGg2eFvbQwSrxWeABLQtqdRGYe1wwEX+uiAFpZ9p+nDUnv2ytkxeSY
2QDttAXSX50O96FMku/6hBR+jYfusuQKCGQCi+VdqeyucaPv1ocfpuAgyyJz/gIX
nMXX0KVrdOlAUAnckgipXSUbZEKGidFSV+oafR5ghmRRUZ/DgvZ1XVrGrHelK6K/
xRnWlMMB4es1Fsk9nl0uqGvH3H42hk5ugyuWM+4/dY0hSNoehwXHjKAZCEurctpg
SH3VzozLxHxmr2VpgwAqG62y463a76oHIey/h9xgpg+0wE39EeLcinPDWmZf6V+q
MHT9pj7Mnjdbqljgs/OUZGkPz7HJYOYMZ5IRbrDf7YbHz9HBwdzLi2Lj38uUVDPm
4kBhcMnCXlw1DIVSfnHw4fbxQsfaeE3On1vrPveGq8NXCLpvyeET04OeY9Fwx5r2
yZP1T6/M8Br7hq6wrE76FXuOc9EuVi5EvszEZWve1ywYOnlue4wAr/VaUWB4o8Nq
pl3IW3e0dkphdLxHADuddkzYzlVqtqFV+VAiX4AnLTZ4sSXprk5fYHWK8+lbLCrC
Nm5ZMwBAuTaZCIj2BJZtPzlpUH2dNn0XCVLl1mQV5+agpopSk45YulHvQyM1ZrCC
J/5oF7JV54IzZWoTqyvqAWvyotSS2TNFHFI9JI73XlOrlxcwZfNVhCZUji7ZmSL8
n1VVYO8g6t1jMxeKIStGSvGIxe9yaEBEe65HxOeRcRBGixlfx9CZLW2eek61+4uS
AyU8PorA+442wolyE570Xb1+I5RTkkAGJbt9G+7c6adaVJr8LEefrwMArWH6ZUdd
mTg92jBHh1LAEsUYDj0CXgPw1YsqhsmyI2UFh6LQkdD78gE2s3EVN/3bFaJD/V5N
rdhhnAPHNOTDQZNf1slZQBE/7sQ18CIZO/uB5I49N1z0e+qKUBJdmm58bCKALMZe
iVueVe9k7z7EGm3QP5rEteDB/A6P/R22rbtThDHqx13BjAS+SvVwBpM6rBLIbjA/
z0UINv7Mq2RqZKYqPpfepruFiF8MzT1p18wlY6WvvS7vWskf+7SNY2EIJ2T0+0f7
FXuZ8dlfq0Hrv2aOzkVkIQjel438ujxyCHmUB51oBRANP0/xtG7fj1LKEt85lWHq
RjXQWVaI3zFxsjfXBUYZFN6okHQYddc2X35GMVR99hW1wSJWlIreCchnp/7HpoYw
+81LQCKeoSJW/U8msJMm8Up36HTcbRNpyZKHe/Baj7RucWY5LYwMOoO2y5eUPopq
ho7CcE3mNUU7wujl5ii/trDV8j46axQDr6FTlxulxka8YKxzyw0MymMK3J9oXEed
/yYE2LzYw8SVphNIvXt6erDVSfWn1mvH45A4ufyk+AYPrbMYn8TNFsbQb23bLlFE
Jh9gziPFsX0RxkrRmAwpn10MONry+9gwizuPfglTrj7FP/XSlChh7ck0wn85yaHP
/sKFzfVVMbbLlIOqWnRKsuWlz0XrqSFiPyJf/HeEppzR97t1FVMaJYB07KWOhTLF
DydhD8iU6fN2+3wW2GMi8xxjpkNZrTGBx6aoJ4jtGhS62oGj+LTBSVDHrj+oIild
QQLrBAXHmqrRTHgcm11Ds6pK64b0OYYRLPGV2onIIUF8O0O1rZg9M6/CAyVBd4qz
ELHe4faziEik0aY7kH6HhpQPCeZ2iAbvUVJnraGbfzy/55lgemBn1Rpc2HuzpqeL
1jEtzIsMbXON4guPyj4/Lkro7Vw/rf0NBdT1/ZwTksVyiQkLvt3oG+jloCAjA9kB
H1Mf0hqWLpE7omuu4hUJFxEbEj8g1y42BY+VLeVUKapbPpHatQ6HcHiSgsxoit8T
6tL/w4kL3RZ9xaN+sjwkLrj3Tx0PfMV+4vjCODMVV/gzRRw7chGzo9H1Z1kEPtRK
Cuar7yjxprJOW0sh+m3WlEDQCE6Pa5IkTOe6VBJnFr4/bP+5KFwNvTanI4QJMn1d
eGt3blQfEugE96wlDTI4r4yJfRaJ0m03lbCypVvXmwYlDVZ3WgtXT6HftVjScq9N
8Rtex0HiJPxDCQoM+lDn82W2S1ARH9NL/XV2CH6zvBsC0uP+RTXxfnPBNJsVzYeu
y2rPJFL6Y4hYVOjXy0Nc0aMAJmD3K3wL+wx6XAYRTfu9uqsR7PuNVpOhvtDbY2/R
2cecg1KRzPX92FoH/Og1KYqiBXzuT0VZ1a4MkZlUJuYtIlYpi1gjYPAECIKyG1rO
EqTRkWUZG6fiWgch9vcDodUoip+12wlATFiFgp3JVDDOXguVeZ8wkJbhXN5SHcv2
uSvFG6VtzovIqxgG7nYS85MuvD6VN1e4RTR3R1Dk/p8J4Wu7NaBT+77/q5onxN17
L/CT/YelVdQX8ERMdN4PNDSVdufXhoR161VpALXLH0CwjoAg96K8vmgysNmgLp2k
c2cAIfPktSMV2xqWCHr//h5iigP49gNquT5ER89kJyaNzUsO53bzHzbHyEYu+RrA
I9GHpyHXI4+4+jKAywwtrKTwsoxs4RrMe/L4BXJr74x1fQwfyHW7bYqCvz3K6LT8
g6+bAPZHuQN1Mn63EPcYRoJp/KWIu5IDiL4SHb0QtbSM9L0KE24k5W9o5QIm/SDV
kIevdH5L0GgpDxHgMIno3H7tZYVX40thcqYfw93BcNXG5Guf7jpXvh5YBdDe0R/+
3tNu9C33NjaDAXZ/Nmm92P9E4KGSaz8HlrNuL8cw+MMC+HYEL3EFP8T+L3nxY/s1
x0t3kFOBcxnGKLuKv4yRTMdRDOueQq5B4a4iAuGAL5eJAR0Ma3hRB+9dNHUdAOMb
2+aab1FrLmy3ubBzEpZXrcNZinMoVDNEuEm5UZfBrJFF6vS3Ien7qN+sEGusjDay
UB/cf3ElBLkwe8GoDolqg2xXrnNDAl1vqn/YFasj8RI+3/1EH/EfG3HzcDNRtVwL
jbp3p2Px/d6Fg1vpRSM0ziqo1CJI8O35hzt4iyOd/CvMhZOBnuDhbtDRug7wyNhS
AguGut4VDerr6u3mByG2tHBKUikN07xHYFVCOkj8jfuhfzR1HbNSb9LOH68SZJnl
3TE7M5NGWL4gk2h+V0R/ma2Oevah6jXgaCJLwXXftucgS6RE7cZwwhbKmmwle8ey
tCtfLvqpCujD+WuOHOqqb0FuvHpik0fS7R2psVFGfz66/Uqi65wnL6/Jfkfzdy0e
KlLgdygj8YtXjJT2fDZ233YHkM3yM17JQ+QDvAA6NGJtANJTb+H64tMJrBPqERU+
eYTwmpkNoeuOUbCA5EdOELYO3IQRg3ToLPhqjZVH41Vb9Wttu0kOlXdTx5oPRRYx
9mR+kfvXncnzXn8PLgPN6b83y0pSa403wlARLf/4FObUBZWc1KYr0CFaBZFCIP8M
wsg0xPczQu2tMbDs4s5fOZa950v7w4DtIA/dt2YSt03+eM4wxob9cy400cGvZF2n
koMLnIZEDHXW9hJAb7ffChu7dUZFPW3APWOL/rcRxWkt0Mz0xRVykSWKXd2AybBP
Mqd9DAClcz5QWEywUvXDNkDikm+M3yJldX3hRYheZ5cE4fkf51zSlGJZ3X+P2WDm
aiic8RY6xUtH1NYafp9SQhKidE8+HRFxH7iXiM1iZRKyQ/nHu85hQxV4b3H2o0Fm
iHoSWkHMcMao82LgXUSJwMImLp3IgQIphleXZXVh3XjHD0HhOywONjTvcn5L29Rz
zdXGh/PpkNHF5Ya8p7zeF2kw98G48kxWIF/n1cFVYsMoxCbLYeEgJX3BNuq+q88A
MSWQzaBUgOwp6MaBGT2NeTKPjZ0wH+R1czvd1PpnYb+lu80/uUbk+C+zDhBrfxcj
w5DDz8hm1BrSTukUXpVMM/nkc1MNaYLjV93w7OK6bgSCk+hL8MOmHBrnTIAPrbuh
EcFZJaj7OzIlYxExShvpXSS2lxoQGtWWnjP3Sr5NkzJnx4Wxsdk46cg+Cj7AH6X/
cNHo3eDUVVHaJ7TFAB+KmzooCYYwSFWqavv5oMVSz/LHsYnXPHLobSk/Js9+z3/w
4vGxUN1RRDqtU6KNbeI60BQeYgs+8zjPNFngB51iOweu0MxjlgM8ifkRKZRQbRdd
XrXiwb657PsMQVyAbtcrOOdikZklAbwUhCPoj3krtCseqx515wN3oZB6cwvhmhpk
HzfxXwG2GYQ12woVBhkPU2/Ak+u3tmBmNEdJLKvkh7KIXMF0DLG/mZyVljm/158J
p46GCXrDBtyzLmNy2M4wNHlwXzuesV90HM8ZDJ4xuXEEWee7V4JKgB+VetVSPJNQ
ohzJS8XMopcoh3jKqDMzeB9HhQ2s5ckaxPOnjdTgtfDPVKt3GGT4Dkp272HIOpgU
ZDdy6PDTUVXRNA1pqQyFGXnFvLUsKIVTcDbvRmEKQOKnpKV0Hkx0dttV/rBdR8iy
2LZdKrGOQGsqSxRqhyikses33wriz6ZQek2cysaopxAWyGofwGBt4st/8F/Ga/au
g2Z8IoEHoJ+Bj3+humd11eayZcQdhxs7uTzfkeZjVs4X6fJYAg30/RxCM9E53Dt4
p77RrhePlyM5/SpZPW4fwXvrz7eNk3y5NzdsAy8+Ek6nBVH6aTOTBBlJKJqlD3Y0
JMRWI22BJf5HN0BozPH9Cbt4fgt/hvqctgxvIExJXelGjKRk21N1xeJrtueeoVwh
Js7GOiE+B/Z6FkTnM70nbMJ3RALdFAw5zOLJwd+A75E/ceUciTJaDpG8KWpOmeBB
0RN8mHfijEuVB0Tw529jvWR2WIqgwhnAsVyUaHmGLjg2qDTQZDvhNdz3Gzy4bffu
cwWCFKpyqY1ZAnCYf1gt/5rYNhjrSq/TFMbdzc9U7MSxBf5hj140ccy26NO7aOa+
TpHekYBC6I6D+wqsGMslNglS963amQaUENvMB7tjOIrVmFKKthjckK7XdpBdzBca
SOY/NsCeKE8BvSmWhDJw0lLXE369gUBDAU51BgvH1t1HrFyHdnTw9rGmULzeI5Bg
fpmEEKoLgIwoWC/aNRdEQs1nfPUeH9UaPwVayMhOYMXif5UAXeAQbxlMKwCsjocD
qA9KH5Aq46p5X2PmdppvOtcUEQ2uiCQ0mkEJvrhUGDg+GDsATGL8wArqusdwb0WY
sXOR9keNSceDwRN+jXLJXsPIQx8Gnf7azjeOFbLJ9ouc/ICx88bMEl+NVkKM8ZIB
dXq5CdIbIgRacCbtjYJBsADJzNC3b8UGgUdNuWRzdVRtEHo4OpATwL7t0/n+ZTTW
U/d3BMRkLY+en5raMBdJ9TNHvvZ1SQtC7/HoxeahV7Y+Bs6ECQ6McTlm43hW0cF3
3XikDH/6Zvif0DtxrVTfBywqNlN75D2pQKc3ArwgieOQrBpdh5dOfyw1BAD4FKcO
WaJ6U8UW0mBMuauktlqhJTKctBR7o7CMjJi4+xX86K8v8vpc6moOes4oA1twXJfC
a8BJKGzOZSQwACCUWCHwK2ToqO/sphp/qKAYxo0NI0+jezJ/LiyGAxBPaYhTfNac
/uhl+7osK17Ew/N2jHWdZ1q0oqP91G7OEAhKdUMG1Oi2FpMmd95/NyYXa7xSlBPF
67C8+TRKY14cSqV8EUi+PN6iIIE9J3t+FiBAaBxysKv1g8If2Rop/SXJ+ZXMlik8
4Cuf91/j7ZYtMn+3y2SbuJYw6kj46Ej+295CWOj0NFpcyKK1pkUz5VqHT5h+EbsD
p5VIGsOFABvgtpqjYDN/oqd1wfb1LD2+xlu9CHMgOBUmRtpNRy2SwXzAiT3GdDYS
xJMcwcyHV48j3znz9lNmrj2w5sn4To90nbq9PcptUcpwzDd+UzbQLVr5kpcZhvGr
oDdDT0RkArpdput5Vk1dj+5ILFTancOB2ZWqP2fn+jE5N8omMTMzbqID7vbv1Ghh
irC+BzyC/ADXTiZ/WoIZQrnlQn4rAuq0CAGz1oxpa/+Rim77MlJjKbw/jJZDBGpJ
mCjpdWJ9AEoGzIYGxxHt/mF75tT2FhB7buIzTfaDszcx5yw9y8rbqA6p408ZVwGQ
m2fo9h4EnweLJq4YbPiFVZIKwGOAngd7jD2wQtmrsViR3rY290zVxeEKUQVlW12Z
veboudyKlIApv0+Z0TOHdepeg9V9fXxqTDEpfnq8Opv2nwlg5I7SkMhEqWkZvq2a
BjJHF/ftxd05pCHW86VESZ7+SsG2Pe/JAD0aYZ3KZ0XEjDZPydUByuUxvRiXUgUO
eUtLzQmRxP8SkAZKOYcp0uFGeM4E6innYZduYjfNut6tK0o+E7+XDQt+DRrstH5n
X114P8VJ/EBiY7ZLBEwkC6ZLTDkSfuthnzMQtiyWoKd+GHSX30nTVp3DOUl/7z9F
QTBX6eYy5s2214lsk9Xphj+uIWUAC44TW+/GNoqX9vK/mLQhvPrRQykZ07B3n48o
84eDvrkvR5C40KsM1aJDrBCqNon60vFh/Aox+0CQHn5BfBmFDvKIPshLdKl2RfUL
SyR6BunaXELpACpzVI0tUd/iq7kD0FEL+ovKD+jVbiGwjAdnmBsloTfXCKf61VmV
3KgCgFcN3SysqtQXCdIFxaApAVbdbIG/TvF5nB3Yajzb6q3F+eoTsohXpiK/gxzE
BSCecm8aLNaswhAxK1aejUrHrk4Jq00G70lk+iEnZ5fTJMj2Q/VzIcZ9roFzlJ9j
e2Lh5H7okqVEcJjmkxjKnEWHsSHoSZf7HsfLBr8zPNxPT8QFysKrIwflK1By1OQZ
q/GSfhC9MuRcheus3aPO2fqSfjDd5e4XPPfyWhLJ7CRle8P5KEG7ECa+um+DGzYF
knouaIY7KBMuGnncok9NOpu7n2xzN7uCplhsmgvmLL3jdD62ZXdqkFjBls3nrc+K
jDgsXCV2XDdfXwq5RtUoqhE+3emlv1FEdcid3dsOdWj2AUxEITS1sMilGGhuh06l
Bhc0BVQy/R64tWNRJihSN1ZBtt8aAFCqnLopg4BL1ujolVgYxQZhy3kTy4NbVVbJ
/SLBnZGODf0rClvVR6hezKtz80szvubvWgVjw9PC4Jl5TLBimNUjGpPyZDGG4+rW
mnB1v33Ys39iBxcCoQmJDIaiNbMPma1Hd7i7+qAKcWZuOTRGeRk83/S3j/Fge9vT
NvzpQN6A8LUDs/pDN7+mkKc0AOdC7vEsH4bvGpR5aI0Lz+btvjqi1Hz5Uw/WA0sc
PnaIa9GmjpvfReLF/HjBiaLq97fRHUVFu7z3ZwF4U23DuEn1wxejXprtdnlgaGGT
WKzH9hOjG4iYHrtN+hpsFfVeaRDQbccc4JNS47Kw24Rmj7+sc9PMFFZLBlgkCuRh
BDD1oxW0ow0ZjbEN5IC2Gos7hRMsft0ssl5Pxudm9HVk0LUaYX6RZfqhcMNobqc3
AGlhqYo2JHdxIUEUqkOzHAHwDH4LiF+xGHH0ZaqUA7OGzkSS7BXmwM/XeoF+kwve
FZlHBryhZaMRCgYF99qPe+skEWW1E35sWHcEpBb4XNmMeN0bNgV9E9vAYSEyT1gD
0H29a6A2LQG7r3WRZMr3K2spI51Q9FTK+Lnjg5UkGGyBI9rc0dZL9MJ655UPA6Fc
4rmzhSbcPi8+7PKk23Qfr0ZYGUNyJeRYBOi80VLP3GYPpIRjblxsPihVUVgezIaB
G6bbzaoCzHCxASINlyap6yDB6gRsYuo7qHG7Mp9/dADVd4Nl1TtrTcZUpTRVB9lG
htVn3qCzJT69mJeVIFgLIX+ZKD8LHlYiMLNDCLsxYLR/N6XJ4N8+0P+CTYKE7vn3
iQFZOuqqx7cUXKCNK33u5G3lukoLnuvH+uSxNfd+pvvqddRLAzqfRfydl+1nWE18
FQb5r9JQqXiMCXIQ6hYF6pK6pcLsAd/bCb/iggW0QkMeNKpadYMZDInU51CKkr3h
fa78WRNXr0zUdqC2AyjqgwLx61/QkPLupoYV2q1VhmlS5VyZSqxkpkrM3qSnx9a4
ZbCkaD0cTsNgljLqNTFqHcEPNxprZoHrggADCBu7++RrpgBJowYDFMKM4UR0g5JB
O7G5aWD3//mmGCi4MwpQ4pHPrxjsyDn7qed599mAbwN1TdfsOT4ZLpAmvciIrw0R
ifBb5MK83GaVlRYZSdLE3k3+Pq8lGur/mbZkXRZe6vPv7iDK8JHQT/No0NCdEq0I
TBL1yBzOQpM/GAFvbnMbDsRYZJhDEADT6oImecH1/Opy0GBOoey2z6RyBDUh0RHV
BQQbYtNMLRM0CyfXFQcMuzhG6yOZQcRKQjDYq9VajtXB63hFNMTDeQsPthLZD1i3
nJhqRmGwWnkwXnpjnqPzI71BQVGRfQd+T2LnO0uxZoZgLqI/+HDc6RQYvDXe0Gc1
YoUDAgtirjHUuWs11dLCW3+6VN3Q5fwcV8jMCLfxiwUTN2UJIWOjDeO6lSg+aTTM
1FiAKBauEOnUfbwKTD0sM9gaXquft3NnV4g2B0pGJbue4V/uI0e7GfGQVwqPDnLy
VKbN5qUNxPlMeT8+fnruONaFb4+gPg8Qr4FsEpJ5I5KkX1sNYOg2WsC5yy+n/nZL
FfUqlZbH5y2AO2GnlvNu54vEkE4yxQbvDi5wKtjCLnWvtSNI+d1ZUnCbJeKiHUdS
joOxLQzsw6tbTAETZtvu5mQ3g1tTohr61Wdj8q/mTqcitL0oLaIRvDLuhhf4mY29
QjRVlWaohabKwu0rba7+FgNGSkeerh8Rpm3GwvukIqO7OfPX5j4VcVPrcZrGBO3H
Cx++z9yAtUR5bTEaU0UgmdblQpgsWplxmvnSONHQeQA5VBZPJJiAoUgqxH5ex52f
8p9XT1KOQ9sqmfRP5N0Q6tSrjl8piGupVJpoyxbBF1m2weQvuOnSt+ajSjku79YY
0hxuFpaBqEcfPzvQseLVU0r1Yw8HIjaP4hj+6cYldtbzEmEPHr0/v4HVX0bx66eC
MeCMRYO4/vlrLcUT0C6Ew43bZY7sF141CsZo6vyfZ3PqZ3PsfAM4XfHiLJpm3CkP
vXccUTMQYcgEek0PbUhLd3JLj/3jUE7Rnll5E4k2ogWXtNNUQ27FCGaN1l5tvT7A
Aaa3P/0ArTAiu+V1errnoHlpigJ/y57tldna/Dx78qZGmQ3IvdJk4Yy9Fs/GadTo
h328vxvu/bIeDopnZWjrLVmLe3aYq7Ocxyt8t6uk+5B+UteFTtiJ+LzmuROrZiaV
GWlf8aKw6/QRDAbjitw0/6sOmjeBrhMm9FEq6zk2B+44skLTKJ0DUHZH3L/TjE3a
8JyQxlv4h8ALFrRHEdPfg8PwKYNOgjzoiO90hdtCB9lcqaZqJij9ZS5nhxyDvaBP
7qQUDUFfa1Q3fM+Ph1345aWMyr3Qv6eXgBmqb/g8MKqQsqp9Zt96/+riU3/rrNNE
NsDdgjNr6xIk1Gko1RqmX+YaBoydp7HSxYgZq6fE5XYw23xarMjH+s4TKLkYEXw9
RZ75eTf4tulpvLWcWd6MDrecFsbfeYLXEH1DcJDMl6qZSFsWHY5WqPJJJG+KgyEY
+83TrvSEIUgIM7KyBVAH4cXIkMg+n4tLstP2zjJ4yEmGrpUO45WWtkPEBvuiX+02
cewtCgPSfKh1G1I3LoeUdeI/3Yvfp0HaQPc9xHtXeSQ8qXrrNCL97gWC/5lfgVlu
IIXmm0WL76MAGhxuxf8v63bFTNuscm0xfgeK0Ez9F0sdtkwx5xy4uPrfJHWvvW5R
CcBkNIzgd2hzf5+fkGPxXPWzn8+skFfHbwW0bpwAcb0wAdtPKhiEMB/ancWGXdDy
jsoi+jfJfKX5sC8x1JHwK8MWN4X1EreUu3G4tyjIsON3KyQG+ZP63iHfrZTtvChz
WsmlJYxOXtfaChhsHHeIFroSmw2IhqkE/LHupmGKigVl1jkOgDzgHFTygE7mb6s3
vhbavtVusZxY+PBDlq18d2MgQUjlfuJYAFgW2vm5f682g4FOlb87CrrXhx0V/akL
Nod1WBCD9dzQLzHDDIWY8hl0kfwp5gL5yxUNA26kdqci9pv3O1/eegLNTJskrbsc
NFxH/Z2Dlv/iee6+PToGAYwbB+c2Xq7910WbUlGOT1qssKzgmcKagYibKaRrfQMi
OXLKmAm4N9iCEjPnfFPJyHApuQzksXyE+S1F68lrLbI9CvwxQq4pfKR7OwxcbqN/
kPdlBtD3RaWM9+bs7aJZyu4WS979331NLjY213UmaJM6qwYDLBcdHU201eg3aNUp
Blz/PGhoi5rcKp3+C5Ig2yz5AaRZ6g00yJ9xii3ajQAhcajJ2MAdYLcQJQp7WyMC
fzlb9dYmPcwkce8ZnKR/hyDBabomLlvPWHKLCPjQd+9+YOEiy0atPYil+1VeGqh/
ruXGxcr4eXmjctHKxinL0l97nIMArqMLDAbcEbMjbzQNraftb4fSPvTlYj3s9E2x
ft4GUoI9FTCYIZ/7Ab6vChoMZkoVNubYmFMVIf1RV9XRUvjNTHRH8EPDUt2yDu0J
S1wbxtaiJYvIF5QExJUw+vnizsUVIxCZTnUNWZAS9OBUbPLBfxD34QWl3NN1XaFB
VRaRbvI7G5W15gY1P1quwwv5UclNvRQurOeXPVRjQqCDidQnoiZuWTO9WVfL+dOL
kJLlteLwJiOnEXCbkdGkcUK3w7BFIK1c6e25CGombq5sPkjipVFO5pCvETRY5SfD
/qHHwb8IDBh7yaCw+0EyWUTGNBuPY3g8scI1ggGe8/wFKnVE/XUEbnmeLuISJzqb
Wj4b0WGbqKm/6oN0E9ZbqmpKSiuKuWE07YPoQg0uUN83wzfm0Vd1ZrOzMSVE1g6M
i8qq2yfKUiBP4p34ZdJf0Il3yRQJ7L/ZKTRvSZ5eBFztAmTO2bu9yaeEwzwbAvlN
Mbg+BOJGSAihn/5/gtBpMOd9UnFVb97rs8zDSiKLDxPVkHU4BO2ombM6jYzzrHlA
T6WiORsrEamt4FVF5mWNy5ADV2LosjHfOuF6mopWbSB8aPiorpR5Np1pNEIcOaU7
RKLRV28sTAqhcEkl0L20m7X1lT0+mh9NIIYpqSpXiPQ2Zg85KgRICDvjKNkci7tW
bIT053vqKbjVr8grM5pWbZ7CVaT08l6c03dIiH0hOVBijdkyL6psSnnK8bdJtgUf
A5dEG8g8MT3IdJoFIT2zSIcDOYUI+cbkaFf2z6Mvj7+/IxaAGiy/PWPbNLviuVQw
v2RLQlXsllYlIdeeeO8cX9fDTQpMP8wOjX+hWblEXwfKp9rDM024WS3gh0apA3Sf
norlP1q+03N+e7Rh4ETMET565A9mmRgiZ1J+JtPOMSTAxVU/KA1CRFIYjhDU2tss
ZEtEfufe5N7vcySg3trdk6w3ZoPcxcbEZaClfA4D3xskQB64WSDpln4ujqaOgB3W
kiHXnkfo/1Dbg9p8mlkoe32pZ1der8Xk5Uqb6vh4Iex45CEsHVqAI2che4Ewmgbc
7f7VLS5Gnnfinglw3tL0DuO6eIMdt9YwgB4AlJUMxfT63c8b/z0xKnAaXbEZqXvQ
vX1Yqj93U0GbN6VwzZG6sjIQ8b+Ukt1i7j3VBXiporj4NsS6jfxcL91iSBlW+oVQ
iTHZZ0FsWjY+On7VYB0xPCnYZXPH80i7H8PapZBnt1njZvnER56pOMkYf12O1fND
oxsvw7BtrBCyPmtnegW1X3uQk3+PIhoT/by/d1GORp50jlSC/WofxQDykBKP3nWt
uq6p8WXSNqb/0GQE80BQjVOfPlZpHnKNRmKusnMWM94Cz/W26jjYuy/Mbz2ybZVQ
lEe5juZOWQDNswsHdX6YxXD3/zNJQ+q4bwdrVbqtCVlzWra7mDBjFk5fvcgYsTI7
tGwRZFd5Ee/60fv/ABMJUwDRfylW9rg6j0hXoq6pTRMsfhocaWQvWVS56ZHuUaxA
UHVnzQj69Bn07mwVrO1MJYzO6GkwAY8EI4Xs02Wr/sYRkKQU39VBHi8TTOpNvR+B
N2xa1sWgs3LEAKQFhGjTy/gxadTRW/xDbey5sLtaqTJeiFcXGDbxd8GK3Hh5X9Xd
KxSiEz6ussj7ND3l86alRlmcWuYWl20dB1xTv/YyHtEwytq8gkNb0OzQ/e7xLMDP
vhKgR5kJizG2B6zFio2NULaCrwRp//C7GAdb6yNaRbyU94uRsmeANxHEpse3euhv
IP6ypAOIA1x5ic1+QiGBPuOagxafKiDQ+rKC1we08EvAVTI4SfB2AdHcoWOQ4Hw8
XqY9BkF3xVBFwoIhFce9eT0PBHG2vL3orjfjkk8+t5ddlS40DdmY+jxpU5RodWBF
Ay3C8JwdfYy3jOT2u8r+RVkzLsQgvYJT6k3oKt93wUUOy79DLrEGZxlKQXPGFFf0
K+L2NX/M8LEtAM1SYPIseHbl9LkEd3hCXrMOJto8hbEkcQFf1ctBghPhm2bp9INd
iciyS6H9MrL4vDikHIIEt9WighwJny3tNnjFjLm31n9oNdklbBsz3WrY26ApbNsm
uYQGq4W3T9NaaIOxza2fSUR05bxCIiTl0wyzz5MilLAnhcWkDENqlxa6vHWb6sDX
ASDP1y1pIVZ+zOqC7CP/E1wT6cfX5q5vyGLHpQI4dm7iWK/axhUG+o+oVOqV2z1O
wTFQGWvXJrCPrKRVAyBYY58ZXegTlQfqEnHlrO1kNMbF1Bxd3GO2YneQa9dFTg51
fXpR+BlHsLFPZM+RQfZGGYWrFBzXzHczwML/cEaspFZU0ImHOfbI6O7YqMTJ8OjJ
15V+xZGAaWrNjBF1bjdI3F2TjVWHlgj7JRXn/uDwjyy9rUnFuz0W4UnJ5Mbj/t/u
goBGTGoXc06zGuu/3zDeBgvUuN4EVXBCwgFYw/sK8uaazLwSaWXSLOHcE99BaNdc
CINO1CTekY8ncFBHUfVBOghWrP+xbrw8P4rhiFrDblriQ5Ep906zP9Z3Uh7ps+Wn
5Qv+L3IkJ8pvcwydq7zgmQq50vAdVPVc9Jdc10xxCTGppWcCAH0eQhCzY55mzoZd
pTHWcsj9nE4hVQfDO5vWJUPyDPXTyPtKs5N6oxmlcorRoARY+id50tBA6Z4+mGwJ
fVNhkpjipxBkXxJTK92q9OMdQ1zDSYdm5Ow1xIlMOcYnw9y0s/CA4Avl38NxTG3i
UoxbeuHhK+bfa2LPHlpdvt2/C0xir5Yt4dyhBt+6FCLwn1GpB43/yfIb56gaD3ue
hZi2O0Io164cBgDtjQrgh5DQ82x02xdrbIHtHUC+ztY+pDLORMSKb4GbFOCzOnGt
yqOkpbQKrtmFtHWxDHBiF2qyEJ8D2SjUuFeT4bjeBSmFIqUqsySOu27JNIWKQ0vf
zBmxNSVqpuHD81Ab7Q1N6oQAyWIJC2f/YhqBBrquOX8deWEKnKQ4MyprkqT03bBF
GFZ3wwpEtywi+QhVahZ7KLveC27EUoahci767otOAqMIyo8NigLqetlI9CBc4ej5
JsFADqXx3ZwrWQjeFcFZ6ahdwcVucbJOjLO34jHQdFKm3yqH2L0rgy/RDiIUue0o
oudnIqJt5dP2l8MbcuE+ACuWile6U+YkHb16H1CF8vRj+O++WNt9Px3L4482RIkV
bRNZ4FbhTqj2nJV54/+ot6cs5YCJuqQ2Gt4T1ZrW/ZNdoOFCWBQ9gHhPF0BFqCFO
z0scrUkzbf6ijkO2LnVxlMnRhoX/Q5UV+Dwku8juG5PPKnDkHCpmANUenBWBxlJq
TyZh4yv0Do9FBMB86TG6q9J/uy8U38juRIHyQMEvXNkp+G9SBCM4HjTbUc7DDrP+
MrNQYUPTwEgK2UDQxGX2jaihLpbMPTfBtaC36HMYqSg75USiSWdyQYQkyZb8x8IS
pEh+jfgsc9oPbSvMf7rTaPsJgvbtdCkxvycp+ZpZfo1gOU9P3u7JUWApm4vl2CbQ
xNrO7O9n1SkJNyhBjt2t+huCb4g4weh9tOw0T/OMvkeT8IL4kpT7h+4MEkk81SEz
/K/tZxRvY5B3PH0tvtx2YYFZIOhvmZtK9liZqI5n6QFOepW5e1o+JXJDDKKxIrxh
vnq9oLHil4JIK4+xn5RHymauscJ2TPBvu4c0fpZZUDoQExcdRhAM2XYAeS7AeSMV
WmU+FuhAFDBECcTQbyY8ljdNvG4zzHilt0AIPa63tCUnvp8Zw1nLoUj1qIiLOLUb
S9vGr50OuPMhZPtQZb8cCmuq6foN2b61gMbsWcRFsANJNMG7y/STc5OuHXtW2C6x
ifGR3ZiyPIc0ZHIMjdidphbV0O5RWkF9UaFowEBEqPmi9zXWYlSIztmbgwF2Dh7a
xpWblQWP2goy0UkhKEuk91p3xLppFfDdKrsgZFUc9Ac/o6UnYa66Hi2lFZ9gadEx
A4nLQWs1hqBpl9Y7O0W0aaa4ItA1c+B9N1/e+GzhDQ0ugfSB2Ahs3dBH6pYjbs6D
1xqqJzPM4Rk5nXEBHOe/8IO+PWGZT0bPbF3wyJr9w1eUSL8A/sTOvonM0wyxhhse
Q8Dk/6sZmpmR+LNZsTjrkVTzmMoHB9zgYiFx8a6A3QAdyn4uz2eLB8WyN78D5JHc
DFSf4yPAUJ9HjqbnhRY6x8A3uDx9rm6LBCg3JTQBkJZvIrpJp76NxDtq1a93aOHS
y5If68+QH7tJ8MZDKwznzKIigJ/pyh3zYTANMwmmAdRqhQXP5juPjZ7NLH/T4vKL
mPTB+8ItAw3DtW8yj6mc0Yaxhf2ZzFNBx/7jJpx1cgM0e4D4GNrOFVEeHCPa8ijH
NBwBbXeTY2WXYjdhDYGsHUnqq7BpgPkGdTjzdHRHMGhFuNmN9HYNjUQR7JBcH8sU
s3zpCjVR34jQhWsUQsDf8yB+UjmxHxFJBXl/cY6usl82bi8HUIvhZGK0GIMnmHze
c8l/ij6nvI3iToSxK4I8QFDwQP5TyGRxkS/CKQArpWnIgtxRUWyo77UmXy4+TkbS
GDTdeCbGCN10HvBEC8VnLuTdmGUd1O8ST1nGX4XPkiUdMDWStIL/5C0stocMUu3A
CdHZfCPsJzjVMNzG81UnJ2s4ygBbv1T2Sm12643vY2hIYzZ+YsIq0i7rTDT9Ry5b
Y9rHjMtxjliSnbsSeTcJI/NKBOUqUhHN1n1Ti58QdMFIn0bQ0jTQyk++23TbbInv
7sVOB/b8bBXyPEIX7XWCdCIYK/o8RLIeddsBTNEbTYqRLjCJvUziaDufBPEE6B+r
rHvZtrVdBkdTUfTGaV+ZjifNfkckpg6YQHppMFRq7BNBx6SVJ2w1DH20ukNF89j2
f5dViivwM1QP1p2DRTC6EMAvAK55wMkr3hEK59ywIYRtQ1hkZQP4OLmIKXAusuXs
1FCeEkZ2hP7ciqE22Zq0Tel7BP4i+H0gR1vDXtDUOX7qA56TtuV03gPR1eEdQNpD
5PiSksIW89bFegvfDycwgVJx4fpGanlhT92fn3dP51qOcUYbb+OT0RWKgyD0bkx0
bcBQM2bGkRicywIb0MD8ORj+ZHO9kO/ApyfL5fX1Eb1u2nwI/00mplr65kX8WRv8
kq1L07xKywf9PrG72mW09uKUNs8r+cSN0xiaJRGicGbU8qTMpLiqeWTX1Nqe2aA7
FeVBEV1RksQJ1yinbXj4i7gN5x3zI+aGvLskhwo3CzOZmihSpljHXqh+1hNH0Yp9
kEN5gpsUubDFHWR7ioTlkePDRP0fDvZlaWGlR9GXTQWo5uUmuhuoZboyDOacoEq3
sYDtpVwdvJP+n+7hk7OlVlPW7AuQdKMhNYxKSzvcCGnOhqfLqF0BG9uQUnaHW3/G
PnoyzKqg51GnM1W5GRmy0J4z5XJDV/VblWI1amkZe0suTPfH9IQMkmo5TtR8VAPs
fX3j2vsnPfi1FYW2n0kaM+D0UUB4xISj5ll7fOWU0iUVZOwB8qPQB0ycsvJuwnAn
1m6SkY1FccgRttJcL58eJevsCWpLmsHp1RD3URO7EJUnpAnUOPPh9Z/1q1AEsUlP
tVg+afFdQsXcTfZQ+B7LLdHkdl2e9TJuuXf5pqKennDPnXIFj78IVbV2+ckS4Zli
UnxlYePoEjfmBHq8UtxPVq/x4wYJM4eevfaYYiP32MVpa8QO12alYsbGRRruTau1
iueROetztM4fqJQ4gbT5fyvDDVsuSo18t4PLtgM5nBe2cpMaJUze5p7XVgOpcB/N
tfwNr+5POf6H4g5kSJF5QOxC5leJ3ZIN0sMofl8/IdTlxg2pUE2OO/wVyBM7Pnfs
jS40bKPS29QcTRGKYopw4o41ZI0MwNuGKbRs4bgsbWcFMhN9eGRmrS/xHy/Rw1fc
1LI/bdgsrTQncJN0r4EK8r1kgGv/RAoiGeUBJUM7L7pdSXpml7RU37zcBCUVv1Nx
PYa/te6Z8sgeJMZDguSiIi2Ie9gsiriBqTyeGnMlacGrdifH5nSvuoWQKE1VPkB2
VAIOHQVXHfqynQ+yxgQSoxBoZNm+5icoGNHW1A2/OSYHxwsDeLVFyRZAEJinqjxU
adnT3Qfmrd0NPryTnBL6dOyF5DJUuAWboChAZHcM0OtsZ77nYAXBXgxwWOQMcwSS
I3N8UAewgSM4i2h0g16qbuVuH89ZCu4FaUS2htu4b/qbltrh8yw42TP2H6K7IpvB
aGcBDKVVKoqh8G/9rXehjjyZ/gqU2PSgj2YUzF1iaUMkBdjO0mwrsIC+WMvHdnNe
3EU9cJjedA3JJn1VJlfVA21IZECpHe3gHChYdOb8LcBaFaa8eMF1gbfDEdP+11y6
YCWuDVD8ZYE4yLXyKmr047CxTNa5KckyFzjopxX+vecbi3n23uNT8PEJ4bnSzYU3
SHlezBGpllP88VeJ5A2HJX+MVtNG5QAdDaPOVrKcq6zph/WmyvB0XGqD2TQOgVfv
4NIzmILt0G4uc/rgaSDWK1SPkVdfQkMhNA/nMUddnWukdEVwj5tuSr8d7n5mg1uO
uVsP2IqPRUyGBock4Q8d0U93ApflumBEaEran9aImb+OhcFiaQEyDKx95QWH7U2J
Cxhv6RGoMr9zi9/o/u0w9f0aP6Mq2KkKXCxVfKTLQ+ZJ1e/N2PCe1RxUv+yHd1ZT
IArQ3edgoewbdvnGpPKemQDiazSH/J2HvsZ0I6Cfw8vrMorZ1Al9LxVNHFh+vFOh
RpBz9e3RrUj6cYJGzuJUIalzFZrLpQds3THUwZ5SgVT4b/twzBvH6mwBKfKTW57F
8m9QHeorGRFoWxtAP6SXYbvypQ3FBWH9x3bo9Ho7YPAZKUZnMRxUFQodplex54fx
O0SKRoWj374IXCPbSqcc/HQ8PQLpdUNX0C2pWTMQdyNjQLY8YXf2KMwNNJTrtM/L
nOh+SbSaC0YBLbafdwoJoyIAlG4gFgw232AfqATC9S48PNBN6DnEvyoMa2XApCzX
hUcf1txQXhFOYC/aDrFgsRHmgFyFifsrEi3tlDokIdz0VVrgv3cIG+9RfGKThQ7t
EpEiXYj0sL8rLhQt41ZZpabdV+aB7vkpSQhxaX9bgyiQYXmfeJQKH22ZO5lyu4Fa
z+y//K6Ph6Jo2CcA12wyqbR6Af4AFOpn/da5RtSngmFLAFtUBaaelwc3d7GUAJP+
b0BnL44P+Xn2EBVSPP08FhbSn8hQ6q6fBqyO0jCmyH4AJrn4eN6Mf2REMwgfepi6
KvWSpnR+newVnxeNZNYgk1w7o5UrFb3Wtt5cyELSBc0r1bHCGxPtt0n7EtMkiGRG
E8gO+p8ksAbRIjNC3TmSj2g8FIG+jDsIEnSVH2bQVsxnZZj07XFqgEuIdWYZvanh
+ov9zB9E0jT6qHMOzpEvyfYa6JvDFT8Nz5d+CQW3mLVdc+CxXNNof+Jw4wx1HGpP
gA9UK5XYcGUm37fd6BSGKr0sd5EOJnyGfQeN9ihx4Bs7v8Qj/+9M3RtnhapSnNqn
GVNhMB+P8Pp/i3L9Ywd0tgrKXpgEF7PGW7tfBMjUqPuKVo4Dk+v6rGIPXwqGdgNt
CSpJiwvnpXGKU1JKbOVZdqCJbWHx7L7JW4ACst1kjzbssQQvMJOWgNvn+C87hheC
vzAFt5i012Y0ykfZknV+nxoP1vobC+K6I0pM37fbc1EfzILi9u9zBYwXMXbjpR6h
2/U6A4l9gy6I8GrwaL7tvmb10DZyo2oyrRqwbV7Zob11ncC1Y6ry4bas11+Yys8v
SJEO8gsGxJMSoKTHdH3tFs2dE4jIDEDQzT+0n0kicRSeTsSX6b7jveQLwM5hdB9g
Gvru2NOOalP+UF+OJxk7VJjY8ZRyugGZGusUlQppwzAmzHuKTHPysgQF+ye114SE
sHVhdlsQG0w72hSzruFhzjf2ex1OzvUFsG23zUlS0+57oa6NtO8QKnB0ndcQtFs/
TALyeHZq7EkrcyUEAdM98ANbDU1X1ZELHWX3RlA7TcY5/oqWBnZiwTMIuoQkwA9r
mK0Ylls9oQQV/gAcATrr+agWQLxVEO3BrcgMfIwVNqrZUp8cq/ndACH7e8+RcGtM
qm0VttoOcftB8bEfJX+gfq9hMEyEAJiYEt4+hZ/QTAdfr4Wfq5/2obRS7enIeSAI
54ctCZ6R9dP3NhmVc2EgqzMgqXaopuu4J37QSyn1QIhIPIQiQtGpdobBhObtwrz1
yTdxQlQ0PgyQcOcwW56iZCBJkRDZqqdu+8VuESGCwAdh0ngkYohvBRM3V8HM5YAt
Y2wFeOFo22+AHbhTt2OkZoiGP0QcOBhiaamlQ2CHKSga631+HroMFMZSj84gCPRD
aEG2pgHPgQEfFTy2kUcKkCqvRv7zrICp4VhCJvjGw7SSL/fRFn1fPWv/z1+agoqi
083gMUmmW4P3b34CkAJfdyADyrsUNvhYArR9iwnZ92oirzfJIhv/Cttv7NmqNLG7
sxvmEotc3jDg1dYx5ZAEywkF2Jz4+h2KPEYKDK8DbLCJsY4B2YSvyxpTT9a/tHW8
GTtF2KyD3/a+q6k6wAS25DTtTLzmjuyWuegerPgLJskfxTy6n9+WpO4eU3LPvoOA
JGazeP+VieqiBkHnKiJdoXP0aYDSB6ZpHC15WVJzN0HjR7f01Fc5CEcZYKaUZYZb
Dlw6S/cbafGJ/k+TjxQg7RQzN5jgxTehMjmx/MrI9WLybtK/KqL7eom+B3Y9vYHr
JTlOiECU0pxM1Tid/8//hBtb53esYqvKb8YRUHbWn6VbPmBqh+Ax1z7ZF2JGIWOR
xRWZo/vHiIvY7qdqhHa2tVWh9dxA1D0x6g7oN7xseAm82h/1kQcBPn3d9q2+tr/z
gdL3D5M7lYYeWYLJsL9lKB/VJmtdXAVxbGs4YeKItAURko518j2KsqGgBeBWnkUZ
mSOx1+LtPStZK8KyWG0aPGKayAVwUefSQjdrS3x4x1MWbHSEIqrQQYL/A13VysBA
X6CIOfyG/f4brqYbzv2RxMigHxM+nW76GBiZG0Kd6uUDSSkJF95EOvMhWxDMy2Lt
YtUx6zmpv8dZ39UsySF59TQPzeE6Whj16TlcF1rpCqP5qKuk99XiOChv1Et6hbSM
TrqpRrOpryZZAbJyPnV8msAMHN4O2TDt1ChfksnM7RBh3fo1NrKGnq+efUM33IbV
WBqyTkq7+ALmSD/mTlb8BsJJXWt7+6wymJg8leB4NVpp50LDE5FDGTuXhN7tmDgr
YhHkpN2s5HzB6iU+M7Fjm05HsKEa0e98bkBQXztTLVPobSsisBwuTAtBHVhZgvKW
fymYbbT9rgkfJNsQeHhAh6ToJm59ru4ZEUWCwQue8tIDsA9Ds9V7+D/6s7/8100c
6/8aQ2uagcZz2b7AZqcHpnu2Vwec+Q/g3jAeERaFtnJtS0JeY+/2by9o9nBXAGaP
Rt0ui6jEKfoTCFOjj9hRRpgiNt/fwBtnjNKwgR31Z4PaSAMbkqKZ1U6lA7E1DNay
WSfZtrYognIQ06Ti/IlJgDbDfoyvoR4OVfUokp+Z5e7znCOSyho7QMCf9NDMxD85
8Onw2gb+yHBkLBi48Cz684KtJyeii4MvoWaGWbsQhxN+oD2PokuREONUa1QXiQW5
sz8vuQ5lKxPQVvrEr7RYI/E4vK6Ww+GyB8MaWmIvKiXnYulHZGsH4IbmSA3Ly2g+
r1LP+fttjeCkBUzu5qqPimXteUoboKFGYNxLXISARPEVZuyQxskaks+ed4WJ1a/i
ibTAMLlflCKCXy/qxN+51e6eU2w2e0FfPhspkxxVKHaIV6kfg3kxgrJP4P6XIYLC
z7s2GSJyn6zcQr+bRbZwIYvBzf0oIdMru+9YiXLKVBQNBknOPn6vg3z1LIDA/zmG
0yDCn02VlVOUPTxCtDiSF3JNKXPX5GObovWUfZLr305MshpNzfTi1aBrxyPPuYkv
FybXCvEMJeqo2zCu65qQ8fhVHhtYI7a7bEgWq+vMs+tFmNFwGcZmw7kkUGwjoe/y
GkSfDLC8+0xwewQTujywRixtLWcsjKQq4+LFWlYkz0E1IJ3CzQliD3ygTSahZuDI
`pragma protect end_protected
