// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rVkoYaLaSL/A9rO9sP0m8N7pcOQhrmiEQVbJR7Oy8vs+IacMK37ncMVL/1aqzBI/
AXeHj1oO1rGDsFG1e6gEw1iIgOnuVeBw+Llj2m9E2FdMa1ZpTJX+8njW8wdTE4D/
P6Iie5CSMckei+lCOleOKA2RVl/0eBrERSKksXS1SwI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 123904)
oFAMnz4ycO4kGg0Y+RTjlobJ5Uau0E2ejvV3k32OAJZ2s2A+V1YdAd2/W9l8JBQC
qlpbgZsHXkNqLS5Nl1E6fZOvVysoY1C/gpdL3NDiRUXHe5JZTrYEP3E4e93CrTDr
TpoolIMZI+A6wb2A4NcVhWDKvnST0XdvgF0fCjjCfygQ9CvULCqvdClwZk9wIhGC
4kgDjZuLMd/2iLoyyb6cXb3KB4lRKvX4JtiGtR/uQr3j2htkzyZU0KHnVBX8SAPa
Mps/vqXmKF4MuKfaT0OZtKyHwEUmhTx3tPH6mnNrPnzTDKmsRp1ZX4M5WpYvL19G
oqtwMVEwErflGAkoyk8O0i6gVZaVXVi3GmoK/PzqYeRB9FFhNzRwD9CtEfzKQ+9H
0PnreIoS7FqhXuYmMCntcGIuVNnG/ChhaDYM+PgD08yZJQxF4zktKPEveb2RWIBh
1luOAxLkN3GwGdybUD3AN0dOFKLJDrnmBEmn56kkhRoMM44PLIMxS7CB0Zgr6WWw
dkELeqHcSUSkNyBbgTwd7RxMmWatwOvNkXTMpBvgnXK7JF1nU+2akMS1w+RAYj66
EhYHB9l6XV/PkD3+udtazBTTYZyHDh2GUQIqzs3rcQRKltrkIbsW/ld5sMJNc7zS
mM4rl+EtiFeJulMJDkpVM+E5glASNe/dAb5lTqwvLhXTnXqNuPc13Fn2gx/xZ2SB
CNXlZMbC/Xw5Z5DxvP2npuYmEJIaoC1kN1LdzACUGac+VnROrHdDl6V4iJJWIr50
AKURDE6U6iEIoUR/ZGBz+wi3kapXY7IBBYPyhbiL1DMX+w0FYQkyOuDgpkslAy2c
SGKdvZ2ca7kzOB6g7u9MLDMebE7GIUjUpnSpTp3Yuar8DnYpwMP3ZkLDdhJ8rDUm
xJkHVq8bf+/bl9kU4MHXUoXTeNeLs+6p16z/EIke0OpactFQ68WmrvbgClyfjRLC
MHLWl4mp7DKSusTiNU75CCeYe24nwrVWF0DC4Ccj7iiBsPf4/pW9CQTOqX4xVBT3
JXFhHeA9ck7hfDjO2SlKKqYPW6Rs4fBWltF5fSaugMtf4JLkDLKJU3gTRffIg1sJ
eNLY8ajyZkeHSGmhL06HjuDAX3ObamJwpznwnjYcwww9R1tKWJNXC8TOzO9X+5Tv
v50MKhzCWaGp0C772cTEo4GwMRdT4E3LDfAfvVOujJzrXqghRksV5dqNQkStP6UM
3uSHZqEkWhVDCXsZ2GK+wwP8YkDmgPtgbZM5dsxbwJ0LSa1a1qi5vXfxtg/WFMND
aoNCSLGOijUTHTnQ45kY5qX+jcPN+SRXjAUjaaPtj00V9+vSgvenEQQQcqx+VRnl
BK3CAmSIV2/6o4KllZvW9QRLj8XpigcWw+Ol9yJkDOQb2ysX4/li+jjICgAbggJb
+V+nAd9di1lPCnIElKCvceIKvnDVcgZ/ZUWWBLFfWRzUwfHlPK80hIE/+eWE9NN1
28VrUQG2n3+97x//cth9oK3MKlJOOwfe88cmdnuAuCmIX+hgbYzpZi2AWRb7jfNI
SOpC61fW0jotX6Is4zx+bk+ez6wvq0ObYB7XY4AT1+S41pXg0PGeQFZyIjFzINz8
oD2oSm7UPoyxrbgedD4dFeHMpwF8BW7K+ycWFgFC130x7PfB97ScfNCJ/I19abYK
o4xvU9mVtxfykxCeKP0+cwx1y+l+tWBa9/avncjB+7HSKKtiuaKypGiG9RMoONF1
3I79nlTjUqxBBmhAoboPgbeL6cmgtil+zg3x24nL4UjC7mtZaBeXP0ENerV92+I+
Smk5lMFi1A9/+EoCXi9HtPo31mAAxfW0djLkVLK8/me4sHAjRtqB4lli/h04kE32
sc5JZS5O1X71O++iNQk6N4dQcUGm8aIft4R1Jqu99iPptai7wDq5epd8oSJhTqmM
UWPXHXhtOxpTndfeFVivEc0krYFLncHFQbO7GmILVN0I7hvd4m2tdQYpeTHWWV6x
ePiq6pdoEAvXEawDsXwxkb5j1dwAZkI1JoVBEAWUouKOtttdvQ3X/p6LJVV9fus9
wApx8jQsRe1otY5vmEqfLPYH0JZz4lSZwtPVblQy7otQBbFLfIeZZwdnJBktjrls
9UN9SUzvlNY2Cp1kdkim3aNfhFzdniW895jnQZO3NheV1ANPZN72lVEKEYDJTOZn
LOpEVrkSSzaBnvO4Ob/8frAI5rDgkCWkp2sw9um6EfN/HWgFHTg2gBQQJmp5HFgP
xNxqh/ABDonh/Isfah4Sqt0lE6WPZKetbko4ZodOqLJkvhg/3u3rcdr2oKnjMj56
Dk+Z/+vEInFGuiTBH7pCH65FxFVKfGZC6qBfqp9B1OEEwtX6HFrfAlMiKK07idxX
bd0k+mCsXK0/YZxtrNrXOKbyrScT+n+qFOE0ol+Pgn/AtCAwB9VBR+8qHCtJLQ34
8DhrZ4zooD/kOb6IAA2NtXWMIO0OcqJr+c1FhoMspLfGIkrwI9mRyWcltuci84sj
3P2o+gHh653G5CDReGJ/wsWCkyi0LZg7NUHCMZ1otgaXMSD59GBOW4UCRtYlu/Qm
VzjJNE7y79GGyTGXlZsbq5+K2VX0294Ei3DmEl+quxcIO0fPDOAO6lcuMLesltFH
qAFxafvqffog5tStc5zZTHVrlDp+91xuUmShT0TKBPwUsRQ6mhgWi4i377huQv2w
ytFghAjyGx+tcubq1vFVNQNlDujATvrv40N6K/m16uPPpWriBEViKcJJvrLg8caY
JGaI/tvqD9FprQAwXWkMxQbP5JDcqqwl7M8yYWnQaNCrAD5FBQM0//eHIzkqQChC
4VA6D9Qf4nEJBRfGgnIDbWuBzXSGy7AoKIGJGee5kj3BFUcox1LWMuK/YrkLQH1g
f52PoPe7Ug/PloAwvOAs0uAC/ju6VGHzq+tpH1tD8V2X6TLZ0q2vBO8Da1Na1fLV
lOe2kZafQ39N03Ui9C7R4mIaZKQcQt3xBdjm/3pQgCje6zWXAZvbZe4ICKwgF2uO
uswGl9CioIdwynyk6tZrbjdL/llJXkxc9Y3mWcCQHqG3cALdVixVRTpVBONR8IJy
lt2+t7kJKJH1g/vbzIkRygsa7B0KXolKBN5ICpR1WHXODQ+arsyEqcRAZf93EzbW
bGKTR7/fBJPd/hgZ3pwa48Ql9SGctix/JjusDY0LLELk+iv9NXsHhGul1hrHfuwn
qxnvD45IvgN+vfPSAA+WBFEJaXi5GjGZEKsTNYpqO57O6sVAURSy/cOe2q5NlDJL
fzJn6AKRtOzB2AUd8KAnt66BSoIfjLdOZniNmgsYXYud2z14htPJj5vbi3vmm68/
Rc9ODKJEga8bdNicD85dU5pPEGoBRe7MFJe0fGtD2i9vLrpFbQ+R5EGoKUw6tT1I
D9QL7BM1iqw5UHPoHe0ag0QYR4ASnj+qXib5ZQ51rd8OhMBlPa+HnmLNigKPkb16
w7pW+coKXMqf76JHsjB91tO36HS/Tn+oOSk64ng4nDI1ILqRla61wJclM1urwypX
QufXM6hmqUdGy0HE5gIlB2IqOoDjH/L/LXo9Ea7jD2Znjh+Xwas/OKmskH1sCCNj
OdyCZ1R4NAOUaArCG7KULsaS8R0eH/pAF1D3clma6p7i3r5fy6jYY/r7yK7idKhq
ArueUTwqvY2pODKIZMryOviqdzSrhMcVzczochIFR1EDF1Lahf04fLlMwKiXnUsf
7NIAla7cO+04UBdco2ihXOmw2sPvUJI+r0jWKa0l+Cfrq/Xf33w8GFfhsD7T6mOW
YxgKD0fUuOEBpVQeWWTTiwRJ9U9bgAtTztZtXWbDZa38w1Wp7UZkXjLCZWJiALUR
Xbt8J8qIjtlWy+RIEtXbfQ9ZEhxGoMP+I/4g0Nr1BybQCUDCB7jpgU3QMHI7Ybz+
pw5X+TjC2JTExnVrxEJgerw0UCNC/qlxgy4C/NHYJSzZ0IRkMyaT/ZlJxVjGt0hG
PJ1PR9C8CbYLOUw5K81uB/NcawRiStJZXgBLbmcSywMNWmdulJx+k3ElmYsMUGhE
CVF4NHyi1OKZo1JQSLXOyomZEPpKieCVHrvEOlqyRFWuJratKY5xsuhldCD+wHbg
/HtVxqEMEMQ4xHvtAtTbqhEDjOtVsLXmjd2nHHpLd3sro7epF1SbKcfCUp/UL8Fm
gYrK7UVIsHh2nEyBoexnLNblPL8kGqHVint4JhYm8T+ej+3aozKs6t17AAwsarSk
srmhTgauNgucq1ycitsoKBDtMGuKO1I9DXO0KZau3//tvksBj2fGC4z5CBDIOhbz
RTSEYmF70YYHZuRen0hIiWI9a0REfar1jG1gj9jJntp64ZU35U9MkNKgTGVufrj/
TtvOC0V3/8075JRI5l2rvPL4e+NuanqNpLkbU9qXFKyIMTBU3aqLJcAdHaMNkL8T
y1i2WOw1R9/MTtQESqNnVy4rWmq390dfY2oJQ648x3FInS8fkR881St01MKPvdbc
5VV7NdFVWEo/lw9/b51zm+S9ThFep3rO5wf11CRsqehoPRndYPu+apaf0G+dVlCK
n2+Vg4TW+ZPtCDHw7G/A89SyhoYfP9fVPKScV+TbOUj5zGLdB5W/HoH8HPeHFPYC
6moXZnCQ0+ZSsbGzM0gG2d4oRX3oAmStIS1W1UD6Kyc6PzcPTUfVpmLFUMlVP5Kd
hix+oxCmFJ1SFGkLP5kx6lgpDV1eS+iC4gCSJN9pbDJx3e5YMz2/HFxEx+RtawCZ
BREmydPkcwBKKwzJtkBQW99ohninEUn9jWMv1FbXhbMtV2D/ggexNQuBMG+iqsok
DjlIUoP8PtJf1uSObi4X5p8CBdG/M1RaLZjc86iMp8zyVMSlbgUdUlFNz7ur4kK2
MLVx29gkif/BZGPZZrxrerERsiyNlX2fZmiLefWrYT4uZtp84PakuANkHc6Yh3XG
hykN0eqrb8lLUdsjt1RCco2as1F8BlwwRvVJF4RO+QbMJjfpKULgs1ZKtB901ozD
NUSLOpzx1WaXlmBZOLdqzfsqXPpqeLxkM90gPvszvxxag7nC6MORoMeGucOcoXk+
f/3cwFraodFDr4GB2O77R2DzERcRsPN3DQBuQHVuzsjg3dQ2MBI2pbc8K0jRRMg2
K1ZB2X7K4/dvlGqF7iEAqkoBiROOGxt/KiRNqXQJDsbolj9lgbQ1vc908P/TuHAb
42fpET5H/U52FFXTTho1UG0OHyI17n/3+Y4lkQEA05SqD50ie6Jb0FbncGYOxUK2
zrvSdQHUq/rljQQZlmiQtCqGFEHUk+VZqWYPMOvCR58HW8cKG2qI3qXN6GALbw2F
qGGZbW8/057P64Vz1UuCKlkRRJzzM5i+MuckHMccFMexn7Zujis2WVPOp9Ft3S65
SJgLMDj5NvgkJ+Vel9cf2+1IFIbf/yVBBkzZDzi4d485s7OsnnZrKR95aufktOiG
vf69XdDWpGZJe8lxHMP8hhfsatJMcsf1H4IaMrXJu80HFodnKoaQSd1eHfP9+vWg
0rreu5BqWE8/M/eAL5Cuwn0KvRigRVcqOSud+GFZK4A9z1wcOLsQ7qGU4SxGx3on
xDsBswWGqbxOMAuW8l97dq83UQIA8rmxxn8AN359axob/6DMDcl5GSP9b3u6wzlb
bHRTf6k9ohaCHqMYFoGeynABAGhSu/LZSD5/LqtYx2aCY/gvygAjtAdTLUk1aJQs
DHtmXp+FZM4zmN+KNdV8A4TLt+nHiirEbbYhsHE0KzlugjW3I+zvBXbgghlA37MR
6ygVmB8YfJrerIk09zQ8qZQwSZRVdevWaI/TXcf7/R8DhOy433PEjiAcZAEr3S5j
T9o4lrkUxjs9O0VlsqAo43cMl8nR9SuWmLZJJ52dSTolqL8Nud91b50KWxhW29Ue
GliPQuyX9VuOSm4Xc77Omdm73claflMMyTn1Aqkt+vq17R0eK+aKVF/Agz54tDWD
/GGr5sk5a7sIPUU0SkPZFA3XgV+c0WNOudXGeJOJ4rFU2g77Nv3ftR0Gtlywxzzl
K0p+scSLSbC8RO7HFcL37+pTlXnLs44uOslFnFzdvN5IztjnH3z2v75WNuSFOY5f
URaAoZIJ5bKttNHMF/EkGD3btz43GMWtRawSvPZTf6VhI12dFxB4MNMRHRq/wLKO
I8haTXTziCcoe09bvD8sNAJnJGdhuxG6fDw/GDxq9Xz4vYCxQk9Zhonl2trmSPTc
7rBXxfeAjUKQQFiOhIlupDI5XFaaFw0vfkLIG1U8xq83UYAty2Oom57gJDGXXW/0
EHnFW1riiNYuDdI/YxrZRGUWjdRfEg73fHcEzezMA5HxxohXo7E/PEVv9mW7E++W
VMrPYsn11GM2onn3o+GI6f8vOVruEKNm9rZPQugFVO5eAROrEzNwyYkZKG24Fhdr
AWo+VA6Ps1/ra5EGEZi9nkNpQCtg7jQdVPndhTy2P63bV6SszGToH8BvVJyyn9RF
POncdhdzQuUnuqpB5g8h97sWvhJkTAsTUoPWnxfMm02hCVzurR+FJAt8ovJTzbC2
3WQjl+0DTVeNtJf39tUpDqpeQIplR9fdQalX5yFJt1tgAqzKZ8viexF6iwdOCI84
/FXGRF044w39bbfSR8KGem3gFvikXvDmDbNenfFTw4dDWrJd9VxUPRoZmRHcKviK
88JwoKX8o3SOpfNhM/ENTSZFRRFblpLZja4yxkS5pXGF1BkrpAxfDnbaVkW3+csB
vk1m0doh0jSBir2WKnLsNtlUwvacQ7ulU6QWsoK5QuOu3zzskBebGl94+7bRgYUF
zIJe+WpHT9BwiARO9g3afKxaXT40Wc0ujtOX5fhkfh7F9sSXYkxo0Jo+I8X1Y5qo
nE+oZLZ/OL3T261VF7Pg9vlKoi/N4OOqtP+wa2tXemeQva0IZTBbkYJ0soNUI/74
XDIEGP8MGeOBpIIRXLKWIg6ZAUvS76cBbjnin/hRCrJVqRnjppEjNeN4xB9pIibE
JYsCNXqSk9P5E/h9OVBKRDfRYxJ523HcEO22UYnWoubcQIxtQCQ+S0P8H5aajCkH
G+w/ViprtFX0wQipYMFYBG/s3xJRrPV35vmPLo+dIZvhkm5/Or/cPkX/YiFoIdPi
JRzjWRnj7DE1G4zh6A2vQmzcGYtJT4liOSoPUUhgmE+O1GfWjMLjuNIpt3lpG60m
qRYFLQBHAInMoi/M0rSMDLRzv40xbOMwqHfY5tvEtsjYuO1QRi2jDKgnUzMmr5gz
/scCIZLsEvFQ+JPnleKMpn3l249eY9A3IJkSAZ5XYjdYV1/FURk0pKnG/5ZMMMgj
kCJhYNaEZvEepL/UWXhK4udLWxFeaPurwpYZKMxoyPJ4mX7RIXbxV8Xbemmdyern
KG7uAO9AGrP78gEGyzruxx93MADOi72N6JANyPSUrzGtPjltFse7qlrXBGhERXM+
RHqvtHo0jk9oDXa/lFgUmzxbUw+s+JF2vyTGcZpfLd+In9io3OrWzfAoO0weXdjH
vW4xruhmXcNjd+ta9MknBtCxs7dbM4YLIL99SxB2ggM5w7vlEYouAiDyifwYxJVv
1Hl8XJ81FSr97wM7RutETSqKEtTuvXGFabJk0GVbXvMfbjtYWQ6KiG6fAEXgho5I
HVDYbYViE26xc2o2zp+2y4Eu5ky009TvH1gPeSurHfBtKQViRUI5sSMjY3ZpiJxl
H2DZm7Leoe+3jtnkjFhiUt3u5sK+cHkaC9PdbNkp4YWKM/P6bUiH/5IPE8IdOTqS
ntYliYSreDSg+BsytSsVjGurELTPJBcBpnb5IUHVzuFWgT7b/fAbuO0all2uvxWe
6wIPRu94MBynWNyLWccItB9V5omKPUN9ZpWKtKsKjsIMMJljgYt/OF2NK2yE52Ae
J4oXjYZ+RW+V3R+k7S5CdCb5b0GbVtHuJHmvqmh3sBPINDL8BHRMzBXkdE/bjsu9
BUT7CyNLJ78+Yt9URM1Fz471PNnrxGH8tEfbMF+aVWwPD5BS7UFu7y6LuCa1dvMl
LOgG1rOqjPEXsUxfHl5ewzORjPzPPtF2FoKGUNx4lqnvE79s8vlrg9D1mOzrDLpY
lCsgPV4MNsRSJisjxUA6xb4hXOrxwtDkRdE8aI9HK+NdoI47CNIXqN7CQuiHfX9M
Zjv0oS/6M0d+K2IKBdVpAZHQDvMy07AfPPzIOvHmmR5DVUk1ec+cxPwsq9XJO6gF
nG29I3cV0wkd4iCeNaer+Rq7eJ9zIQDMSyyLiVCMC4UhnOaN9ZxAa7/aLd3pVHn/
GEAe6X0tlf8R+f6NF3DqKiBxDAJJkceIyyR3qyzD890XIjAT0MC+JfYNihz817cR
TCygFpG4NsGK0dhNzfmbGW2YjG66TMYLlEWHUVlTaWDtQ4gu4FsRVRSWtkQIXY+b
dy5bhvfNlbJM0G4ph1NxrKCoryzpQQmvd/GjWa2QZmhWi16b1E+uxVtDu7ijLEKU
IP2gd16aOvdls1h7p9xNh1TQqGt8qsh1xNS+T1K8/kCPAmPSn4MhMcFzEmZWmN+z
SgXHJP0vjCzs2hNV6sWb0SyFVKxXPQhfKDgBVoGJhM4Tjo+5AG0XQbaxSUmweu61
Pl6A6Fiv1dUuap7xg26CX97HxMBiOENDFMRiIZx1b9axnQmgW6TcySLoUs4giVgC
mJhO67LwTGpKjHRTMRSYXKCLLZuMZ0xHG7z4eMtc1MiUoGL3oM4JaKIdjG10qCQ7
wUlvLpoWzu10Q/yw3LV7/zNO7JjKcbqZSBaP8snUmx4iJ9BQR91UuW4mVHmqzmke
a9JpDWtzffOfdWZcmiXszTNIVMA7PU6fQIxh/HaYOwaiFjBMDAe1UKNN/jHgVOR5
VJhuUv2kwVEpP1jLj1mr+JX5sSI4r+KICJ/rmgz2XoGQgyEEAYTQl3L7dqzRjug9
rO9Cf7yJzPWp4tzdDbB10HbpWJNj54eUGzzmWGjapSeKrTnICi/xPWkc4m1GpExw
awVZc6CQAxZo1lYTC3ByNO4q7x6i6NFNlUpkXndDRYPwjnCB5vGjM+y4uHeROoMt
NVP0PJhKtAcgRFef7o0T7kOELdnqEem9M78on2jz1HT+ntMNoUONpawOGnkW/pu3
hzS4fXkZSSUXaPUPylLZWJvHGB+S8/o+I4c81Yn0Pouk1S56lRSVVHR4EUD3I4Xk
KZaewDqEoThh5slM1K2KP2Fkrpirv20j7VLtW7CTtW43mTNheYwNkolie+Iuu90Z
j1eOJyqU0k4MyhisaYDyAXrinvLQB3FOjCf2fzbSyaEBzgMgqDci8/4x4B6Nn4iK
N8tTbQkIEvbPOovzXe9BinoFw5xEM74BYTFxER96YWVB30vS00LXKgg2ARJ3G4+w
HbNRNHHughleK1ZNUoYAyrF8XVS/XrMA295saIbjjgfmLiVFpWnPAeWrhoZW/gx+
nWrI4hKiDnjpby+5r677a37TIKoAWAIrmm6l5Gxnak1ihn/zem2LYgeR4Tp7yPgA
l9pkfeP3VhuRWQ595f2/UTa1eP+QQbHsK4HgtWgZOdgCf3ObXuAPQhn1SFNfYw6N
uFaXr0PVAGzpsqySjCXqvZln6gyj/Vt6x/8pGA3D+nMeG5VkqeiNfICSJOOl/aIq
pL4TD9EIvDozWS6wRdt74xpSi5CcsNtD18sUqjIvuSG8jHAlwX/as6LlRO6sjZRO
R9YTm/IHimzGMGY0YKAGTu5shP++2uibujp6W4WXSUhLIGZK+sTmzPJmzNLE1F0d
1KeF9lJylEbOLXq32qzD6SRhjs6Ng6uXRJ4qjuQHO2atrnMZnNDaCSfmmeueeS8e
HSoRMGBuJ3/UHEHpZ+311LdmHFmpZzTdlFv/a4xjxBGYIaxuR+Hx30rwXY94wx/W
q2NYFNyrGLwfP6bDWvBw0RF9LQQRSg5wGaOR8wSARzQN7RwXfziEO8on8xj9JTkd
WkK85JdPCEAKEgyL+/cKKBvX75ju3dZJyUgOMZNT3a+MQQjQpFtbJcCLHVtKSgm/
YLwdi8fZVaRWps3KHdZ8/z7BcL0W5SyUiCa+PmoWRs2ufdWbUBbf5FW/hAVCABdJ
ip+BcvTmKA/w6mD11rOpeerPNNSsibzMzPxbFAu37/AC8E9TxzWo9wsEAZQy/JX4
LwrqxkIh/W/mxOVMx3lfH51P0FOw2rBOOACNuJ696WzQ+cK9nyth0cx5q5ss4QIN
ag8D1tivnhttYbh2nnCTE3jhl/ozjyvDpNctxiii3ATUsBp191jVuZs4fTEdJ0kU
iK0mDLmVFu90MbircTUDiBh79daFTvjipilukaxPaeHxgybW2Zv/znPvPZicxYF3
7jXl6odLhU04607XvJ/6pnRzbqZPpWtT3HaZWPCtGow0qKS1eM7vRLNiOfHm3igp
O1Jpe/uGktBhmgGPn+v8PYLkCQj0gRx146kLFNAj3+olJgjFEFHkxAllfbGuR1l1
lrwYG+cX5nnty9RfRZuVAhY8hSSl4V+E2j70h7l+2fzgfmI5K+TF3XiadHK9GgTI
l3p8sjnDFEeUFdwaNhyb5bXL5D61cB8b+UHSbcS9cP4mT2qP51pFVFom5IjyQ9G/
qZMgJq44aA4u+kEy3E+QST0m24zSkeElYntU/1x+v5MyFKUZs8ebmgMmYtMTV6QC
ZoNx7wmMJMLBIQJhliM9poEhDJLyuYO08+EvaLoEIr3ytG8lS8KslIDVWY3jlxVf
3eWxul8opZsciLdHVjqctdAaU2RgxsHLwnfb4G2NPQ/bnwU4d8mAIaKcPMQFnyE4
ldGOcDH5ZQKxuAbMCpsbOaP/44hCaClmXbAomOH1f+Ub0WGiSfLxG1ljr1AHv0OY
V0fiO+1m5nccJ4i2ZNMVSCpvRL6XFnlULfYVNuueo84KimtnOTTKMQyU8xjwIP/D
vGjNHEwO4hGvqba1GAmEEWIeZoKq6qhdT5JU6d2PhJiZIiMiuoqxqIRlvGglsPqr
bS1eIhXff5QfF+BxCPM7PVwpKFVyETSOuEDXImEucRT9IQTcqJnkjSSPt7/lth/l
oJQRUUQhHyGrRRjLAHPFm9YpfWM+iv6DEN8xyf/W7uR13/wdKIT6fAMU4qonbfLD
HtdbAY+/KJxacdckvW2nFCpZFSiMzyxM7QSW9DVlrZhflfZU7OcbVlCW28EypSrf
A8IS/6d0h5f5owgwgiZcf7da1LbkTjF2x8dZjByK1I2A3UPx0PH03kwz/DOEkQtI
UJaY9bp+lp8AU7tvtCvT9WYTyp1sfzZEF4DZPeP5g/gavrJDNuU4cG2k0t+MEyi0
daX+Ms5qRiacwYpsrjss+XXMzHaPYAubP/bAHZULAXBFyy3wNDuJrpHGOd8c1Vr7
9KRREHtl4RvZzT1XnD2XCpUjx+SEE9Afhe4J8Qrk4WMAVbqieFKqpVE9P0czck6D
iZG8HMLjTZS0QBPRojh8LpfczslaOLcJEA6YPVTDQBcKafScTaVt/gvWdpbvuIaa
/ODgpFFwNWyvAh1ryIo5UxUITIUGIUXBtUgzPC/TUgsjueKRTz/9HtqF4ErDADPh
6wYJk5eOZXFf7NGi7oOS/HBEeDxb9pKCKmUrULcpvylfch5NoxbKCX9v/UR/geMw
WlDiWjZBQ2u2JLWq8GMDPoH0tbKuvQ7hoTPhbpOeqeNivWzoBqpUUEWwuBHees2f
zSUJqCIzXn3U/JrHsmIfLH7m8HoGtLZgNvEhOOSLnG7mabe5kJfwn5ISRhOS8llT
DxpWfkgQhCp25xVgq89ycQOAf58GlYQedK6/ue+ggtBFRpf/QD/YveA9uVhWNJlo
2haKc6lAYRONP77nnfzcJTbSvz7pQRt7MKoMNCFYJhOGvYLIkImJ1gpiYlnRL1sy
FZuREEKeocqZvy+tVArNlJ5dwvK39nzRml5rctVcouD/H2zFJKodyg1VKw9u3Yx8
yzYYH8no3o1lahGUD/vHO4ZTV7Qp190H8aFsSa4g7ZLoOlSMrLDJBd5JZRLff4Ou
ZYvut0j14XqGOHyqki30HFnO/oEyQAM+qiMIO/ydbV24syMhkvRuWoT4dgfcfvaP
IoMeiTcMHYUoJ8wNC6kYzPucOKuWT5iRh0O1ZPtwTAQ4an+rccgWCKhL3YdMEUBM
RtrrGNrv9mBxaWrQRJoQlDmPSCg3eCzLAgGKKyMCFEfGyTdCti2apRI/lM3jNkcn
KY66wz8uEQE7WUuWfjq1WXg3WFsJUS4gN1WdlGiImW5sByVg6W463f6G4U2696mN
wDQu9fXRYoj3pSarTwqx0SzMkS7ZercLFQE7h+KSLdKqgtf3AUAlcr44OOueptz/
KUjMQLc0m03Jt05NRShqgiVUVNEERsSu06jx9/0YPg6bk1s2iNW+18IgveDqs00D
1VSVh1KF+sYn5aaC4E1LZmiori7xwJAC2RZeIPwdboVFlqsdCyYZx/Xf5zcM1gcp
2WNJAbfjTo03eZPnsJwE5BsiCcinC/hIhdvk5JjKj5LYJYkLOA5uGzRzTMXn94g9
E6KeDy8tPhpNWa8k3VlonBtFCY3f1XwfM6r935UbZldtmJcczyLYFPPi64se38J3
Sd+u7sEOa85G3aZJUDAFrl/l+OpzAWI0WWBpPxLOFZTTE7Y0tmfxmOYHMRMAra3N
KSffcs6y/T3N7xG4x5wArqmoXJfpVJ8fPGdJbc/Y8J4FE4cTiYMVdAE7Ce7hfbEW
i4kASKbjD3XO6dhrcQrvLE2Lr/fMqqNk8cmCspvBBV5UYImmmG0KJyPUz/7Tw2V8
TR/8rXc+A2VYptpJx3hG+ECAtE791Zxhwzpucd30kTNfmIS4p+L+NOqm5JgjNNwq
7LVi6NnErYloye5IXg/TA6MK1ftcY0bVtxYh5viAKjUqu/4Gkwz8W3ipeCUNFdz8
cmGHT/+Y3/0g6Q10rZNf3ru5nuITAknx+Fm/zSB5sDiJnbcnxg6s6EvSj0HMLQSx
Gz61nzl7Ya/dVQv8hhr8i28FgVFM022J/zXoRovlYQLEBnkIgAztS6kD1+bxLmza
lTU3m2yYEqiHT/3aT9Nsn9/aNBWyEM3OG3vLs63QOvwKMeKvHSPJeO4ex7t1XA+W
FdRp4M+BDktHGZ82NjTSFzzVa11fwlDilsUm1cur6h9db1FXxvp9s4VC28MHn/5K
WwzLgUfOez8buYFIZT3/kQi23eaoDYRc4netZfnfn+BbW37zCbF6URvpkfWF6Rj0
NI3LVkbVLJ5ooOIWmva841BKi+9R5+pRVCz9pIxU9Sw/53xm/FpU5vse8lT367D2
7RjHnVFDI+aVEamxYJ3w1au0n9ZvTn83TNiUskpjaP193CnGNvKV0o2SkxQyf5VO
T0OBoxKHcvkpfvX8tiMfF/FUAqXmIRFiTz46pjDNO0fh3ETYVEv0fJXRWutNzCw7
EnlH3S2KB1HeJ/TeuOhS0sB4dVOqnaHUnoDf/2MRQAlbZvcASPpDqPBjj/i+M7Z1
pNByrWiXnADaDsDI9AysBem/oXK1O4ojFwSfOGZR1ZelhPzN3c/9x4tCcgu/VlOD
+oEFG7q1jMgwwyx/iZh+dpgda3FMAdcz62K2Qf36mE0bKSwW8tTTdGJ3Fynndhhf
uxi82teir+Q9Jz13JSK9Tdh6mihQ/mt9sU29NimNWmgQ2fHowXG/lVQnjs6Dqi0A
zJ2VMZiASOIbUExk9BHAnp0zarPmt05hTvak4coL9O3NwE0KyOuGRbmTRk2aRFdH
dXohR+b6NYySFb01xmtKSl3NJ8wvQo4Vfoj96h59REilHYfq5ax1y0LkbIYx4IgJ
0BEmhYtChEn6tSVn7OUaQLc0g2Fj31wSntmaQmVtXEH4nu4HCR5WHS4I8hHoENzs
tiIGdW0F//ipBJ/ECix8sZRn/RbloATm7rVoSr5WErSBkaNS+Tq/UIkDhXJQk4X/
qD8rSkodACU9zHsyti2nhjAmMF+L1ouY3aKL8ACs/huR9RISyAND+uspO2TG09JV
UHHgFSZXoidS+BHlKugMtqoowlzwqGR9y5Sk4VpISai1Q6+tMo2QwfciJBiqYT3n
jpxKYtLqbJ0DJvSyCl5nLhg1Izf/lM9WtT9Rff2vZggw3jPaMgfnPYrFtWie/hVP
2QL59yzv6Igwn5HMk5h1NFdfV648tMLeR7NZixFfnnGcKZdeV5KZHraOA2a1IVoD
g9D1HP6S/K+699PpHy/5a2nrpZPOyMJKwe8Rbrrp/KqeWGu/6R57jxli74MCTEtd
l2LVVINqZls8MekFJjYrpejOZm7EAT0uTcFihqk4uLeLMsqq/ZxUGn4UDewxnqhS
+lV1YUhkGfmMb40wRQZn0pB/RqhDt/rXtZSt+eAqUhhYArQdsJwIj9X+m/lELGJA
f+XQGN00xMpqJrv4d4tLse7eRbY/hK8ghflXr50xexVaVErvcSHur7fhClegytV1
IwFwu1rVr1Gs3xD90t9tr81qNCtqcX3INE49xLhfGs8X2MG/6JkuWVP7IFWfPTF2
lkWnZXFUpqWaChPKhtQkd9yoOcLbblUIDHh8MXMpcZ5FMKiYxhSIa1YE0SmJjjRH
ZBpqSDtzJp4SN+A/Tp7GwxXAqesdH9IVfNGoPKBOtGGc/0Co4E6TOCnQnpJAdBuk
hsjCNFoeFA3Q6BAkTyp7RsUoABJjUCaL4ZNLFlu4z3FdxjMctRGYIWwxESvtE1h8
DJXSu5fuMkLhtL5r+/7wK5ym3V76TvD4JfouhEeb1EcHb5z9GRkaS15uKenv9Nwd
DdCWu+nzishlNIwZhT21u/424VVI9JT6WtpMNFoYakSXdn68Xj/ctrt5Eh/+Lf08
rKdLS9SNenCZWThe2NVPB4ex59SMcu17ihmUxeDNgGbFBNtD7zop7LZVrmHz1b00
Z0KqvzuEyklGg83UWfMOwY74Ychb/JLTby7hXbGQL3lj1qozGJRRgdlkTJgD11hZ
2erLmuhlcWNgLDaNNm5r/tUvSokC2bMLo7KRSASCXUjtpH3fgvwvgNTUKdUTNpVM
QTWhw+ZHaXtMOmxNwJfaJC7ApUfet9TmRZpHJ+mRDywt2vLK99/voD7bt39M0YMq
EHNk8TI9ph6lQR1Rg/D7WtJMtl+pegLxA5kCVNtjFJffP5OXr/pSalGqKhocsUAd
eogcO/hykc5DFrqdZujoYURC58n/QOZv+zzDZ4MCE3Yav1+Uzu4i8tnL+hKLfi01
qJF28xQZ4uLCdke9mu7QECmjQl1LBni4m0hijN3HeCjAvUlhIDr7UNuBkY+grZCO
c/IyC09h6Xx6f7lnATir6ej+bfZ5Dx+FIjSvtSnImMGTgNVtmL6AiQ2VjrBMlCTE
HXt/1Hi+psk5TJ5Hgz68okZXFhEN0b3w/S/WmQVTQ4/NNvjRYQ6VqrA8/tF74Ms5
cRDVwFsVkUUPDdjqQBkRCLSgPmXMGFfc6Aryc1r5xvh5kGGaTQafgorPyxo/+Tp0
2QCTAATv+HbK2lNpsRnMjirHH/ERKfEI7MLuXk30ALV6tOBUBgAhiG7TzsPCDeZ1
3zlCvNTlAam6rmIwqM5wyReiMyWqyvcp11r2QuIZdqI2tI8wiWoiF/+zEknhgZMf
q0eCHt9GMbqZGkgbNlu3iaJghqo8m54AgfGq5/oNd9GsQcxsR2PWjHIqyXjXirLN
HQNrbKA7kiQ3/0RYcjVzMKRqkJ6rLLsBPzSI2WMKXZ/dc34J8CfOn5aDrPH/LG/n
y3P4GAhwtwKq2PookIYSkkkRskwgQi+9sLl3zVBj/aeaeI57w8/f2VA1gXjGHuzK
o8A8QfsKrDuDYihK5fpiwQAII5XC6CFGxgMSRe+Qd0v3XYo/L7zXemKCr+F7D9lj
i7D3zBIFoh9J7IQ2pxc9PvdXnpeofjOw9iWoHnN1wUpE+GetFPUhNOmPekMCEj9g
OU9QfgJnZoAeT5s+10askS9aKymEOY8bT8f14aOFil2KDA7V2O9WEaFPH5Cvrd11
cTN2RWGICt7Z3KLI4f0H7WqQR+0YX6Ym05InWI859ZTEQB80RTSWahWEXDQaPoBW
k38pFmp3AOK8tiEzLPoqMmED49rcOsj3H3q18VmZXLoVCt3xZBxZZ7WdbNkm3Uq9
M9I9dpV5wn/jt2OZ5OVKH140fZndaQStNvCG3bf2KQ/kAclRHYzkhHq8tfVQYs6+
zdbrKycDNGlmDfH5EBGRDu9Xdm36jJEyeDLt1oaP5MMQ6yVt4MfmYx7BODclxLQz
86+SIgadFAcVFHJefWg+gNQEgEvPKeJI701obsvs78FlDJ6bHR2ThLOvRllgibg7
JMBrB+LAyLIh8169+O5obnAupBnzRES/95zYYrhGy7HtZhs/AJ3A1Zy1lR018LZ6
d3VjdFLiUGrbaygD/z7VveMp/jhTI5YRYmasqdM/x0X1IqPYhdgFCpuX4A5kLrxW
mSXVUwlDDKbL70jeqz7R8X1Sv3N4HOGh+iuAn25y+ir1m8TGiK3dwZgTyCiH1Tl+
19VrnOT2TUlMCYFveBXzKB7qSQhPJPV1iM25Ei82F7Jmt2X7Ddc3RYu0HoWjoSuU
Bcx7dPSU9hML+QbnwLYiEGhu46dm77sgM6Bwpw3OFwP9V5aViwbtroI3UhERgf5K
P01uDR1PuxITbHXbfFxJU1k/FeVQI12BkXaWrMd1Ka4pIapDhea5ASUxxVjbs4Sw
EHGzcgr3NDVJUI8QEE+d/5Iicc5eyrgaFVcZwcONBCqpmKuzQmehZltp88G82DDV
5KraReKCf6jZIOlQ20lYqoHy5nc9uqYz3CUZ+OF+8vUYIfArgsMSlCuq9dkVOjs2
xrg3m6K2Wqbr566t/fhPjrswdlofiu6b6bylK9mIEgbtM49yx1amihuQNEQGQ53e
5N1opGqB90mp1jwGYmVWjTAk42aVveCLJQPcrcSExlEPWVRuQ6y3i6ELrhi4XHMe
NCEljbmNc0kMsyP4Bjo+GiCq/fKFGf3Nky/qrN17jXpxpmer0ma4rlRI8Wzagi10
QvHdMSYdCjBb4HTcKQud5BlOnISwigTIf5J1hsOoOmzMcRSt6RgMcCUrTDbWP6oe
obDWbWCz75ynGggc19VUdqxwu1uSJgHD3W2LXZj0wOOlINhfrpRJMyI9tgOL2uV6
3hDLOja60uRaBexqfZwX2BHDdSrlfN51MxSxHkP4GqgwQAeKH7Y5DJTBUYCl2hA/
X7RGCpnIThr4fwCbBXwde2Qntbo3JqDLC2G2BSXpo0kbdBDTITF2JbU5kwQVIzB2
niWMKe8mSD98jSgt5YGkjYexXbb0iV3JrXZ/E5eGF8W+R67DXBjXKGZ/i+ZR4+bZ
ZOQjjt1x10xffhilu+07l0WFYNSRE/Tfjw5O5nKZ1Ww97jn+4B8oELV9Qh3NK/JL
4K5P6b7tNkyufeJ+tAyMq64chOtz1aopt/nc0fABRH+bmR7r1JM2WLw14YtPU64w
q+Z+cKlqrqi93pIg0XOw/W90PnJgq0o1LzbVlr8jdWyYBgKl1DkFAg5QVWRvCWUa
Dan1pbv4BfPz6SieOxPzjVeidB3XvRj2hjbRGh6KSuurvzfit6sqdES1K5wu3RC3
yAJTDTJK2c9Ab/0FnUFIBNCXKqbwWYsNc3l+nllUt7BX1brrFpwG5NeJwrWcqZIJ
JZwGo5HKChYP7GYMabGLyRAWyfQtUEqhybw2rU6NGU9P7gaznZPgGm7ztUJFi7gS
opwj/Acv9GIOSXqr96lyIB9pEdn/yyaDEwpwgQJN6aLLIJwVdRQEMVqb23hkhx4q
uo7p03BzLXPFw4wPdaHFYdlCK13XfaBSjYYBKh2CbKjagt2Tc3iz6bj9AOg0RCm1
Ea69a8hOeX5Cu8ha4gGqg+Rbrd8BWv4nDPH8sUzh+4qkGnCTRRHsaYoTSrP9bG2M
xlkuhTIfV2vs151bCBMZLoQ76Ew1bFcfecK5B5qxteNGk50vTgt/BHqsYARZDxdj
xods3rIiZ8+4FB1i0wXjWR5S0NX5sv+ESSye33O2iL5c67SF9Bn5e692lQYvD+pQ
xKMeGCSgGUdwO91JppGk6NJTVLstOrY+XAaVOmnw8EL/zveVWVRfXWtzhK4RZb5e
Xrx0bnONwbvJ73MGr423tkO+6hAOt1k2Z4nbRgKPXkrqbhLTQKeCnjCtFtvOrKH6
hCG0UaySyaj0b0HwOMRWW0/+mOmexKm31VBhA3y7uh0hLPiKaYi+H5yR8dyOGuO9
daXytUcTKQukQh5Bw/6bQfdiCgnRmnEPdfDw4USef3JS5lhyi4AS9mlWuRtguJ+t
N6DGbqGnSaAZFTZ1K6gtGF5ncuuWr801jLsWFjDs4pz83IpZ6aKdMZCG8ejnMFuE
byiDUgaUWGD4Bk+cvFdFQsFsQsiccB1WBig7xpoLhJvbiI9/Ed1FObtI5PkcG3gf
9A1/KACl4s1oIEPjTCX6rPNpOhrE9qIa2FTYqedqCrrd9G5P0nFJtUL+/you1/2h
nDaeD3H9Faufo26v6PIz0QK8V67K01zlnDWRrrjRznrBtUYtvn7vp91kFP8p43R3
f1jazf7zgBw0XC6ZaVHnHp0eSwhcAHCrTTsTAvqn8j4AB594gboCD6xchJREmweM
jOOxxw+zZRX93cWOfaAQn0+3UDoSEjGBqi/JNbk+VcrQ2ZN9OMFEXXvCcBvjj4kD
HJs3XPzPWae42y37grNW525NrB8CdU2AlwVNj3EGxNzIBigFZfiXq3g/23cIr3xy
LsnP5AFzieVNC4M5PrEPdLYfBmnJROcijr9aOXBjWGqyaZXFhJzUXEqRyDz1AUWT
Ke0M3BoVUBsSQF5ZCQgK6z3aCZvs9b2Vvz2SDKq64nbMFasL3CUnugRy6n8SEeAC
/Q2SJ9XEvMfh9FNEjVBA/bKiYh5/BdzQiU24Fc3FLstwDJFnzbMSdaOgKLCHLhHN
aNj4bFs6DCt8JlU/7NBazM91x9vYuBb6FyJhHkeqUHOQKSajKqR5u2losGCQdCKZ
B80ShkOK3fuj3M2gmCm3k5GPpfDCAKqwsqM5EzuZ+5Q5OxTY8uo/CL3mjJp8H9+c
9KB1P3GeAr1B585vV9ln/L7Q6ZsqoTdHBaTvo7LYMdOLfo/wZKobz0jZwHAOe35v
JSCu4Rt65qq5CaCx92fKzljWOMHTfpEiWthL9+OYwVtFLQDEKvs9f/nZPO5D6rtJ
O7FBTemZ0TxFBP8T8LwPPJEMFybDpgIZCG6xaZUwAyyYN75Id9m7WTCgGI+oRdP9
gTX5RRkBhKWT6hQwXX5tY0VjjMfKx05TywvcXIHe2uPmDup+H83PSYUomM2Ov8a/
srdsKNZdcybdyZoCCcubQxy7WetiAGGG0ACV70bWLcOyjpuHoMtmrWq4MbxT4JVV
8B5bCKtVOr/Y2QLGQipcPX6juJE9nJKycDLK+9cePR4YxVR1rCH4kSXvZI2jWW1B
Fq8AVnNTb2qzs5qmM2AWMx0TfnHkx8ZLwgG9iRQuM3lgBU/lm+ydNFvmLKF0v72B
Iuy94ekPTEzXp6U0c3Eo+BBPyPcjjfZmTNtDOlLNKtyNDa5Vi7gUTJ6IwmLl9k2Q
cUaekEIr6LgWZWCxIm3MkqLk7RhAo1U6TR7xQSNKVUHmYp11Z8DX42nV3w8pfbrD
Pv5k91C4BjIlTMJd4pE592CYiECipoQ4RghDoPKFPa4CKtKYv7kk/qPcFNYyJCMa
AqloxBGmefFHDY73XJq+lIzKy9K9m7yZ4UBGWuSKkllGAOuNdpa8zalQkSjsl7ay
sHrSjdZ1yvA7DdyZM0xggcYWODsO7fYqqn69/daj7Qnw4psp8gniKljtOfgdzU82
eDaGa0fkmH7wAYkjgmSW1vMmG6OK8QGQXxBirFbrZBB126RkAV6EGEBlNwghUD+x
7GP0Vbfpf2IG7V6HmgszNJsLIdEO4xeANCe6XoUeNV0X7sV3fnG+cJAt4vPMfjv2
Jd6c9YKFs9yY4ZIBpfZ0sPECWbQwepihs1rkwYqNm1HY47US0IB4GVtaCs3gN+tc
JjydIC/GCIhMSSKFDr2Z+qYPoNoq6k0NtbcxFm4po81eNmoFbWteQy/4ehz7yCSa
cZygXqy0QNcrrGyA1cuFsMDMKJzCd4Tf2RF1GBDAqfDUL9Acv63Mp+TPswCvKhJh
swLnrrKPpXXVStMMbYonHKy/0zaffZBW8MovBE5Xzkty6al///ry5k0hjHdBE2ZT
uX3d1nlBD+24a1h+7+IxVHa8BPJiyoko5hmWZedzjyD6bk+8Ym8wp3Flr/8zTHQl
wF5fLFr86TK4z0HsHTYpOE+Eb+c588aH3z/ieFEQRa2YxZpemCTRsfRgqq/Rg42h
A9JGsxnsQNjOtMVEUVj8Fh4IIsc9FJzDzQjB31Sf1kordRsGQiROX/B1IvtTyvxv
Y98r317Qwh5K8Ymt+b1BD0oDTNWqnFxmOV5T2WdC1LMtImv2txwupK1htzfzv/+G
mfVdC+es7NOymlRiXZdIDURjOV+L0w7/ym2uZpMXcMn2XvaWM6JxakIA8m7jxkO1
Vp86dQokp+WR+/53R2MbM+9/Xjn+W0qLs2MrbKYpNh4QMsyWLZvNpubU6YmGM9FF
ZN2aAwV61FMLJ5PHXxzGsHbecKOrYufFjbiyA5eYS4in/CBnPg5KhO/Jixo8ZIV9
Bhlv0FzSi99X0abYzbBG0ldFt+KzpY6K3HPWgF+LbWh30DCJjECpCIW02m0m2/UL
FxBEvwd2drrLPvMXk8llR5kVGntLnxstH32HFOQwrwJA+AQ09rAzDTtJJp6QYVH5
ms0XvpAdXTRAWjL6BMacKnyqSQIuzlo4nVmmk48cPeahcGrEoNUnBht59zcVvakA
BcanPz/EBSy0ioNgPrm8uD2oKJhL0GVc9b2gff9TLOZOiZjs7+s0wg9JlmUWDOWs
i7r2KvwUryUMh5lsAWeo7k7N8+lhh+kt0XYEX7Wx1z9BUPUeoSlFpGxuAFUR5MOk
BfNbQODOHDdAsm/H/LL1uBpAgbLU75/gjx1OJFk8IIWaYr80tDSuMyyZDtT6+zKc
d3HbTFOoA23y63CuJgagf9lie+J2AzP3Sl1JK4nKu7yEGf2Wt43EHz9eVj8ApohO
b/YNdVC7P7gtrtQ7RY1tVDYh5ZxvP0jVNJedzbYcNa+VaeoQgg1zVXgd1w0zV11c
X2qVghJIxLioqrjKSS8Bki/J1yHHQvKiQ3LWz0Hz7Z/QPuVqWS9XeIFTvTQx8P/U
wGdlKiTAwaNtGDBbq9TzLOtY7hfuWTQJ6OlFwCxht2LYAHdZiLgM25tVVHkiHCxh
iWH5ZmJ6Y2vkD0eoO++pk4+E35txLHnbqp+hsiiGM8hfquseTXX2HKjpanfnVrX8
3sAls4SXAeuMYqM/RIiiChT0qOShxQkzH/dYfqmBPVTVwR2eZfjJNJXdB4T32alD
L3NKxE6NzSvLni55sRZvPXFL85b34h6atIZU2T1YigzMVyChDkvnc1YKs1wzVg7L
csr6TcHDOqQp6t9AMdBSKVNqSMZhibq0NLUBs1Bs85afjMrWwB2puxomcCOUDHTc
VlpZpOi5r3OjqLc6YsC/hGsYtG/MsPlXCMiXKwFw5KQzRVJtsZ3z61o+i7z2vJhk
vvuRHB2UOOlrB/sXdk1qbcBn5u+93UYj/CQpTM4R/oSYWKIEoP+k+xj5Xo6ademz
zMsROVBvIKm6baLXA0balhKoVtF3PMramZxNAO9BvMM9QkP5bbQwlSdnBJQn+7Pg
4hEqre22kXxBMInba5qOi0AVrK7tSH3I0aevUgFEhsEaqF5x/pj0El45ARz5w1gN
Zjtid4O89Nt6zsvZmhPeids6Gakw8kx+YRqNaZ/dH+u/z1pTQGCQt9xwjKEBYa8K
QHfpejVdn/pr2aRmiaUym93VamOEdDFdRCWHXgUvumYEE858/YxiJE4zhOEKdmr5
BmyCA2IHn4LS8OwVjfG6HF99Ug1BQFLyOKfAjdjMnwUnTZbg8QITvv3vPAPL441F
p4bXhzTzEdVX+07O/Qx+XNxTHSE2pKsabkmlcAa/3nR1fJd4ef+h13N+sSTKn98o
YOLVuAxIzcpaBrARDPxh1CBRLGzowN4+vYeRpo3c1zFDCxREytsxDQS4PzF6iBTE
+7sv1Srk21zbRjG3dCh3nrGH1RwQlp2/glagCQNpHEmxLQSkYk5DMPyHKCS0lnn2
M3xZM10IwEVhfLbVSAuwGV43bDg1vaoDX4i4v79WFdztsm+Ag1KIID65vOtEG6bK
wcG0MPwB0Ni7w3EUw0pZhoWxT/skMvhSygBvnNPxlY3/Ker57GrKQleNaGooGdjv
Kxu7OIHAlf6gSWa+2zWZ3y0f7MDY2+rO6U8VIygimS5VU8wceYLMoSJahMNbL/GV
JHerjO/5Z4DLIMh01DrOstIO7vZBLfOzXp5w/4ENCzP5Jj+dYHSrUt2Njyk8tsI8
QyUYEVvIbsGudC0T3UfRTSpl4QRRdHHR9ufkq38yvdSpB7R16DgHuHH9vJ2+p+I3
nJIQX2+r8UiwiralX1HMFMm0wkjpkx0sRgEWM4MwMMl6+QwKaGYxDa32T5rdzxkD
CPqTKqzTdbX9w1qaf4xW9aKNcn9J7Qnwt5UXCCRTHa4IbC3kjzn+WXd70kVRcyU/
njzUlQpYDE8rhMoXMETAospeW4yBULhKP54rUWf+tqqm9tF0/RiP7thlkfT94FNk
r1ds8BUTnGzup33NkD6AoHJGdzy/8fNUydoWykqNq8fancJfi4QXxbrPpG+bHMQE
Q7FJUXEye/mGmHNY+k/nLxPdp3gxZDg3VJVi/tplPQ7gC6s4gB3UTr+3AbOG6sUj
Pz0RSK4WC4cvw8PhJSftOmElz3atltwRhPcvE4q/foCwhvLt45Dw9AFzFl88Wg5m
5SK2kV9jnjm6gYMUqb4O6prHPLGpLd/UOyeMDhla4xw+sxKW8F2VUzJJmdEGaIhT
zF7ftjIxKoZPV2oMl82li15awQ51Nn09KTv1t9UyrHuEEH3hBOT7QKC38SYm5rOv
BjaneVvjimvEFisRjQ//qLjgO5B2u9OmLXpE6ImSaSy6L/6Gqyug+65QlcKjfHqI
wxT39FhepcuY5kIUMKJRQbV1g4kxpd3OxR+g+pGIQZ1reS0bP4KLYaro1lV/MRjS
aNR08NN7i3dB9n82JYEdujs5m+8avpLGvuqAs3ZBtmvbNth0N23/MjsbRJXdNge3
5Qnh73a0Cs94qjKNrgnLDkAeTaqC/2+H90dJjMxh1MXApp2gau4XwqQeV/w4fBms
U8SfcC7JcUWeIGJ1kXhUTIP3CpmoC7x/QlfsW6RhFfHZTOIerazN4WaQPl6Hwfy+
HrKLdH2L3pcSYaVR2geI65TRcXnjtMWJ1WCiCzGXu0BS4BCK8lWst50cwqkcWibg
h8Ra2E3XBRyuPjnsfAUxisOdj4x5cmdohSBuY3I0m9Z2xuiPyueij8HugmBIWGrX
Pp5+lpBLcq8Kxvmmi9lnmcYbqm9jjlHSdKZdwnav/NsJ7ibehX/Jfrte4hC4JWyb
5yIja2B/HS7w+A/klZCy0joPvxfmNN1bFNi8mXrCB1u9quDeV9RAhY64kKkTfoZQ
FxW2OrRBe5NjfpLRGZJKHjzhTlpBSKJSjfmH40SQlFq1J+XZl1HD7joBlSFxgMDU
yAeRWgz+couEeWHpYFJGw1D8hXzg0KvIrZLk37IGBdrQKt25lW1wfSU7P4a8ljpr
DKXu7J/0G7N6mue6XNyGBIjWEMJpZljYLvpgK+5Zvyl2iOq+qUwliiakYbFlT5Pi
O9TXmXuymdHfIp89mq8lv4XodogkLXhGFfHOsDWStJZl4XmC0vISbaVfDN/SIx0S
0NnVKBwQny5FLb1be6N4rG+nEDZxy5y4DV7qU2KGdToGXOuYDCiciguydqIZeoZm
90b5ZryMVGYF3fl3RArSc4mz4fSoNFaWgr5EFgic/TuhbRQFaDeQm4Jk1c+h02Sz
NfbFnqmwAEPlw5Twy5JaJ2nOk6bdFOfHO+4PP/8lIEZlDHR83AxVCY4r1IjbNu/u
d+Ah3onec+tcjxnO1qLiJFMKzaZX7dY5QpfBIwelvGmKxHmsLs62yAD96wocUOnR
jY0bM2bfNC9LmlewsUIrtVya+3IQ44GZRypw+R+PUP/CNXusDCg5/dukfOBZT+/R
ZOIk9SULxsRGVDoE/VK4mZijtNVVUMcY5to11PBU/aNzX8feSwVav7vfq97H+BCe
QX823pJE7MI4auIcngT9YbbFfLr+SEq+1YLg3XJ6Tq39R8DaNQxDnKaTpOVbkJaz
h8tt8BW9bjoPh20MBJLK56CIoZRk4pgPMEJcmOm1UBsC07qO0y56cjhOKvqpJdlm
upfMW330XXAOzOedudB396n+rm2CtB/55IElafXgaFLylrUJ8oIUtKAxMN2LCbNx
fSGop3mFyXeH1uYIcLl0aTlU2nFrYmkC3fKzn6wiJIXlPPj7bcPU/AH0CnqUtIYU
/G2AXFABD1Rl7Dwb8QAHQbAdHdmR6Tmpxf9s+c9JjQBDBWBd0EhuwAH7bgRDIUB2
XdGRVz3GoUoHnRC88QXFzlJiw0okRnsGn9UU28+wCg3zaiac+dytX9QLr+ZArQX2
EZbaNAg2JW2Q+S4jNBBB/MIDzbBQQ4BJFa3Wgc2HxH49yT2ZYKGdVecXKzYYfHeR
xHUNwEvYOFcxPQDQmwGTRGc6K8FCHIeSSDivLCgm7xRKKSWdUuf/VnUSAchgoUV+
FkB90GVGs2tvoOYKrEute3i3YVEruLCv+E35W+5Kf6J/T+Xe4bwhUvYvkpJMgfdV
Zm4iEhOiLw1KKN7XuziZ7miG4QVdIVMB8B2Dj+8eU6RMZOW0ZzDHBnD8qO8zku3J
dQ7HNyv4AOt4Rjx8Xj3eb3ThzeDRK7eFUR6NGTkKOsr4jnMeMbm4A9DVHCOH1NRg
/BBckIouleDDkg+vVY/2QDlF0fy+EGX9aT5vnbMjge3PIyZEkIEpy9TYWx+lKT3n
BMx4uaaMoeyuuumeMEdt6nrNGudvTMbZnac9ps/DMeFXpxTAo/cv3o4JiwLVt81N
SHm+m8cvDT6wVjbEWEM9e4ycJTewZ7ijjV2AAeqQrtHmdpNQpMindrWGVyMdqG/D
CK4pfIc0l7UwzFTKloDUrbX4aBX2EUqr4LCRmQef/s/VOjaf3ApWla9Fa7LMaPwE
9ZpWyxyTKBmRjxCwv7/zOlrIPD+9Ws548e9m6EXqVXGARekEGJNR/Ns3R1jFlL5u
iwncoslmtfvMayD2Afn8wiKw3bJJb8sXQewnCXSgfdrUMq4abw/1/YJ9ImzMsSHm
R7S5uQTaytCq5tCRDbHCA9SIcZK19ZT2oX0bDEpeFmGZhijxk9s9BV6zD3m15KMQ
6dhdELkoRQute/CdrH5eYu4ZP8ViVjQ4dBl23rmSBTq38lvHq1yk5UI/OuoZxbGR
LID2V+O3mYY+1+1Vosui6Cgz3Liwgw1zUC85SLaiBIbzZj82id+bPVhSWOnFK+Gn
4pAcISlnN8ymLdGOmPn4ccYaoB7nGWvST14jmZ/6fbp1m4Zf8rla97aFGh8eebKe
s9iJ3T1tshL9VwNqRFYc0uWMy3V6s8z59AeHeeZweDPrKPQzhsCh+l+lY0WDGRsK
RMwrMa4ac/9Bxg1oVxANldTtkHac0nnqIvDyc+2z+7k6InbPotGSWjob1fFCmQoA
MwOziSNc/nHkh1xThH082K5gSo17fKIKJKEYu4ZN/eh0lZK0QUBS22fXK+5N3yv+
SiIW4k1bXFpJ+XHRUjrhT5FFTYBcOxUQ39Luh9IwHalRqdEm6H/u8HQowER53pVK
Y4okI5EdtS0Y0DL9UamZHMvNXrNBR5w7OKWsv64TeLpaHr/TmY/E/ogU5p6S2NEM
duH6nb+iRvUeTMyP88sS8I1IMkcCPxiCYDff/cHNxdng3uEiNODpiGsbZYm38oCo
27dmRZ+iJYmb89J2St+AocVyTx037rby56hRrKxiYBuBE34yd6Cx5x9ZxGND3uUs
XqiwVhW6mKu2fcfn7RmTsoXg6l5Xo2K0IernebFz34v0A4NZdXRUUCX2+wlBNtk5
q5WIsQRv+LEqs7JC6AhOe2bN8cfD1Q70vGVfuaG1KnIjwO6xAZtxNHsm6lsViUIb
3rnj4DUuSzvTKd2SKUaQopKiLANGlgbdKrzgPZj84sksWI03WjIulKYkzZD/E1Ve
0mA20LlIDXfg3Kd2Q9U+zYn+GbgE3IO/YW9/JPb/9WkhcCd49LUrH/LkCs09Rx6Q
qPOscnTCCBcTG820IOII/lbssh4FVZu/S5VhyOJY7uXxqPuLxJraODy/7WsILTt7
Mv9+s5XllCnibcvGfb1ZLTlQvOYwlGq/xMHe8sF0YgLS+PpcfhMkc9CH9g4OO9Lp
JBcA3JExwAB+FP/K346gPpiA17lFW4rCe6/ziUKvREm2J7/kQK2Icdd8YNJ2La8S
6vuGY60PtU98Ijqs3CY+/uI+DesOMV67zybQoJrxqF55Y9QSJ7D4TJwMEfVCxFHn
vZ5gIqjdSYp0ujpWlFatu2mN2jlWPCfX6dhqtwBHjxZUbZWlT8I00l1U372YJ7Zj
9RCKPGftjtMLJaVY8XbrfJQajOHl+UpFntlQJwkzYC51WXyMsTJ0foKLsT6EMcvi
QOSlIZz2sBUa8SjICorX7nQVhwNXeMq3wHnr3YDnjX1IWgAYXsjT217M+bJGt+WO
mOOP5Bbo2mtsiB63g9nShmTjuy/BWrrAPuzWJSiJSL6p4UbxIwBATQ+Hyhhf1ffi
0eGNWQwtleEYp0jGd3PXCOiEMr/b+mO8UR9eE3Ie8DsK726l9ZVJNLLTWU+fIs/d
ENU6oOeFsfsPksg2VNa2Gt7pzp5pcjk7rALOxA7MLWuucZtnhgF4Oi126MHp0Ult
qfPtVKRjbVfLLL7gxBS4/eQnUHleD5LWBar9M+VYz7CTh5BUsgjAKXD2s4mGwhTR
qZVGoW64R8L05E6w8cpJdzXz8+nAiSfjwQTBTMM8UR2ZpCsNnF5RyGIWL6PpmBH+
DzSWSIx/Sn9KH8k4pE5s7SHoGFs4CmpqwSLgTdjwdiw04/wBAKPIcIwf2utiZwPJ
pD9Cd2cS8aqy+Un9eIBMKwsOflcTO2JiLPPk00Ef+ArznMW8yCWEoF4eyd42zrzc
lk79KTlg3Uvco4f4MwirH1KeRLVQfxJLpCLm/pFjKmyJwxlnfDmOrDEZANiMQBCI
NyxpC1YcXQ4R0AmPf3teabORvFswL0VN6S2bR8uw6n/wcZFm4swaeDj6uwt893y+
u/D5+UjnKcuCh3hlItgn+40OvLkTPpJgN9YYLt/VMevXKJlk/pLxEWQEzZWePJ2q
ISsKoh3oVj53iAiVlMdUBRSiynPfxEGIVTzQFfCkwpl/g7TgI4Dai3hz0RjBD9We
S8FN8sGlklouGcXgkMkyuZxuRG3hChMh/8vaWEB6lmVNqwcEwdhnCXzVYAxdo3m6
xD6ZhUgACh9YduNoHHOl6npcpQIDcjqlMiysI6JucZaBjyrCUpLMyDmWKq7dvXQo
3grubwj1e4ZxhxCksyXK/aRQJ0YLXwF/jbRQQdEX4UXXM2V9Ia+Upumn5H07cSTW
fO+ne59Ybk1R0aC55GvTsj3TksR66mNkc2fOMp30cxTyMLTAdmu6i1t3wUJfAEno
2YuuSy9mTMTpsRlpXWYXO7NoM6vAT5oqESnppfxp4CZCoVoPeF+Qm7qNpe2C5y6W
+EiTUOPIK2NKMNV/AVA+gD0PE/R5z7s9VbrRRAKhsy93SVuI4mrUsZ5mzLcOud9K
R0T2FXG0kgVbfF68CI8X1S9fKRT0kHS/iCQBG/8bwGFisrr7BaKaLjOq/N0A6uzh
tmpuYjp7KOTsIV19OBzr6FktzUsTWZzLphg9agnli/6yKztrVUZJp/EYl64pcRCZ
r/W25fxh67xmvie0S0vJjWFk1ch90ubg3JXHDzplo4OlMEaMGVg/XQWq3oqb2L5v
Gk5xWiQWEeznawLXjRbhIL5YxmDogZ8j0Fvx5lJmF1w2FCPyjjyQoJwlljpDz/gb
k6OVhFBC+uva6BGpEbT9v54cJvZPRzQEKt4ectI9TTmFHzXMDRrkeHSLnZjA/3wz
k/UgTngbnUVsgJTyavQaQJBy0dkmH1q7LyvO8tjF47xNRMEFtR72qAk19vvgiJpZ
N5ukJnfZAW0C4oqKPIlNX5rXxSHEzxNONPqJKPWHDPHPED0Y1F9aZuZhST0WAwWX
M6J+10KPoVPYCkMQwcPpvZLkiS80n3x+YUHHLtClr4n8MzLfizOT8qATBLV5KNAn
z2MDsC8i8oRhFrZtDwCH4v07Rb1nPt1C0b7lFpV2jXkI17gp51kUyrxSjrnQelXV
2vj7dtaKsWt4Ox2YyDumJvzbDscXVxqu595cYF05viWLpK/MTpt9HyN8Jdeq/UTu
bErf8CUgX54GfDNE6nUK8mXCktzcL/mOOmuD1vC0aXimhhQxBj2vAml+vJLRwKMI
nW1uHYOc4zn0vA3IrylgEM6mhwxaAXN66y5mMkkX1uKS3/+1LVq3pNngS21u1g8f
VElz8x8XBt2JaieNSDYqzhDr/WS5Bd56HmB2XySkgpDEN85bS3i0YonleBccGrVw
6KzUhUfRHZhROZt9zGzx7GWm3WUPsPdZLLtSQEf61OpRrvOt4LsrHAcVRhiyFzUi
PQdf/8nMf7qJmLCr+2y717R4gRwLCI8WnQkJ8C71PQNU50PsgFVHA6KYcqw32ASE
deaT402N8iApxf1Pd7GhaLn4EBzIJNeNZ9OFJNKJlHNFpoVU6xoTHlQvCbuSDDMs
NxSF82Mj5f9YbTIkAXNKoEtgVr/yQJi6UF4u/oUzhpswsjZhTH5MSFo1c3rknFee
tvbno2IRmNtQ5gA9PaEZhdULh32+B4Lh2coxOxP30hGqDyw0f6qnOCA+iBnF96us
qAo1lpOZXLoP9/41r6lh4Ks8a0+N5y4lkLMCCa7CbEL1/YS7kw4w9ZLzcUhmo72C
z3gnboUU4V4nkPD8PdH416UCZOb20WiiBf0jKccl3Evhq/rpQCDZICz3PyO0yxwZ
jkJyh4JPQJVfOL7Lk58SJuF5NUk4p5shYrS2xaejmV5Nr1BxMrWzLG8ghzSWxurk
wK1y8QGMqNTSizH/jWsNRzaTsvpZU3PXvXxQPeTrh7bTTmgP6onf8S+9SC14tLqB
pTKDqNjN47l/LmRx5v2ZAcrzyrr1saTD/igkioZnK2lGcOCr3tPTn/1gKO4oIifH
O0+eisgankk+8sy3LSDQvzyMjkTsRbW6I5w7foajRv+tBt6gPm/uKb9PT6aN38nf
n8FNmNfjQn1xjz3oZMl+yG5A/IB9bS9ctQ6ZW5MtyHg4tuN/7WX5MmRH+TgqjB8M
8cQfUyUh3NcyJ4+1RKuCJu1tfEzGlBwUtqD/sgkWaOxHJSR9Fo67RmNO+zC8srYD
/sAuwjp92bNR4mSNuW6YQY4cSviEsENEcW1BsvT3VBvHwyhHPlbCG78LudHgmp8r
uJgHFLn3w08kc3e9N/s7809wluWH8inUHvLPu4hJ3/gGPhGdkcnnhwnxKyty5Hgw
AZbghveXrS2Ecv2yvKjaAakXqs2c0vZyjGImIuJ5zu9JKv8c2TW5hCUPc0kdlrFr
mqsf3EWLCalGvC+bF1SyPIFa8pqVveA1+wtzsLGDzWLtUpcO/qsF242PTVROhRx6
+VSZRlFnOsQxgCVoaaBr95zO12rKGo72Zsm/EpfAVZhLAnbZiTfVOj1YYDPQG2ht
K16IfueIoDdvLtiV7QQWehbxlaeQNiOLeQinFgJIoIJz4BxByfDGeuwp+NdNl/U/
oA3ZN0lA6+pk32Nq6teUXa8qgH9J9A7yJx8TfxKTn86qGBueTfFzfKygVmmoAOwA
/G/JOeHKnFL2IrnE8Rm6ciZpCaGMrEPmr5+MdskeLvrJV3NI94HC0mNPex9AqJLb
Ty90KilYsR58Zoa07huAzVV80mWTLpCtjYBQRh7+qTxizhGX/XN6oHH3Fi+u8KM+
B5Uf1/+8Ksc3DmXRNI6O+1tsOtx1jNzqOUPwH/0Mb115jOaNQepn3JC36D5Bp/o1
6T/n73kbw1jIhwPd/mAqT3Uc1XSCHHS20mtacdLTjrcNi25LsYD4tI/8x20CmOW9
6IAWgy+PpthdvlzVZL+8ewAb6YgX4DYkUjOPPc++/9FBlBBNM6zh35tXmWro0lvC
sT+g2lvTby5vXHWTLcpyVErQ0zIydiNpNOi9vlrGQE+GBS6gbh8jMIYGOwKRJxoJ
juTIFlnagxBbXYrlHkA8BdBT8BORxx5hyHTvFO0ZRWBwFBUyE+Al5LvNi+KhnvBV
xn3aVx1gM5E3WJjdmzU68DBEqntmgJOPV10n/GAW6LuYgxkTJBXDl5NrGJekZd5K
JiTP5h10iKn8RumBChdd3+tTj5QKn/iRGl13dXf2qlwOmBvMHb4pkdtCHD+l+yGx
GQZmYM2wXgbDMMxEGPpdLVmsayVVh16tszyPknZy5sU/rC3/yItjmKeId2VboskD
WrLtQeZbNTlfPNP9ijZIAoOYnpq+P6ftw+8TjsvUAWBMMVhVSQ0lhM190hczbBxz
nNgc/lAe5tvZd/fPV59iUTaslfO0Yo4yW45StPBHaeWefwmb1QxpkW2NxJfoOvke
JKkeWE4ebfUQQ3i87dCBP3cBCV6a7YPEdAGP/ldJp82BkZA9eOUmdY/gyIsjx22A
7XZhlCZ3nOfVJ7iPH3Kjj+zbYY6DWh9QWgDwQlJg9BvYCTHJAvw2dFDjQkjkJSrp
Jfu4+lKawaD/ArcL1YgQGWLeznSRUL0CUCBZjnA7QuV4Zm0gc7DmYwx1bzf7p2Fw
ov9Ssp/xIxjAboEsqSFEGoshvOBka/11ok4pi5T+AytStMRFN1h1cGIZR50iBmDN
P1v/a0DtUlMx9T6SWLoRIor6CembdHH12ktP5dfIJdMuGe0/3MvTKISl5Sb9wk4+
+Y7/dQRk71t+/sSt9oc5W2cVBswSNoKrUlqsqJM2ZCA2+oVonBCMk5Z/HbSam1KK
xqkq5DjpNy0wrOGKwSyFmYdbYxem8eIq00h8U9j6KoDKANHiHaazp7HXx5DBIflF
b2oGF9/u/hRh0ojIrGU0nM/EJuBgtAvu8xjhy5wt+GlcA9tCCWv0uWdVW+zfRll+
ndnxqXUQPPEgr1eBJhyPqGfqoFw+I4t44VTXR7pKAXPLJPkud/HrQ8CPZKCbSJJh
uI6HOrm3fIV6Oqc8JOXr1xbAiaFl+8/hFcxjnuvYDvK9EU8X9GXRrwjwHSbS7wb2
PMVEi5AEU5ZLjcsZYTIsKHh6NdpDtuCJtmmin1+nlUx4xr0FiyGcSJ8kxYKLWwE2
n3jD1JHu4NiIE6UkAuatXBllgbI87i25wUaqR3ag9/WrtJy7v4knEtxfnjitGyPd
U6MbezI1p9RJxuZkdlvWuF/An2cMbUvsBkhqNdLqYrzCzetdVlQbRbUkqA7HKptl
gRZgzu8cPobv9fOqo3aor/YgC7f6Ixo0dWXZzYMobcKZjcMZvQN4CWP7we3xpQgr
IBx+bMQ9elepAJ7a2O5UluV5T5CB1RCN90bS+b2W4MZD/3XFzqFVPdpNgCLEK6SS
RaOzOTpKwrGhu6EuEEu5YZc6NrzhDjAoCKizj3Ewagn5EjdVp18etrkv4S6lbIOx
JNvONMNdiClSwlf/CK5+PY31VrWFZSNZk9JHfdeHS5KA5WWHlWwvWhutAPq7Xgj5
JVyraTRLrxh3o4HoyDSt542hv4n/EGFTzGLFDrzEr6EbJlHyosh5Ct3Hr/xap/3t
oDh01gfgoH64tOWa7w58u1N8OudrDav6XIEzx0aRNIBmL7z1mZ6qOo0pmDGHqAUR
rxcAy7hB9gvK7QdDa+og+dpwDQbTZQIIFZWMrV0JU9vJlBIcl61eqcPWgdY1ZNm2
P0yf9DN8VJC8biw9TGhXiimPaxiPuUyehMJYZl3o89gpFAsZIRAO1VbKmQ91TQEs
gUdVMeJ6WAdQWEG3QrRdP58ZpxgzTgBrP+yg5X5W4VClL9rvMqBEJnSBghhqpoLG
D4xlwmq44bXabpniujpvGYp5Prs6obSH2o3VViY5oFVg2JNAY13lSLFfa2kOxy1j
LSqXp4Z3cfcE7PYqc+dsNaOhpxJDAnWamNpmk1LKwM+yPHxDLVAi5sx7AyKj4Z/P
XxpFKqvZhldHfUnIcA/JLaf5M9mdUWM//B7xT7QTuoCCLRb2Q2lnUyYnQQHdG/Kh
CNo/nim8H55R8Lv3xT1QKeSoj92ML8ezWbubtt0Sibg+1MHslBFY3krn95zSDzoq
NQU7BJzwhwCRPVcg5E6H7w8g2TEA6TxP1ft5aSnX+emgc5XjAuEzEzSaYaiudtgX
KThs0rgY8PlhxkBZkuZ5lIN0y8d2HAUuV+wHSKeRk9aAKpYrE5glnQ6NLijPFVNG
uLTExm8gAZb6wjZFRFwkdMtMhWC2VawwpR0MuUL5ODfUyoL/8bV+ghJUVZkdZrGC
pkyXn3K8vIBaBpOVSPQIL7CBPNZzzuvJBbR+C7g3Bq1hIhat1j6nDydVaQFdrE7y
Bju9/w8Alpb5Dedh/VR0mUJhikixJU/K0rwSlHD4ByJKzi2rq6jICdkQwpnMvKbT
ArniHbft2qL+gGAeGlop3Wxy7xI2uYHDcc6Ds5zcdjr0toWdIu+qKdnEfp6wWqpi
82sCi6yLq7R/kHh41pOKt/DeIAeQloewyO4dU3Hl0+pS0nlLWv9gJ6Oni/gYymLY
T1cI5Mf3oROWnhn6H2vWYo5MjidagzoD85fi9XtMBp/K2z6S6qRcXaeYR2Cl8cK+
3iIwZ/IyeraIZWBePQo71Gu/MVbEfeqiP0+x7twbto1iycsPPjiEPJCLjMiJVnln
KgwkhNTUE4O2XggP6fj9ZxpFKxe/S3imBEfLN8UZRE4rO8kbqcT8A1mXuvJq3SK2
oBjq40/JW973cnhWi/AymNeyXJTELzFsfQz5PswvAOLwPOSCTi+Xdc3oUBCA3ogw
p679rOFmJU3A3e7mUOSZqsdl01LaKtCscTM+QV9lExUgb6Dim2ObsoIS+rsBrOy2
exf0XBDFIlIaxEJAbNZtMWlu7VJ0RKy9U0/hxIAXbZcQOIPD/poCUVgeDO+Hw5h5
80zP7a31n/yfrZOZMWjR7gw5Rpws/JNCI7a5TQJmuSLailM2vfInVRy99NlfSxyt
lffhKOhTQJeaCmzov6OwvEuNNW3IAYS0UnmXH1PqAjd2BK5sYo0M0Tc4NgjgveHe
OrcMtuYNu2sXojSf+zyzsuHh4p1wXPFhKOxb7g8nXk9udpJPrsLePoITdU0Akvm3
FCItBQ1V4kBBxw2jn15uV/yDIrgYtSH5mbnBwPDN6voL8v5AmKp5CxNhrj8JyQ5F
mfLmwyqq2TFqAY9sELmHe1MP4mOvMSITDe/GDWgkYvMqNuceWGBXEDpU0ur70jtw
PgOd8+dl8nIU1DJO8AEHkYt5a2FAOZVetdL558fUCobHYhNx4yiqKDGyM2gwYT2L
gIwSmlAhRvpmHz6V+ziiVKP6DAr0H+57wP56lh3+PGpMVHz2wq4iUCJavGQY8/R3
uPZeny/7YUXuOIZTG4NDcxIV3TpDBwsHVoY6+DQwTzKWgQucfcAu6SFYT7mI5Yb2
OKj7ZipKqNB9J/rzfLQrpHoDgoFhyrVbL5ciJeSI6YjuBdGIlH9vWRiRtxARcUX4
upAjt1vDTqTXyalas6ZqUAAelcgB4NkD59VFzLsEUobErEa7ZFBU7KUczEmlPkLA
wxlFH4VmB9eFk6E6sdM+R10VV0BivXZF3ysdCvaQtdDYBuCpUjrDN5D41MLUana3
X8wEzGCXuxoOX598iemXyHKdPzbP5HD56BeJuaY7s+WUJZ0pzx8XC+6cnS8GFroY
1jVZurmTgEJbZyHaNgD896Ekl7DOLLmn3CJrGwS6M0S4Yf0FuOA1LhvkJea07Scn
G1CnvoWt/EXQblykscFuzjmxa2aUvXsP7l2UMOi/f1l5qJVB+BnboJV94g1vdn5T
xIdH2b/x2NNVArE4kbEz1pNy4tEIXuAWo7SMM4WxwoDJTynBAgSALa1I6j3kjfPp
6DlrrXFLZiP2rVXQHcUYiM7DW2Bhkpx61T3Omv+mE8NJNW1pzml31Uti15DH0c76
SR4c9C7GB3Df35UBW8prEwc5kQxTaktrIRT3oTPQl1zuB4fCB/PS9qoV3pvJlqOb
1AQyB1F+DmuNVM9MeTs0/x3hZI5+/CSb5Bti//fGYfrztvtM5DB3ZC335l2hYear
eNxfxJA2wBcXf3g/EAHHGoYNV7msj0f79eIZWVS2ReX/6cDtRX9hO6JDnDz7qfy2
c0rhUHsHwmmTmFAIzBKmxfMu9Q78n5KQfA9PbuQGJKeNRtLoU4Kmb55caueM2BYv
lOiyKkHl4JT0xLzfasHpigjuSwCcIxHAGI+IG4plgJBaZw650TJ1gAgWRjERnTHv
SPuXG1y6uOW15Z4VbIceY4oIK4VSpD9sTgpAEDBj5iNVrxv+5UefXA8GNvzo0HDf
HDdHtwpf3fAkyJx2DOBO41Xsr4EbMFUrE5vtk46ePLouzBoNItBOY92Mu2lfCfMk
jrJ1SpzUEGqwJaEjB/4So/KZLIDE4CcjE1XCTedgqNYMnfDYUbYcoQLFP5VeKtUT
3AcV+KnaF/GOKe0yT7sgueftUD06Tb2zA9XrDU5DjTM68QneQkDqywjO4dFj8iB/
0G0BgVpTEXzuyrg1lwaoEG0CaU4vaFTRB3lYfLrMoRXCoFLCvInxkbZ6BIYFmFAy
VhzKwC29E+v9UmRQpCpMmF1L737OM6hJHemX3ta0buBA8KzCK6TGVireRcyI+H2+
b/hezH79eqHElRe2Xj1afSkwwKr7f51LohcWJiUq18r+RP1vMCTbJyDWw9ab99k6
I/HPThfishOqSXKk8cxIbOzsJycNN2JsvJmE0FB/3MkG6k9B+qPocZkNVZ9ARG9M
knb6++XJZrhWF0Fx6iU1Vx6X7x3Z7TsI0UA2mR4R4KgeFrFB0v0DUSy92sn+TpcO
sCA3gpQeroYhutfgcGd+8chwfYO0Psus2zsVA76ExWAVpxwKOOFm66VAfIP7nF44
xSe0/TEm9Cj5hqp8PjzDNrRcPrRbiJsFwnSkisWtWu4fru/1A79emK+59v5VePmn
iqRnf7qFkCGoC5a8TXYnLdQbCIHbeS9WRsTE2mxdsMxK+Dcaod+Hm9E9MfugkpAh
OJjJZu6AHmcaa20ExRFh4b4kKUjGaMSrd+UkGfYFuC7wUyPNsUbQuSUo+dRBBQ9Q
LXHluKuW62HxSbaprlfgIXTXBuCnnUU8eVYtF28jzDx84/b55eOqyGW3sdkVsuZR
zPNfR+IS17ufURDzx/FmnkJdGyttPWVLEFFEt17mgM2TDFpAi5v4rY9vuKc7o0pr
VnFgElDujfJ2/qx0LIZd+onuuUHASenKatetNlN7HaIvulIIPopSYQfwDm7Lb+cq
QsYzhHV4LskWslHEIpsT3Q06Pyn56ApJqVK2TK5F92BacIP7OGJ4NntGiqlXhF2A
xis+cO/rS++sx3n27yw8gbG5NMWqySivlwiPAvXpu5xiElqm6e2SPO/xrWHS/xsf
5Wch1Zh6lGFjyLxy0OKMCr5Yr5/pSz696O+CzJc7pClzL19I5OAkxsLNQS/M8Eo6
wMm1Sw1nbD3G80Ysn7JgpTrQgq2qvhjghUgRZ9EUgdeB5dm/CMDsQppt8lhwutyM
2BwHe3WrmgBBJIWOF5Q7MC2Ag1Rry5SGTnXJta3IOs9LekuVW8BIVd8ysIObiXyh
pyNyc6fvHZZU6LqdwBEmiQ/ajJY2fqkTpNNpMna5ehuXbe4SMF/hcIaJFlY1vC4I
rXiiX7we7nXJQAcQ8+PvlaE2DkpnPsEf64GfvibxXipt2RMA8e+WSDaGmKIFZ3yM
drH4uOihWhnhUqGhsNi/adqqF9w85TVduNqW6iMhY5jiyQtCFLWRNgH6qAJEYtrb
zdWz8dt9dvzse0lC7t2NiwvA02otGnU+gUa5VvBtLgpBO9N8irhQcUoLcjgVDZAr
d+wDsSqLGQykuHup6GhuC/2hudit1JtNA/Fd+ZV4/cDCroGcxgIf3cXD6xv6uQ75
KqYby2czsJPIXGnfr7SqhRgSUOborHqEsEsb4iSwP5WfWp7eGVv0CgBH3QEZKA0a
heUlniJ+nUmDN0GTzsBQgJNFrt176yCmMoyHTxcwD7UNUXu7/SdfJF4rKUwGusap
YHgf7O+EVy/w0jqrawDej10/vcW2MQZ/tjBVA9yG31twkqzAJ4tYkglzja3IEb7+
WDcwYVY5Up+8J/M1mhABGx2LzE9f147G6D/j6Y61fwJM5g7VwRE8ZOsStmWF9q+F
bZs1grAmhOi1HFO5Yn+d6CTETAUV1ZmysgXYkWEnu+X5Zx0eU71ATNoPi/0gOeXT
pBb5+6NzdmQvvX197sLm6D+1BdNfMpRdDWCyIUAPxIVzzZtpcr5ba0GOKaKKQngm
4sFifYdOH3LDjRr0kFzUK2sOx2ipvVLsG1BN9sGPmWGw4i1L+UfakO3dUluyhzNC
4yfMY+Wycis8FRfVQHQuyTIPET3AJoXE+jsoTD+GVHtZXJKrEvr2wOg5OeZPhFoh
G1i/EX7z6zS3OKsSJ16muYVGRjLSIzPSK835/JGwDF/pLAwd0ltgyFHd6IeMCXjN
3b+Q0vgFnHG+dcr4KTA9GkmSJ0yk9BvdP5USf64rdYftKRXTp+kjSMXMEZvyzPRE
pFCmOW7zE7fWriVN65KB3iyFzbA6qk04/LwIWverO2K4s1bY2+u0+0qI9x4U8fEM
2oLXdKzs30ZJEkhWHmlIakBfD6f4XM0eRKfMML2QnrLFv1FI7AidcmSpxzwmZNcY
eb7SbiMzUO6/1FNoaF0iPvqLC+G7dfqj4wa4towhZSxwsrP3ouTvJhAgXwCHNHjI
XtzTrLHrIqTNM7pX+QikMwqNzDs132EJH7BqnqGDqRKuqk70LtIOCqoxCkqQEz2M
WLAHtcgmJFy2UiLyMwm+qJJgpDvKZlisg4TC0Qa/+sxwmYJ0IiQLL5Rs/s9pAYgI
P16zU6ekBev0KUZmD6bfy/FMF9GHsibd7UNZJtru0F1qYDvDXpiiXw2nahovelSo
X6mhVT+TVKpQskabJKPnYOdH9USgp2WmIvSeoIwupqSehuL7/Wv+Pch8pDcmt2gr
j5bIXlk4/UmXQHWMnyzAdGovAIbWVGYTjhrriKrnkIsCP2fNzXhSQR7rVR+v2k+W
RjbYdol5ZhB4pw8ef/Yz8GK+72s8c7eqcH6rgqf3uITiTIQlDIDxsBx5nGojw1Fj
HoWggzobDccVNZaq+8StIvzhWj8S0jCrjtFjXOr/3PRFqw8PXmRN+RNgQVKXJ3rD
AacOJfLy4U0lipjpjwJXYwisa+xis/48HpilLuNbNiFhTyV8juZIlgZxVHfW4rJ5
uSOk3pzkoiEyKxcAdAFT8g+hZqj3M8NHKlxtUgY1vNEL1DJ/V+5puaPQLhZI/8Ri
fr8t+aS7X7w0JrdJGQ3MkAV3bi8+SSy0AwetJxLoSdRjj8CXHz6ZhvcIdk++vlW7
+NYtKPKzT4rj9nj3cjSqVSw3xrZ9gcVGAM+lCr6fLdeyphRy01IY1lY4ehSW2bJn
ZG2QVrqTsMQxnXX8w9/MQu/5s/PntgrhcVCg2fKJrhWHtsmqDiFogicbs0WAtbHn
ACxV2Xl0DRbfLY9MQ2Y8gWqiKDvwF7XENqQpM1duEAQ/aCSQZPPOOvbZ4t9HUUBV
5m1spmRSCtQXa1ZiA+lJmyhU3nfnltqd0N25PxT5j3MuP85EjSPpR2qBIbQyQWkl
aWn+NVZcNytUsze/rv9dpYiH0tMqfW2gBwBa85T+j2dl5O+LixjeTkGGwlyNgZdX
o+TC6qY/Bo5BXA2PJ+JudwBERuZKCPOzruUvse0NtXEMEzRJHCj9TcnfpmygOdhC
FGWGbs5d6bQ+BxDcW9ElYb3UUombAjeqXvl7TDU9vnb1e1E0Je4d8bzxL0JoTibQ
r/7OCI++wv8+kLlAi4Rfr8h01Qu55v8sGPLiWyUDFxByvw9UpJgICQFzxyw+Q4No
TPRT+53RYCf9vVca4ewqoW7F76wpngFDhtnyp9rkhEY2ejtVYWA1UXUcjBDPANdx
MNYEovmuJi+FvbbwnAcnpY6rmgFdsfBJ9in+8B1Rl0/5S9qG4WFWoiGGIjwuqneU
kn+yZRd3f/RQYFXq0qq9aKPr3PssWYp4ZXZu/ceZ8Po1h9NojNyict4TL7QYuSVW
sEW2HV7XIu57L41xFHWL8/bnSOOu6FE2ckteTcAPZZDFKx8e08BXnZ5P/fbIGPjF
cHJuGmG9mqpxQ2zlqIcePtZlXpnM9L9WzHY39r3n5v/sjrBIDb5/BCzUMz39moQI
9VkPDA+sC9Xow2T4x0PoU3VRt89gPMEJNwL1HtK3E3hv8QKwSKPEo7xh7XxY3AmU
9HXK/rzXyyCTyl9QnkDn8/YR8XkBCVT9YiRJqeG89dHwzIwVoszctUZx/dGBDt0i
CknI5CFNlciEIYh/VWqIET9xmyQLPhkT+KSsgAznpJWSeT2Gw0P3IVjOwgNG2yzT
GE2nUZTiJPmXcvOPiWiqymnAu6V1YEQaTCWkxy62GHvc999DflEHIYI1jCinD+sK
20uWC2xztWFYeOS7tBL8eqMM71nOWzkUCDN0Mx880FCvE/lfgGp7VY9IduBXcaZT
fHGPVTBPzHrz6D5ZLLRrFXbxNma6fKm4PVJrUuDSwO61XdcdHYz4zNc8g41JzQPg
1xJQ/rhy9Ej0+hanbBdZOJvLdXPDwTs/A0C5RXtnihT801maDcgBh85noH3yKUBk
LwOnylOEvB5CiwcttGZ8SU8QGg4j4X5s99+0MzdZMwLN/gwL0isLzLzOsZj81oX+
7zVXp1uWRZ+YZLngq6uMeJ9VdrPaqAB4yUGPg2V5Ipe0g2HC3PogzfqI+5/+5k5x
AbzwOFXSYrBNI/NmkWHsz2Hv8cnPG1rYqkeWuoUkBWPo9Pb28mesajdkVvJ/i/j3
CZFo8LZcPJ+S2/fJMe6yLvxBnH+os5F/xhhAd3s0YG+XyBdCNWujKadQYbFGMx78
eFgScnd3iXw9mnVwlqTPK/+f6X3vqD7HIwwMTFPj1S7rr/4LncYl70BmVzd3BDYL
IC5yjoq3QseJTX6eK0kckSH2B/hQ7OMpCKotf8rtoyYgWXNs0ORiqHlKxVxYwrAk
Gu3K0wBEcxCjqV2003/RDyqvm0HhEBJbBY0gsthTuJOn3/WoQ7IpDNJ7MbRkajQt
O6vQpPcXxpcdioC57nMYuJmCLxfZowPz3SuJaq0Kx7nK8iX76BPGcoBGoHcAt/fE
fD02syvoTuwQDJ6wYLP0X/+Hl47z3rR93N8Z68g4lb5dTBoINbfp1fsMh2jcKBM1
0IziQRfCmpJHX21N/mCeVhNwa+6QV8Wedg+/Ry/zRY2110XrHy/EjC7eTP5V02zs
O6SnhVmpZBOsPpcKLHNn9P6D7KXemOLGxLIolqi2gtjmR3vNKqgwkn1zssLecYx6
IvTvHTBfQ4INLJQ8N8C0FD9SyySEvqXKqb/wtLz/QERq6hnrbdV8cSzjGnZfhI9z
5LMTl8eujmA30rG0kjqYxusnQvAbkQjs3pi1O4NeKxCypoxVQHWnmPZX6egPTJL5
GmWLoO/JkNNQ+VbpBaecOwPB1vyYdHLCFM0AsW6cb6+BHX9XYOSQw7vYIEZm3BDb
rd217Cm+CFWlNTt5AjkpKcjZFbnQjpMniQJDBOa5mO/bV7o+bqnfBKk22MUZbBjv
ZnIMq4o9QJ+BWvW6SqRM5upBCD9LKa1DQuToujseXvVvvYlDtq0sROrYN8YqTQZl
d2U3k9ROa4JtJt5EO99oq4WxYDO/1L5U/A2zeLb76zpUOeUtxXYFSA7jJ7bdT7pr
P567Zo2sJhbi2mtK2fejLNxuoJ3Z4r/hC0keW/rZawjBPkZpbA2C/vFzGxgGWKIZ
zFSyQNqcbRbTN0PsgJ5KFNGBIprQSQm41DYVADjs7w5mS0Zsfbxw3+8zgycmdwou
XqjeREwzsj4WW6fhg4JUeKPmZgOSmbJ8GPKb3A3heR5EHoDKFlgukGOxh9tO4ETv
kAYldZ9JBs7uvT5IraoeeOvUPAZ3VbiBkzvbcfjEpMMfoUOXsLR5lAzeNeh0sTEy
YD3cKMnrZDfQmpMYzwL/6pmajRLCA9n4eXUCsowKPg5Linp4dGfip0JJNhzAuirx
a2sFHx4Zgi1QcWgvdTa7IaybQmLd3YhCqJTLjYTgDioLVq8Oyvno+Z0sPGRa6R8w
HW14ugl9kv/oFJ7NLrEC9mHxT2LNQegj1WPz0eICa4ifjz8ERnixfaSEYTI4PrBx
iL4fvElSyywo/oITOsRid7+vbw0xwjKH2btvotTbUGYmvmgukVc8v8DXM/iRPHIU
3o0/g8hNHZUVhRl8cTExcCWt02SDf9xAXAJrC4hgtMifkywETCG6r/CGDswh7Iwv
3I9/T/DNZVRAjM+lKTE6BW1Spb/Gix+xQqPVVdZQEZGLjqjVtu0U1+jnG5RP0527
otEj67HdEj2KpJKNzdBvC2OXe87tCIUkqcuQA7k4tko+bqOnopJnabwKAA4+rNUp
nuY5b214j1mLjX01+aKB61/jsdOx0zX63SGmoPI+7YTn+ezmbrx8paYQKO7vrWy0
iRFPo5QUhE+Pgj0SclnKVuCbHzmb8RTQKXzF6jKTKUKQ9aQJqLnjG2EeYdCl6j+V
JtIXAA8xiDA7RuhPzHAxw9S4Z9NAk/fWiuH2OOhxom9UlbRkr9MnSmwce/s1AMLO
FJmXCg/Lkn8GvOQoOhSlwKZM6H4jEbgTE3Rd8s/tddOmPK6/iGLHm8m/VOEVJG8h
vWJxjQZ5w/C4KenDMcjOHT6DgwcilvMSq7IBhWYxUwONjTwjIbHMXh9oEW6r5ycI
5Lh2qjXxvrsdbPdHYbb7dQugn+VwZHcEGNH/LaOcxB0X65hzHRILys1Vv0AMFgi3
o8+e75XT39dxmyaP1VexYpyTSirCHZ7cPeFeBk9HQxEPjKwvKBDA+3Xo9BcmWfQw
yvXhKHRfBwUNJvqQiAGLFmzqkeG5XS8VgiFBx8P7qtan9a6m9RrCrxNHjrNo4FnM
uNjLy0JqU/ED0C3HfgfN5mPA+g2sCiw2CFnEPF9wI3TvUCcTjwq3WCsaqh6H/W1s
N41UQLwtdvUS/jSxunCmLJykCvmqCkYyRZqafNYV/KeJhu6uw+3V9hDg+4ZXNLc5
KBto/NgMfeusjkBptgnlCV46nHlLLJKVpLraTVFyGaflokykHq90jvUBMBkFhJ+I
YIiTHMZPhDm11dS0A45O8lG+SoX5m71vRDLjzY4o/asTmE7gc619qBIXYkFsHEWi
bqHKjk0W5MIqDodclwGFt3x+yqLe2wFUA9w7XXCRtOAs9krCUmAlcBc98trTEIp0
/poG4j+FeU6JUpjdCY0mxlcpL53YNrdoPrEVVNUSkjjcrK1u8jXg3QTNFWejQgnS
ulcQ8EPnMh8NCXv+Ps3DW0K0yGYmYUIecN+YuVh8t14Av8F0QDZTrxB9FdOeHl2U
1xvHYAVBuX39FuCtByqdEBp9+0E0m8goSodFSwNrKn0VmJlczqHnAk3aaWYJe0Eo
vVwp6EtFz7ab6twJhTYOQHvSHrGspuxq8Ho1BHwBWjgUXlLGiuO/5XnT7ThfjiMF
I6WovBe2YN5rEZTFId4e9GH0RhX8QgAQOuNboqnKK5FruwXRR3mTFQAxGOWV/4b5
DfyBZitRNb7ptzOpc3B04LFqFL2PtuwGztP5Uv55GHVKVYVYRkkPueJw7yU6nY7C
15O0zlABQX8qVhhFNwRJy78R1Yq5UppqZLYNz9UaL8zv/UpvQMBnGtue9z9vWEio
vsN1Og/JQ1LruZhsQTbGerZgpi7TxrH2o+79L83rSAYcq5PtRuX89D7MOGh8F9dm
GdUOBQPYiCluHKuVAfx7MzS7XHngfMSy7ysSoZN+Ba3DrFSFyNYE4k/62E1e6AkO
JwupmjPXCgSCkrTHkniA6iW/15hwgD0B3xAuTwx1HrD1G0Sji/IB9pvZ6dIErgf2
E1xXfgYuWXeOTavUyMq7KkbI7/JVCmZhbU/O4Y2CEE7imtiF2NNOGU/QQk7z5hW/
mukLkzAA80r+hMOOIloD+Dnzd9Fn5JXBSp4Tkbi+AOe85urTbwg6NPDZDd8ecgOa
iG1Ab3zI+yc26cXCdykMlJPRBx/IuM7i2XstaYErJFjjxBE0U7m95Efa1mtdl1lg
VpO1xIEvAHqzTySbqOxZcHccZNXD8sHdauKeDG4cio+KvZd+NYhmTdJPUNrzOE2G
vnQZYqxJN0y4FODxWa1KSKenw0lQ5jxrnkfLim18hnsK8GuTdwwxKnBYmzonHePM
lpxTth0GQYjrEoem+nw0J0DChek2ERMQnSEods3IQZV7E2McbF5tGsIApg6wLWQX
XvuZyCE932HeM4jsrI73ry/CJOQhI7apUOWY9lep0ZRldsIkr+rzpGFudK3oVZ/t
tay+cSDz3P+jQLIdY9G9l6vQQ22cs3RmbmPeAAypOA1a8FZgh58UqgqxIQMuEjZj
oN2NqOSKYemM814g2vMMVWQmI4hC1Ky5WkRuRlL72fqpGPWPTi+QYr17JzSaazAd
raobb3zfFGA9SdL1H7a/CkQC0Ac6KDrLGungFKoGmgW2TLn+g8+uweMoS3Suqdxr
2deg/Lu81tNEq3/8X9eqrppvmgji/6Luq1U+DdQ5K05/qO0wElfz9lyeNCFGC6Jg
dQghGwcuS/Cn+csIaeo7XmZ5VH1YbULfytRX/Mg2337YCEG+0KC2D+BvOzaYx8J5
IzaxyZDZ+dKPpciaTg+94LMDX815XecTsQM1myx2gy5fnPW7OPh5OwkNajEVHvIg
BZS8F/fdlGPSa6pzdnjvvpMMyLhvcdwaJt3asmDpZiMDzydnCISjzE4fNck313k0
ZlmTeJRs/g/2e6wTmFSZ/doCPcxFzC0Z4OAKs3+xko+MNjPdLucC9fCxATQLpdAF
CtTcwH9l0DFn+OAVI9R9cUT2X+/buaC7QQ5+yPFPjaEXaGa1vIcIbdor0HHlmn1R
29IUalkdSFXnpAEJn7jstzk5oy/Xr9MLqwC5sdtDd2Cwf0+8eXD/FfD7rZY0aKl+
qaHVK7HD/ZvedvUFMXVc8HZDMZVwnomjCX+SO8UTD+oPwAhFp3K4bZVRgvxpryKe
UYTkWynEgL9Sd/o+X44vi7zrFs/kX4eyMZvjKuvNvgOn0EgCxlDbxoPww9bx5jPu
C9XDf7C5NLrxfkUHucMMyK7qEzwYVEMi6K7GteKAEBQPAhQEUzolUUfIdKNm55vN
ur/WJFfTCf8W5meSViEiSvRrxTMblgt+9Ahavv/6BcQWAYsPFHGP6k6VIboZ451r
uPeUMQIDcdfJyaWThlQZacV4Q/sZrdNvtFnH3XOxxPL/eWzw1n3KqGeERHkUpBHs
0MclfknwNUZqTOtH7rCN3xGOTflt+qG9/uVLoCPTAKi4k//AXKB01G9uP69KugX9
YgytfliMMAeeaDG+qR1yh3M4gw3pqa4oxNj8Oa/QGK+frkSfXS7tr4WfNrtPLUTI
cmWWlIaeDeaZM9p52/5nOH8bAtvByJ7Urs8b0kHPUK4e7+gZC4uNWNnIOurJnZBy
UhH8XNFeHCvAq4Wg7W8XnMN+IIc7Fw/+wjFV3WeRRNKYtBxyQhmQJ70huFw9ZmKs
JTJaQqLGO7yy09FbHuTJRpx/RhwJ+vOSkzD4m8EkOrGs62YPe1cZPTbae2s79/Ek
cVrHHqPbZY6sbO9S4vTBkpqcj99Ha0gH1qcbVNMCgA3uwhLKjkbRpgVZfS07JBAr
NbTlaL7wqBvymNDbU6fvhWnQmCGXRABxwm6zLD6OzTMaFpVC5ngCHEdww44GwNcZ
qnrgJcWsCYdjp29dlxBg2GnhPM4lVwSWLPHfng0PUWoiNX3Ai09cS98R2LhoRXyw
HjXiI8WEoSeQs0WXwTD4piu4eVC0EqPWdOh0k/d7T3pWDZSKmPofXkRNPbdiajJq
r/1ygwB12b6BJXYcCVTlgJbAODZB4cfYchnGiLPZZNpqtuYa6k0j8Elm9Hc++LVP
WLJmIrtNSnFMvToch6vYwwwPQIgcfiByISgSKeX3qNptfECJxTbyDYJp/N+6EwpS
vqgQ7Eo2rmoW6pNeYH3ecK1XXnECbwu2nQodri5kHMP+XV6EoXJvoAVwuigorVVw
DhvC/VZV4IZMmUWuEHmkY0RPtDO4+7P6MtrSFYFujVShnRy6Q3osjWBc83UzvkhO
6OcHXiAaTmqpZK7t/SwyPEr17XJyCea2WM3AJeea9Fz35cOQ4Evr5ZTnRxj2m6Cl
y4Kk/HkHdFcn16mupYhnb7YGrlDhV/iWb4OUA8r94URU2DAY58wRwB0M6oHuD2ff
9WrI/jrMlbh3WxWfWaWRkBhRAXmtIz39LUQf+Ft64JumHIX8I4LkZ0nDBbcUl4dG
00/VCZc9Gx+tYsM6Zcqt02TTSJicG0+A5fBUFdQCdL1cvcEm7gETD7Qccjfbh5T0
0AuENY2oOEu8PAPKa5dc9AfAaWywrQdoYsRPRahHLjr2FLbQEGJzJsOwW39M3QVj
ncBEKH4o9XN43mEDEkY9r/tHRt6DYqmyp7YckUOCtjSdVTeAwON9qR4GiZWpfzPq
iBr3Bbl4hOgBsJEcLSA3BsW4eYYo40ZsWBujQHKxs+DXHy3DdSXO1QSwqX5nY6KB
bxq9e7xA/RktKk7vTOKz3srWLczZtxrKW5Fw8T+mqhzDBSHiad6ECFzAoG57pWMd
IMJq3JICitpkf+mVY6EigOxg72122Z4WtWv/dLxCQyNN3Qheq6oNwUxu1I3YX875
i7cAjxplkh1t3049Hahox9nfRcyP7c+gw+37w9EKA6Mo4S/Gt761ORselGJMH7U1
Amg9sM3kXKqYxhdP2mqcW7jNMhwkR2FLRD4VzIRg3eFxDXt2kqJWMMH5ghsT+SyB
KM0uVw5mapSEFPVdr/VkWB5O2hHPVaN5RFEF0B4KVlnk+caG6u/njH/RjSyATqU9
iUP2l2WejOvIzbBFdXv+npUokuUhKYBNmrSOG4cGhyU3JyBzu3/JA6WMOcPa14Cp
athMaLbY33Qce9pWSgjxRqkCtSjMrF8bkX2KHKI0lr/OakcD/ZvSrO1RE3BeycPG
AGhBt2uK+brIZ6dTicAbNzi8why2Fs5hCyh3awaIW2Ba66nJXejRnojVIIiMIz4j
04VZ2KivwajoazgQX0yVhr/T2DSiPQmfg1HYC1VDg98hyRE6QfI26+lba9TRK9aS
OPNKHFDGIVUA98nxNXEZ3o1yAcP3hqBLa1J8Gg7QBE/eqkhSTZl5sw2WJIMdzGkq
9tDBXJIDS76EcTNV15Av3+PlO1xlJmnCg5XTFqlqtV1Sx5hsMR0tcihCuyazu+RP
rpWrNcaRL7CAGPBJNpHDdoHnC+818t1sLY2JWasH7imdg3QKhXjL0X+XqE7j+/Fd
JqHy7BC7Zh6Gur5Py/tHJy+iwNq5aGsIrXm5BcbJk/AdQJNORsdKvOqZL9HtuAHJ
nurS3oXXcZmWTYQQefZvqGTHBU2SDU70Rfm9GYdR1iYtjXR0gMy/pL8Hjh8XJDeX
T/X6/fxTSTkKqHeNKube0iMcJKQkRQqdTORMBLfimhGP+LsyaodN3m2gX2M2vp2T
H3cAqC3AmYS0/6HYBaFy1qNPwBD1sdngsPrQkFzcfKvIZDaiRcEIQYybjcade7Ib
I8isVBv9t0om8pLkPmICLYDamuHefOSN1ontDeH3R5HBdfHk6h/NfXRNPe7hNYaC
M2q/B5bc/PS1rynMG8UYg6nUQ/nljX1xH5110q2xkdbmO262I7v8mgnEw4MECFBX
x1e/NjqQT0MnNQEUJz+HdpJhcygAbI6bl5477ahd5c0z2FVnG7hrWV0414fbvBu8
pbim905iB3T+1ckJHIoZkz0+qmcHy1g5u4mnGBpbh+HSpcX+cD9rLiDkRxS5SEs6
q8phnzBV2GnquLkqB56oK2C0dhfMPaQhfjUUgoROjo7UrfUyMtLiTkwtx5Ro8Igk
oURptCU2wIsPJlJ3YlteqHvlvyl9EprAeDTvyCFuvG3vGbwj2mHs3SV9aee8CI47
hzTqZVqUuC8mBWekvDHaYSJnHm85N+BhLOvuQt0QVLuhqxCw/xqMIzZi9TnpOQ2v
dFbqBtrqZ9eLEJBxYUfb/1kz1n8cDatjCvMLNb+iN1zGDLciZm+2DjL9ktlXJ+vB
YNK2dePn8/z4jZ7RCjLD105CPG05SuL+A4ZWr5vKRkN3LKGlMFCm7wJPRXkFUSg/
veIFkDZuhWzR4m/ly6fwHqROLKEjYWDABrmwThwbvkc1OFDRe6aOoO03TrcNzxjJ
FuVlv76BqBLTODWanaXNA2QPlUvy2tCzbbZIE4zM88T/fa+ghpRD2FPumNxZRqtO
2iKUnQallc1cVbec+adLBdyJ66wQI5uLQdMmTBk969ROYJA/Iavsr03nN+CF0kKL
2JTpLDgQwpuG7Qd6IIaHJ4y8y792UNJx5cbRkxfZngwYW5bwuL/jzmQBuGUYjl8e
PbcqfNUVCOc+58ZjfysEtrVhoNdXgGl8sV01dRBB8etTeI1AjKKvgeNq4SAeVILd
Cwb40vz3S/LVDE//3pzn3F43D6SRovgQddeljLdmIozXJActvRGIx5vHzkB9sqUc
jJFFChFqtYkNuZlE5NSjZsJ+0hxNPM6V0HElsdJenvFhduRAtl9Qrb5qRnfQfAoH
+KkRb3ZqyJxRhxaLRcYfq3QOD4lkg0XTTO7QpKNiEeagqcVX3N35kvMjDh17gyYO
pU1r36YYU+9Nxqm5tq0gZCzOppX+OJS7WtWJPOfJyPcSaRxnGc+mrwAOEVMs+Ve+
tgmx+n2bgtLG401jtVAx8sLE0I6NzWEhr5ThmFn/v8+FGRkQsUJXwqNPWrhcgVSF
MuobvH3VtElOmqVZyl/zuoj4mZk2Fh/a7hOMQA1fs9YIPDCJcVcyXdP1WHr/2rx+
w6zEZjQRonZUmsmrtq2G3OFk8RFc6nQkCf7Ae9RgI8kIpHZmgHJU8K55o8mVcoTN
gbB1QZcA2KYTDDbR+StSU1LoonNmAJuE/Wnv0E5/CTLgfGlbewHKwHk4Tl/fakJm
lt64CzBm4U3cGRI49u+D4ryJnpBRhe9c6jcfJCZdN5tbZh8RO92XGoF3BmrU/Fh4
k+lmLYM6EsCpVWzdMPfGpvUrmvAltDxfzq57B6wY41GW40HDRdD8mBCN60OOoqDo
D/uwFz6qUxsnssprFlQnisnmBpUmFwjyvSJ7fzMpStsmfNcEOuk1TgL8uMvudck3
Vz6e4OQCLK7Fj+OUYf/S2NI+JoOKg3T4OBIEnCuxAAabQjjYUJANQJSeOuQeyqBL
0GL4vax34DrtYGRHKTg5nlbVGstTw2dqkkDAC1Iz1tJNJ+n5elcPu7gYXiJWv9hP
yJeHrp35xJlUR0lh0808lH/XxqC3R0VhJk3h4izeEAP/gpONH7qEmXdj4qd2Uqqs
sXMWiOHA4nw2cX705bx5Ez0uu9c26JFlzRXTm0z1io8WafruDhszxiUqWtUMz484
NI08993RqUbz/g/sHCnDRvRn4H4/vjLo/NOuiXAzSGb/9IggTeEKHAXV+bwGz6RB
GLIGDRD2dXK48L/gYxIMIlfYS7HP4im8xN3dwbpojQPvKWfeHA6yFtM+mZmZJrh3
7dhsMIsl1+M0+Sa2WM6y2Z2lFy39LozPd12LOi/kI6dGvj2UNVIOqVQnnVkB8EgQ
xdHnuwPeS67Vsee3qMI23oN6X9xoOYmpLyhD7trablZpqWT3LLYuCVOv5pS4/a1m
3sxSW9mf3Fh2Jwph4O6vSOKsvsI5WqeM3zFt1N4k0RsCXP0gi94FpMX8Ru//nMgV
jSfOwvEytfy4N40Aq6kHpym72OdMlj/c1HjyYJIjLZaJd0ixhK/0YQWbmjfEGX+F
xPaowWalLi1UbcKf4sv4xhfwEgGETAEq84ryO4pJfpAKRVZn+qSCStyqakJuZuYg
leu/oZMXXWqLQpZN7PGsbRW7yOoAO24I+03GaktHAMbsKG8jZPojqHuJmFWheWfz
KorfpAvOLYLirbGMt6gSMSpcd96XXZOYSjTqcctYwJL9505kgRT9RedlsAlrPmJq
3JF00r+PDQa+u3LhRMcTFqmZbQaoH8MEQ49XJUiw5UFR/nRwOgNSeAfpZI2/xYqV
ncH8yJZGjprp1buRpX00J1Y6tvjEkEawLNVtZ59KZnYlVFsJs5sc6ERz7dwTxAqD
ARAC7e1A4mvSlIFJ1ePfytASqX+37HPpgNVT8xl1McfmI+9szOvBFO8VVacJ0lZY
UYHwJF2Cvi1fGYmxIZA2JEuh3IsIazaF52kSG67ZVI/Be1GZAhWhLv+iMRKmA+M9
VjLteOskVRK1Vkuam+hU8BnGk8QF+WtgjW6gEiNnr6XNQJhjQ4GAj9v/xZtimxfS
Eus0JJyvYFv1wCCq5RnYwdSdl216Et3lvdF5gbR7/jwA1z6ynRDawS7H68lTAg1i
Pw/ADffG6UbiiCr4gnmSJT/hr6mPh/xTLngjmXYGHzDiaFXEllsDuSl1CH944DcS
amBU89H8XoFq6DwxETADGzyr+3R5OhckkUHW20RE5lEOXBw43YLVqXqk+JfZPq2t
ZBWKLMySBtJjvLJpKTv1tHiqLu+8I23Q5oJHALjgqIzRS/tHXiNKSs/HQw4K1Aa/
XkVmFP13l+0feULwnzB4584Dr18KRPwt8DIrCEFuB+mSOsbptD1iLdeyUSahbePK
lQZa+E6AUOZAQu+kmNpo7DUPOb5wmf+T/W3tjRPaSXqFfSt7lzqCH/j1algFdv1f
wF6DGCvi/pTtcE6s4NqXsWWFvTB4iTDxEMViKhQgaKtoAXx6AvyYVGzLsdik04JJ
qyQAxHoFeUBFqtV2ct0vtpnWcNupL/mR1o/cIbQpxdsU+YvQtROo32wAVIJ/U2Rs
zWMcaMqtN30Z6i9vBRRe1FFmFhDEG+ATarSw1P3Stg548eu6pJ7GC2/aaNzvKueH
MnN9fBH15mUo2C6/vvyZwIrv8LAQb4t61j4SY9y/PUJc4AOAsRmYIJI7XwLW37ab
TucqHArLtQFJzwk3XFF1ZOjA6f2g01ZdCx9H3c8fUyzSdLuWra7QE4eEfJXYKP2J
hbIU20YInWcVqoUO8h9Se0IQ5CM7AAHSP/7byUAHrTuTsr7uGZ6ZHPfIjTpUdHvR
oBtq0NjEeIysfMgWyQWbeKoklc0Ivca8KR8u7aR5Wag28ZlTiEGUXQEt9NHJ53Vh
/JPYdzPPgVzYU3leA8M+e7lPdrBdehadI2aApbJSB2A4+G+A/E3Rwb8umq0MzUGs
iyDEiCFgyAFEnfhze14TVOF7B+xihwXIlHsmGRSKmy0cN2fVqm5if595qd8Jgu4S
FWGCk6Dm6zQ5FT9U+AV1yWOgn5dAS0ofUkkNza6pNqXHoAtRV93xbdfe5m9Rgx6t
Oc6NoCiHD3qad5K+2KYtRkIFh5NNPqCyWc6xRS+6QfmKe2cle44R2Ai1tTaDDJtC
26QHxtYMIdKkUAZyy8bebQ+yMbyuXAor/54O+hw7s/7F+02oLGLv0BB2RdZp530t
bub1x5hJH+4pEi2nJRcukuECC5deHxbMpCwGnEuD5y9tl0qjiop/Lf/vPnezJRYM
cCVU8YRTS7BPWAdR3RoQ/A47z7ioWKcfRi2a9ms3bs/2IDaM890J+B5zNFmCqKsu
nvrtYpGPXLvEyvMeaCgPzV2hxP+BVwW2yabVwulD2KF1jGsFSDHqPxqjynFkWADF
nn5iGku8RGZL4J/vaCcCBnrZ8kowSN5o0qQW4eQ/OSAZa5zt8JDsO8PH7Pms3WgL
E9D7OgL55ez0rPrZLZx/AHPTQrsYsZeHyu/b5/V30pum5EQubfw2qWItJxQRFKiC
MbyMhtNKs2LCFWCaeHOx2Vz86xwznWduSRzWLUjSzuip35Bk+57JIYuVyh7Hw4s1
GaCWCYehtZzZ+ILkHE4hDKXUOGRUnlR9KIxVJ/0r7xpH1Ei1+JJcJYcb9/3Cxsv+
G924Cj+5T599Bxlt9uO5VqaJV3plfF/vKAFYo0qzlpH7pMf0B8Oag4ziDl89o4Pg
SQ0Jy/I5lblX9N1Zo6PMOtHL7PtGueAXNSNtKzx4QTqW+bHwxPuEkbLiTNuJrBS6
NQONpwqpa8bpW6oDczEmS/f+ailBpRpjbyREDPa2O76/KgCtj+ksMSZ0uuVxdCbb
Eho+mfC/cojYZx4gizzQeWQeXDvUZtz7UwT/diwVbdrTUUVTmci7XF8H/C3lcuHA
jI6ZHslCK4BPj7YMsTqICZEvi4Xk7bNqVSMt7NciqNJMdCzm9ieY7oQGaMnyMXC8
Jqr9qt1cOYJZZBoxEnD/S0tj8c6rUttgwjaMaJ3aHwMETTCdcJrczFESyDJPC7PV
/LFEqgKijWGURQ1u8s1bOcnHP+hz7QnaKjD7QY+LGZ665rfSCHMf9Y4G7p/zYsCr
0Ce1RAbotBfJ5XCC6UYGCTXzI1Wn3AzmUH7iQg1vMjVMiWuMyZspQiKrC1JThIj/
Tb3Kc/NRIXBsYEbRQLrljNFSXtBFN0SA7pQ9Lum5homCa++DoqI+kDXZYx3gtvfJ
KozX3jUHzPCzyYZm/5/uX8pkOXvGOJm+1LYO1wfstAEJ2HgRDswPUKUxMZWeWElj
RRwLMGKkREiemJeal30LQsFs1sV5dCniGSU8fPEvypFTnc+/5z8stxIWpAIZ6V0K
hnPkCGkZTLmg2zv11zMEBhcgx3a0xJ6KsYCHc0P4GshiUzNMuXUpRA6PDXm5QXNm
Wvvxkx0YyoPtHviM21gPqhxRNu8Ev/KNviH8Z02RcKZH0j0/nu4/M2KkdI97aEQf
leTkJlYzgHy7YQLbL74/Q5i7yzh1prPSl6vws3il6eZB+UgzCX7+fGRf/adxLZgc
s3g3Uz21GBtXGkTbSxoBL+yBTlQqqq/dU+N8zA9KT+yNqVSYqd6/G+5wVg/iQiEh
u3A43DoQkZgWPciSlPlWVdwVlNYI4CKD740LTbLT9lzFpPyMplNK8gRFKGYoiCU6
Vkg8TutxnqRkfvKz5a8OqL2J4GlJbL+p9VIEZeRbQ4C9AkhuWjEcpJgYGKmt1lIn
rvIT1YMBfftWvJl3T131FZlhBZ4RNdK5PoviKhqAz/hTZK8ZAisFjOC5S4DddQOX
+XqWQ7mePd44srxSwMUzYGUB26h52ISlY3h0ACpPHI1i8LCsM4cqzH/2/XoIbCHV
CfjXcMsH/AAkNee7fopO1h1/0Jri6380uJZdirFSl80HTVVwicsHE4aYisd0R6mV
RV3Dhp8mB0h2xs5+0Xx1PoXclKWggsgxf0m5m6Zi7Fmreq1A1djn+2L2AgQqKkFp
SCGoBzTw8EVuYPPMGIms/fc2LRfJfJ9Mm2IBK9GNmwWaMpF9GtJD3CkcCXsEOUeH
bLRB8E8Jm0tKnYqu2Q5fugCiEgdOOTur9EVkwn1IMU8DyVcfg1JWMJH+3CP10cv2
EBGJHzxzd9/KTp68ombSuaydno6mpdqbZyW9bIZ7NsDSLBHdEvGkYq18Dkh6w018
s3ssICkYKC2FWw8qSpJiPSU6NN82EzHcp4Rt8FFir8uA2XldWATAM4N06xd5SuSP
q8WJfEjJiCkmcJIKs33oG0AKHKRlNTtFT5vdlxJQsBgYQYNY1cM8MuxaWQalOKEd
0UTYGDrqYfHSXeyKYbegtVvPpRlo+aUAo/OytSgJ2PQ7j+Qi0FFhBIwFRuONjib+
DFm5Pgtv8p3Wm2NviBbxBlDwkovXOg52Q8n8jLV1uG6mUNita0rIH92NkGc+5JF1
NNhiPiCJCWX/qZK42keZdpzDURdqSivatY6Cq22787Inco2p7G33nuvJosKTswaK
yJciWcs1cL4DD2I6z2LozOYeVFnI3wCzYBotoxdGpAlPVDCJysL7lwt/BD2GkXNz
/qwMRB4g8OInuzoMuXG4HNEb6E/keF3NY6de4mmBGGAx87zQqMh/oTPYmc30I05k
O2cy713pSSl1105Lxi6oEtFp/ZYFwYT+M2sjjG8ffIC15/GIG1L8z92fU9Qw+w66
QsOTmg9KJvZY2HdfGVCWV9ddR525eFfhEA2vCQPU2hz2uR+kcOQQtoFcEI5EePaW
24O1EHLLo/VWV1U6ws6nhR5q1J7FYumEUiezAN73f/XN5BEyV8QwKnyCneuvqtrm
3FAUd92JRqiIUZHi3VLEgoupEorp8NE0I2NgjuQR5yMDGCKYtIUbsAoJoA4qiwv6
wj5TgdFNd30cMFg6IJx2Nfy53XuzMGCCyTHKF1XWAq5CfEs9H0F8wMKV+foFmZRu
3Nh+jKaL/sqIBMc+4fFM9veq8d+JEE5Znjei90aB3TD+5rQa/9zb9er+PNk1FaRk
OGA3CwgWhXWphGre21ztTf8x8AbY1MhP2cL+WcPUrL9Q6kTFSiw3xL+SQ6AJrnOo
LF2DZZ07tWvYQQvhq4aZRqO2PbHxB1D6O9HgB9pldR8/66y04pxZ39SL3vWFPo6g
+aA2Gvn0mHAj59Hm1EQpccKIOY3P618ivJyG7SMBkwvS7NoLDaH+tITHDOJSM1FI
bMdKd6uXH0qfWAQRem+WQtIfY2H/Fwrsn4ubiOpZXxar5F5goQ4/D3lDCERP/dXV
gf2wrHeOjyX5y32fuWu5i2t1vUbRICiYZcfQz1aF+5YUOzuk7kd/z3of9Ok80Tf8
vUCvHWX7sv53XlM04tENn7IQZUhZFDqY1dROnmGQMIeNLQQyx/MCmw27VzDERNQ+
+6lsO+9/x5pNfW3pLzEDCgP0f9BikGqzwZf/MRvWPGISQ2vsqPALPazcHQdPEhkG
vC84dsRKnMUvi1pStPZbu3VE/1YmzmBaxFtcVCPPRPlcigGrpfU9ew7NAGCtG+5t
/ot2tyg+zrJ0WhS5++ksMB/ajf2ur40ymlUS8bvHZcWKsLLlq2kXs8+mfRXa9R01
X4rZsqc5oJ9EZmzaXbRYacd9CnbYwAyVE52TUlh2k6YInim9vRy0i+SRNNSXK0MC
wRJ31AjORhmwsX9BjtHxkvphAnV5gIoSDzgaRRpdHHCAKQstWQipm7OWQspD1AOX
l/ty1nOP6Drryxiq5pPFmJzeMOsgm/plAQsDeHFy651hQjY8WJBYT+GAFdSy5D8v
y/ZO1hNxgF8iqBrlx/dfjqMBBB5qOodJHMnTBIBI+znnNCqag1+iBxX47/n9z8VJ
akTy9rcX8iGlaMjrzljLf/QdQf/ipHE//AgMFjTtVXG+z6O3LNWHMrLqIfrD8VXJ
xevimkM47lmsoV6GZ56BdKz02+pT9+phfxGWzlFNvqHfhg8Vjkc4YJHLCmvhY7iL
YuB+s8ckMO1KHmWST/KVvDAdniFxSAYYIhK0VTGr0Oi5NKpR8VWx1Zv7V0QDexe+
qElT3fc2Okr2P7k0HW5/sRIO5N0OcHj10uSnyPB36ghFazmN1vuJXYa3HrsghDn+
XxVDwXZ+AA3mRxUfVi5fNr8lbPRtU1l2KfHy0z2gPBjr9qcZLkGJezlZC9UrTOgN
mHOME7owb/+FRgUhkAQhF1HvqHhP3fYibhY774hKjaGMJ2aJQROBNVvQplKhAOxv
UGzBdfpPD6uz3oz3gejHWtj50yjSF7GB+WHWj6+dthTmaev3+QmQF5SPwy2WOfF9
PBTtxtqLmQNcTv7GnCT8DaHUrx4ReBqrJyW2v9tm2oSu0YKT7gEPJbcC61hmBgfS
p66gOxOdgOzZCuv9D39M64oqbY+VrnEnSYQzfmTgyfCo9Ex+oaLajzrtShlVEO+I
TsvgS7zNWwf9pfTMd7nQak1BHAlNkyJG/Zpw/hhYG2peuJkZA7Tzv//vxab86yvP
DhnJ/qIGPTDYT5SI5E6o/L/36C1FuxJG2hbzqTd/4RRL4KbIJauGDd5BGyRiz23O
8tL2KxiGRl/LzSXh/IoC5h4O54ltuo2cSRYyJYjqzxFrOxVbnhOyYXNqMiU64mEC
hbIhDS9rxXmdByGQizBKaxqWkszn1w52nKmK38bxWsNIBl4au9jH/06b65mcjBR6
UW5N2cB6bl83fHpDzGdLOGpYijL+HCbl4Bk+ZbNOUMmjZa3vZlAkfiPOs+4qHLz/
i3GOZYRw1Mbws6T67NI4n9YchTC1ICTs9A8PxgVYB9K3wATCqcaFapiCg/yutwO2
+5rcBj0U3yjDp2THp1RgcIT0D4zvQxYMoaCpNLizQ4nUQ+X6M0DVbWAN5AzVfiA7
M2348DQnqwrPgIF0d1YGTKHB9BTn3+mVEECxjnLOCLhna6mbwQBRb7ZXS/90iWDC
mIpytnpNpeU120mOVBuObkYboXaTZ25VbsmqNR44LdqZ/lWT4fN0uavUTWTM71SU
2bvt28HhJiqbvG+hF2KFL4K1fabQR6KCkn6ZG+BknWvk7TbhO88YIEjalKmd5P/O
Lf3L2WZe1+hZQqAnCpP63by41IM6K/unNa2lvZsYdKmE985y85P6FEp66PVKZCPv
PCozwP1zTfQP1IZWdL6twxuEMJbEfT3vev3fcHk2VLp7DIytJ2Sv+7L7w/0WO+pH
ggbxmxH8MmOPcEmNRk2tFuetRWyzJTm5CbTnLihjA4kmSiPzBg5Pne3K59dYvDPq
i8W+GE5pXv39+2NqZsfsUinNeABTSxYl1dawFo85U+M9B1paFAZ+JS03r2lmk0wo
Q7HXKk4pw+aZ4hxY1GH8zakPBcf+jJ07O1g06gjGkT2Z994Cl9odbyyP/a51dkIs
vrUkx+WYgdjyLH1GuyEceWKkayOFZTS+zWRzhHdkkFOfS2HVG4IbMyYZbsWEfK7P
L1AX6+nQ1CodYazDyGhsF7gCaaOB8aZPeuSfwBW/hDGwE3o5p2kIzfXvvgTzTFBr
L93u/1MV4XhbYVQuUaX3g89UbfudYMswfV4YKg7TfMPaJtx1F4zdPY+PDjHLkUjl
RbfVRwOslA0mSVdTIix+CQpt8byptqN/XFL7HehcD5TOp7Ow5rQTYP86yIENIrM6
1UVkBxxROhNWzMrFGwS0ULsniOWJvCAd7SzJlSkTbzX27L4vADSMA5b/TbUn0ku9
cnsqwDP+TTCmIIlJkA9JEQRkbjYHlx9hWM4KIHVuw7dI+MYw0KuJI4OVDmgGXEFW
pmRCGWAtI2fmTJtVVilcEATqEqplfsAb64W4atvy8yyNcDut7q61jVjEeztCq7cR
x3eAk9BGeApiLlhPuvrMd1PEqgEUosZYMqpQNJgjulCIBWjZQWjrCRAXc7vvK/bg
12ECeKjgorPCvJp2PF9YOmmwtfmooLZxDXqDsKh60PgZsOVhZHxDTox7UsrXtf3W
TqJURCODH/jX3XSlgt7jQGpm1sphgZR2n6j+zM6TgXf9fiSvAj1d/siMAuSedjQL
Vy1njR1EcctqiSJSV0PyGchFMGPiUvp6fWGLOa8V3ZXHcS4EVB/Yo+mkOE3jSf12
Rj3ECnovrXrF0akojyPf3g+nuqNInxbZa9QFbq1LxzneYKKVH6CLec1gcqMou5NV
Pp4fs91FrL9B+hHgtesBCG5Ftek5kOBOyBj1sWiXbF6iqUFA0iLUoPWduP01INx6
2HH7R9RxCuNl28zqeFKwFEyP9SydROLzPvp4VB0/pA6kv7L42PA9n6d2D2nrzY5T
jeVMgXztWSSYeTuOmn33ahcOtIrADbOutaf75nwitO4Blh6DpOYqQ1uRsrwXibU+
ognqSM7+iA2OCfiBQkUPXtkbBj8gPsWK5uQCFtpHrNtMkyPE+XPc6B0QiL4+5Kau
5V92L+u2vYZGlDeWZfjWxSx4f7VhAPlqeJMg2k9Gg8zfYlppMlbewaecExqV0hy4
j4c1/mmh1Y+Hr9/5QTT7mvUFIyN0t8bhXi7EXzDh7mRNBdxtE25JnU+Fdu6JNcmH
bh4DNOSdiZNVDZktDrxSJy5yJzZLDkv1kkjHZbYkzxJhj34S1D0MTQkKQc/BcZsa
HssB9vejdnKXrv/Tg/ZoFzZo1yyCHJ+PZm+YCCf53+EMFascLO4lTQMZM59PeIsX
dyaGVpEd3swb7f+99vQo+nVLbBnQ2YJjRGR7pC3vlztm0vQlicKu2xMWzWz41/Gq
Wre4JZRbOM0+5GTkI402m0zu/joDNdHQ/JN9GsUArq97egOxX2mueWgIlE4NyZWc
Aiz5w45BQ37IDl42DnBklRu/9+kZgjCjhzda6NXHssbAwONoM8/+yKKYL1p166yX
bvQ4dMc8obEDXmUDMtjTuRzSekKCZhT6L1iDd5K9Nw0UqGAsI+NnrZn8ti0Bgi86
3v+0qMYRi88zxmeB9/0heJBGHoPNs0BzQFyGvK1N6qIFJImWATeoYvlbZ8gXVJqR
JsBsLpivX4o1cxHY8xLo9dU/hNOKFSZr3hElYfmqd+Incu7rEAJchbRT8yWy1b7U
fM0dDb2C6swRCOBy7uqiM50xk0g/PvKOOR3EeLm1gsI3Aapxvg9WWjHgpMdVJ+Sa
7LuD2rUhKDLTwcDeStSJU7Ux7CTieJ+Ak4XZdYAYoXoaK0BUl/2Iehbh+HN2YVao
t18c+/b/F156UYFPM4ZfE6RtgiTPlgqAXyYfVPnmP97aK47nmXaW9EXjmaX4dmlj
nCWaL4vVOoeTspv9wNR3SfHDSGidqCmHi7FUsl3sQjemz9+WYlKWtgRmdsvKEUXG
o8jWf9lh2pxn9PEE/zmYJSspwfqFA3vOOB3ju2L9Q0HyODzdPLQUJwdZxmTP3fPh
Xxu1sGQZS3IFQrZLMiF+5A+kuZ7StxHxBYo41SGWRQqYYxgUHTCjLSlvYSRwB6k8
Cwn2MR4R5RSUJPm2YXuzDrK2O1b68nGOra55UdOHmonoOg+SUTNVX6IS6pSglGeg
5j+F7lwR/oBiyOtpdO2Dh51UGGoWoGhfQU4XQ3CdNIqW6HT5bXb+md2blGswxd4k
oiFXvI/LVe6cRkKm7y+SH1Fy7tUFtu1LK5skpq9k0TjqKN5Enf6XT6gjfjvAgJnF
6hn7LUHwHIFg7Q+wTCRxSgrEt4AddedQn0ItRA14SzD/fOZqec1VEmeIU/1POCI7
R/LqMR/w+Sc7qETP4kyIjluf9Gb0eR0RuXxZP/MvHws825V833SUSbaJx7LWCFAO
LTn40MLoeiYD2h16RiI1r5Pcg+0iEiJFcVEH3vjz+o0BylVzvGtM+QjuxzsZT+kk
4FeJw/VWoGg88032NVsWHWuslFWpKJKMm0KEVqovjX7QxZSMx+ekRf3b4Sn2g0Nd
RO+VzLAna33hOTjri+dqpaIzEF1FW3wZxxAJ3sZqA/1fbUvvSJXp822oGnijRp5p
C8lm0bmhYsT4r74yoUyrgiBBaMEt/49bvamkTYbm5xopXHaXMc0BF4JdZAN+/LG2
mxG8OIEbBPnAcNvIRh3Nb44REiZErZi48bY1VUpuIWyhZCcO6DLSdeHluiW5sHLU
on4q8EgKJllNK6ldIDGsUklqBkMHsep3unsVzzjlGjM+CsiIHwQ/Qafzx0KIFQab
816WqkB3Z/kot0amsr4JcoGL/f65LrpAq2ibARLIpiRm83uMVC3XcLAbu/pnPoDB
fqM1lYXEhwxeIWgkXj4nBi2hnKIlq4GhySGepoTkV8wkJ0Z468DbOX1UdQnHhEj4
P3Xa2W5OqDs35093Ug3X56y+nH5/BfcrpnavxUOVWIYTv6yKtVyHDaW534rqSICY
uTB7XKpUSABEzL3jb1S67kVTwylX/rnw4Orh4eNNEMcyUGTerGAM0GYoAznBjHnw
+/cb02jPnp+15JQypzMlqSv+VJjrvOAPYWWdTL11US2uqgUufrXIbu/VKCFS9hwr
9MMwYct4zg4vJZLEWrYNXhRKsNI95QuvDpsZ5vBrkMhOR+2Gq/KefLJIQ23pW0CS
BXSbRdV2Fw2m07cxU9pQPdez8NiCCaRtC+Xs5TZsp3x+ag8shzsWdmMviDqgaOlM
ehFWDvdFOQeP9AFjOh/bOS1C8/v89siFq0emX2UneNOhiEIvJWw6GAO6Ol4XaVcx
dpqG/6+GqukuqkVccbpBU5RcQhEHR9VA6SCbb+HOvg/98sr98XznAJ/6yBTA74rt
gcLEs8vmY5qUkw0FDG7JRLVbNDPrsE2gdlapfvoNUXh6G/pBA7LNveHxnriJBCmn
lVDWP9r+tirxtBxsCEsnr+tiLXC6DGb9pNO1AZlHJLHXSPhDIbHI99nzN6r7j81p
81034IpNzD7xfI5s+gkrftiM7lzV6mhhr+lihFOIC9G5wohkJgMq3AMdhuBNeFFx
TFspOVNjqBQV6M7WUKRKohN40qH/jWKjOcenuOGBxVYG9JS7MZ+R9de2VQ5YlhqV
wd6a/p9bG9j8bznVSCOpPllifZdjr47r9HT/Ls6mdjnHtZVpItDUIrQMZy1/plTA
Zn9k7ehLP/6JBkU71aq5H+Oq5bCfyht7XNBc2unA/hCgsxI7fJCbHn8AeJG1z5hA
hw+KH6iovVpSSzuEr3UYqcyCFBXgPBaWYjLbsUX4kPcpGskND/1/d2ocz/WxswtN
T4bgstIp2LeiP9gIhgr5NAvHK1aoSouduLDsemAuVIov9MExvTCq3+hJ4IEH/Ouz
rqpXSQ3yAbLT3bbDDYj8Ei9flbN8J1PCgUJZY3+OupTM0W1i5BLoOsXd/MamIqaC
lU+LuPGEsWSnhRiOUj7e2WAQG6u1YBLMy5lqDGZJGFs3V2q+gWFOuwJz48340v9E
lKuW6+oMkoCcoo1FQ3BURBYR37CoxOjN5s88H3j1Ze5FpXDynikwQdUEkKIDY5TH
y9YxJoow4KWv61X2MXChIgO537cJNxtMB4lOft1Fd9jgYiFKSHNyyHfoCRnT9ICb
JrR/NVyRmYaG6Qvz+Nf4sxYxEZI3uaPt4ro6jlQ0ZaMCZmy6RWMHHKYOBpbZU22a
HPAGaXPSGqxCLrNkRwunS4r92pJXpxCmIml8xZFl2ocdZ38ugjdDfQzv/rh/RCOb
Q7JUace75A6PmIazvsW9liABvpZj4UduiOhQv58UjKHJIUvRz+hV2VXm2AQMHpDH
rp3d2AlcOzOPhpR5T5iDtTB/Po1KlzOuK4OvSgVZerVdtoAMtn0hbkNHCceEt+ko
HK07xdMlwOxjiEb+Mc0bmt2S+YVmTV33bnjLIQGjM+winTR4s4NKgDeVDVuxiRHX
iPKcjp+Pb4GcHg1YQTbc12gWvYK0ot+r2NUDxW+VQJVo3Og2y1zTtyQwd7X4foCA
0HdrXJSqnSFj4KWGBt43d4cyU5D6Q6JGPyPtx4ejPXGGJRb8R8YCxdC3uIo1TUBH
V0mXm6VYDSD2zGB6WxkNc6muGWOCuCJ9gYgSZomRVADmmFJNVAvvkQ5Ft18u8VFO
5hgguqePKJowKj7DlYFCuHWH9JJL+0G33Yed751uyAggHHghTavEA3QOxrRYuNbJ
X1vn71dH+gp5ed9+1w5ngkYmnNk817lQch7aWeJers5uXRnTVuxnU1UdrGSIzNYO
IH/rAbrtQgMgStN0IrHnsU/3Vo9mYyzNannaaPNdOh7n7BXuFUsInbG/vhCb+bAy
jsMXMDsY9gg2PGWXpYePZjebqKiu5gGaenmsWiPABX+kgzay7V2sOX1xPniIiNz8
Ux4AnePeivnnpUdbqsDg1ZaFZa4Z5koMngFHqw3Yun4ay0Y4Cq8veY9bE0srlXTX
Nok860TfReDMY5DvIuv8s/plS+lvTGgF5eMjMeNkNtIzWcFEyatvCzLTnr3RRBvV
2uUZ4HNR5a52qpjycDxsnfZRdMMYgxULvxvdnQLAEHnkieYr45UCStD6PXOcSR+F
5h5HS8XcrVvQKO42YJfbashy0Q0hmZlCj5SxEsqhMu3fZAR26FKTGicGGsaQBn76
/OCvYRyMPAWKvVlrpquAGQqMkdi3bFyGe2hDDc1I5Nv/PPSHIL6atcTyDqwNA+Rx
+yAQGxT71SC0qxCmoPbGv075XvPRrl0p1Qg3pWTWxRKTtwve+TLTqm9YaEq7M7dy
QLT8WewbkJxUF4uoHLsvvtJX97D15G0+6v4uxDKhQK2PF3q8vnm4YWlOYJrSsBSn
YN/zJ2kr1KIrUTLBm2SRQbDsxrww2/OfFmSPmPuisdTdqeTk1oGP3gA7QHDuj96c
GWGAHqHNwwvkCHZ72BA8PsZC1O0R/lTrR1fJ/H8R+jE60iByCtmlUxfPK/fj0TT6
ltges9zHVAi93TU1K+tNvPTVFTlCV8dzubziawZnEZNKT89TIsKWiMz8mDqisMp1
sqIisLhCfjYwz0fuGhqpcKSo+4VgRtMhwc4CEx5GsiQttruof/oXjnWYa2/TAhYl
RLAffMYJrNh38EMWKc06yt6+07l49iyzY/lQkz2kdneX9PMEGQ+mSep/zOdGXyl2
wEcmHfGxcDO000JxhHiZcRtxrkywM6XXvqC2cQAMDF4tTIlbrJyMpLaNFo+QL1vM
FpXsn84iVIScISYtoE8FxCZ2OAzj16TgFbKJwU4/cpHUOPHhCcVNcZy+3aX++fLb
hjAYU07SbRF7cIOvl87LtZYsF9ze2+YqXlAWjcM6MpgN4rAPjpzwwuuMw/4xVG7L
U0uBTUuoHlCQ2+mAzsEUxos2OcVOrT6NLo4y/GPoiCxtJw/rOPNtbtMPacciQ1s5
q4OLavErRq5znFn3cSVkESHwZDpmSxppTB3dzQ2/uq7YaQ/Jh6Cm8i2zzHBHVJBB
9dxfWwJ9VPZDP9f96soRxm2RmDWG1k8Zqrw//z9CjcOoj5+BldD+8GhZaLe+YgB+
Z4buS0ijvhCQDCzcXx8TbTQjv1NLRkDVJS51hUDMc0kiYGkhP0HMY/Omgeo20U+V
hdf3trNklniZff/bb8xtjD+7iIPgmgYidZ1b0GIQVXKk8USaeS86JP+jDgsZTcX6
DTXGKeVIxm2CeTuYlH+0ImoUyIlq+cnurnx/gTaVgv+Dy78CAAH35KoVZKuur9WS
9vw28tJ6YB/wLSE1rSNpb9M6Jk3q0Uoq5Jb/72rM0vA/Be0xcGy57Cvx8hB7RnUg
07wflo4dsrD6QA/AqWdknjapiXO9mTM13XtXTXs2d+ER0LKIcWbNFKcoFHrPmfR8
tgMIplQv6+or5fJmKmS5o8BajsHRbAHIuhb/dOyJyn6XlIqMw/F99qfDh9pLORc+
qmXR6kRQzjzAO7zFPJ4vNnyXygu0XtpZJ3SJ49hDBnryHwR4mrpCx/K/YlwRXy+e
ZUpo5+Oqji2RkKM27qChOpoV7PmNoZda2+vLzaZt3JR6TQluhj8PrqUkfc78gr9F
LEN75BHY0sRv5886v0Oe3fnCGc/vHXOWqhvskRmtxJeEEtUsDTutSWnsTNdpt9ac
JJG2i/VoM1VSH9Ap/tvSxsuLkoTS/Cu5UHePLwEAQlkHUH1PK1CSDtG4cYKFxgc9
75LQAlGLjbfgiALePQbPSAzS08y6OOHy7Ss/jSUzAYo4nyhHaIdCrfn8uuHtzTrG
pDfGWW9V+WGUPVwXVvVkZmTBt24tVC0RonGobEe3GXtk1Z2A+fcn13+ToktEtq8H
8orQ6aS9yDUrcUdI7lLj5EV2WPcVvfP8fSwxFc1BFON2KgSzJfUpwPYzf6ku1tb6
nqkpCHwIu5F4UhzQ7JS6QeXFRXxf+6yffcQu3OWtzKuNKG0CWJRywCNbKJZgdKRg
Uid9J7ndTW8hvlMcwsgc6MLsi4LgPiiJvBGYQMyASNemoIsOJ4HIkoujAQ0a+wy9
EDUY4Zbg9kr8l5N0B4Ws7mgYFDbPTXSGZmwfFlPLQTryVZGuFOtyk0lz6FfYTd03
UXNZ7mjaz0VCaIunNylxcKvuldfN8druPw++1F+7U47XfNZH+dCrR5OvKueCA/cq
iot8VgLzqYD8hxuwe//R1yojvH5T6OK1wV9zouTSSDfhbisLewil0Cazgv7vPkbR
pt6u3jnP+Fawcuyozy7wxDCqPpKdMYgO/jxnqkm8p2OC1puVtKdZBqJ2w4lgQEwM
7gyT3UeD6q8tmmgy4fhglfjzswws2xndpOP4EwjI8/rZdT4Wr1+drKguW3WyJDd8
MDCnIPtAYqBeJRWp3zHA+oHvD2RtenS9oy0cXPpynKdzvXxkgGNA+sBfcdnnut/C
SC1zS1l7uWyuUFX8sDHXDBHC0gNTgmvWMfDGicwTvCcZ0WM3jf3lCr0JR8f9NPjw
/24ZsIVbEbMH3kOui4z3e18q1jVePGE6gc/G11Z1q2ZpxDbv7aEtz1C3+ABkAix1
evSxocq3VFIE9PDwY9xo78HSQKvA/TUp1YED4JRkGE2vIZAZnuCPO9SM49/tgpIt
kFkewlQm+/GX/KcQV0QCTjiMKkSCmxXiR04+AmaZa9yBQOv9qXXnwJd+6axG8nBU
4/Le8DvvaX9pZWLQxZfjJGOEQIuX4bBKRuXhd2VCW6ItYOzQvq5Abwjs0Irhbtix
DAT1+EYeqLGxmxKKpMEfPyqaxDdYbaataMzrKy7sbRGRZxpcreC63ZKbtoA8X6A0
E8YJTtM8jg39lPcB+hfGKIof9XguZ//YznCq7yxRcGRWSfjFPamRBWRG4P1SCWKN
aMdufRfTf16rBuxKlk6Jv5cxec+QrSS/SS6OSFzNE1z+QqujPGkB9lkdOWA1JhoG
8xsmYjs3r21G9bGnA7LuMAAYeWHIOU8gpdl6qT3I0mUnGTxwsK5vEVVGjBDrS9J7
6PM5RsZ+IqLLKet12Aqn/5VLYrZ5YP4sPq9WpFJU12QLNjSPbsa1FvogQmq9eve4
9yottGHEclvBDWFXeJvO1hOfqPLNRpmzKdJAmBimqc/Kx0/leukxS9x/X12UN2p6
w+P3b6/8ksKP13UheAN/m2Zkt0j1oHkuhTKPmQ0nGR2THw40pkLj67OkJ3vAhNKA
x0pv2TpDfBoabR2QhSCQtjrMzj9iICj58FSB4z1gkg5KzrXwR7zrmgYcczZthwMw
oG05fcuAYo9dGBYXLpzZl/a+d1MUp9/oYGHHJm3JCexWKlfopzAQ+4QtyqjdnBdG
k0Ce4F+KmvxBcav/V7arlWKrCPbH1yFOrwulXDHk90Aw68OYtZOO3GdMgSxbJn0R
4xxpEqi3j2QCXpABU0X+OE2l/IAfKFo0/CEmfYKL3yuoOZ4ofKwDCKBA2i635mH3
zCCLPYxLHR1uXHeaa/ESSaiCR67NxHIc4fw8x97bOmgY5m4wiwRmU5wxEGf10PKZ
TxKQX4Fv0Rf4Kcv1/QAUbIZUzMFJ4sPccZOOiWSKeDZ83zXyR2zwXWVDItINWmSK
IiD1NHrGA8EWEQAjZWxQv2Fb/Ru70zItDDFCNCUxLZ/UgWZK56Tjfyf2F3XH2LjD
5RodeLUwq4J1Mghuh2ToEAehVxtQxl423kzs5DpgaG+2Ly9lJCTtlOW/Hw/+7qUb
v/qbzgIbcA5o+0iozG2sQygvdBuwoK2Vg9ULhNSHlVxcy3grsyzpeCbcQ749BAG/
rsCSjvM5/3lwKoIL5u0lCKH1r56PXkmjUQIe6Jd9YTmnIg55w+fXunz0TyrjsJYl
KbnBJIMpjuVHwuMJIe14OjJs6vp6pK4E1e2MacVsfT3RL02o4f2iJtI8A4fqeQem
eZ9QGvw/xDLrE58TZChDxGCjliCP5T3z27RbcRB2lFFS/II+2rYwAo/e/yBShieq
pisIM5i6UhQEXc0JiD5VH9Mm9vp7YbmZ6eUt8jKglWNNPUMeBi0OXzgZLZZtEn9B
Y2B67Nz6XZXyIbnMWKO8+jo/vRcYs3dAYARstOb9uXrRykQF0c0br9IqIDm77ZEF
3zGQaed1Ti8AObF8EJgb326Zv6iTSh729bx9I2JcMNfpqi2Vpm5Fv/VCLCDpZwGK
0jAQp0lFArFsl5+PzdhdMqmM1ls+wHwdBuoqpSRW4lvb1mfx6USBhpARwietB59d
MzqcADsVmB1kssxfWcZ4/hHjIfN0f2LWLjpB89R6majnQTGjFM6CtPzb1+oHYXUu
qcmcgpMLZTbXAfq1wm1LCuheHYe2vOv/Xt4zlXBdbWxJMGylPaHkkkE+F9bV6iMw
tiR6/RirIxL26k/Um5u6OZwJqJsyPH9xE7NK/lq6cwP2EyXmQUtbJooQyWYcDMSS
2z/BhHV8w88+Sge2+8HMsExWJsL5b3ZwjYa5KcMLBJARohpTzgqO74tBqb3hB8IK
StT8awyZwD0dOEQpqD4Kbq/d7S5nbMmVz/fe9Nl+Vo0WrgXAnPWwHvYXqXLVZYBg
K1tPotKlzllfMnxhvfNVeIBuAt77y2WV5IHr6O6qhb1XV9JGZ/y0Ywl+WoKIQ4sZ
HEKP9xFfq0WeJ7hnWPJ5rhP6e+RFEHE51ja9ZBH5ZlVPSRUzIWHtfonJNkIPh9RC
zsvxYnFZE/WY5qG2gPLIcwk6psXGQjiZvl+sji3LLTrDAC4uts6MWl3KDHElLZ1x
yGFF+vAgXRxSUzvWOma3r3DdAOQYm3cfSfUuO3h2GBEMg8fyBRU7S4Mp35oFM89l
qfWbYA7FSf5YGzmJ0qR+15XjkBAUXsOug9yce8Gv7P4YFbDU1o8kpRW+T/UgJz7n
vw9UjBzN8p6pjUIn8wSCHdMK2yRra5OVWX5Cxfg4uoIheVI4sXeKgbLyM6QOOp9g
jT+1tnGvBI5PRWc1YSwYqbtHLnF5R6PrhP9T5GycJ68+jrUVhi0Yt8vto0W6AKd4
cgxHiRlTOTLnAeymH4bjYyKXCChGE3/+7578buT2iI1z/8bnTDrxaTNn7ZUfmlWu
IuuQOmT2Saksvt5Az1oxlEgg/C80wJt7qwRRvFH3kHv5NpYJdwjUiK7hdBnKNxKt
C0F+m9cz/qnNEzLUspIDSU7BtHXYxaQ7F+LxXZBNjmYyK+1XeujXImWPCo6Pm9IV
0GugcVkESGySUHRjipIh2/EMVJcAO6A01nM+woHFEHtwgQZeYIqF4oUhMEmhv490
nPfULqgZAT4KEi9iDqjni2glqKTGBnQGR1nFyOR6g9Ip0rNqeghnS8LHaciY/dWd
UCqTopdx+FYAti80+JJbETWl4mek0KUJJlfJxL0dJWtK/z48oAWYltF16mC//5In
vltRmU9B4qnYmDuXEkGJHUUfzV3ulua/3qbdXb8TYSZCfOXoCUZrRCebx/AaT2Nb
mkg4xHs+Vn+EKh9oDoy9y5Naczr2YN7gROpNfeJbj7Qnl/fXm3W4O9FEzsQCVMvD
whupmYLYg5vBCj/0MdsB1NNJzRB1ZbVLJbVbIXIVBST9BeYeN2rJHKVMmVMgziNr
wZn8pkIgP5Zdie65LJ38zUDKIH9bccNEY08DIryGYdQJzfX6HaV9so+OkD9AhILb
Ybw1UPsKAVwrTdBtwGAHhsVb0iYwyGObNFgFVLbvuxi+C3GfoIuFMK+EGyaLWP4m
9z7+vUgxFDf1TNkHJmLjqmR5JtrSHBBuPcPDSlUjiZmEDU1/TpUB5TiPb79Peg/B
s0aF3p1nRESMHV6KkpflHSdg5pK4gmpR82KGD7kzo412oN7tBTFc2SpqDS6Nfc1P
i/GfZxxS2ZSUJcbM1fl3x8O+1yOrvP9lYqbF6YVnNzxFXo2VsJMkHFQBx/xpXt71
EdnUdtTRa+RYHUmp8G0a8EnNXnNK0c3zWpMGloLlDYLw9/8ShSznO9t/jMnArc/4
+qKJ1ukG89wmwUzsKVWsg/RocTR/TcAotEY2roWQciec7xtxuKH9wrW23hWVNxV7
+lW+uSww9FVGdBd5fg/YHra4WsdMphaduIZS53XoN50mVnKGMKUk25Vq3W91tVaK
/EP3423iIosB2XSYSPEwxgHa9MNINIG+fCsvTqPnHsBu+k548QZfSqGkwQ2WF4HP
FwFcoHbLpDCCjBEs+H+Ny3JuA1wx8w0Nc92Kpr8twJOKGPH2PCCLz7ATfhmxmgsg
eYuKaZbP9wz2fodoIQeK2LqiYqe7hlMhWlytBP4khxby/V6FQcW/8EPRBR+oRr1g
bFgjHt0Whxm+AWC5PwDhXsHSmHAwCkiWQiTTj/ukTbkKm3IeSsg3W3SMZrXoOus2
g/vQkr51o749MeKYgFfVR1ngkPRLAVWrMX2yoQeY6ZIz0/5iL9u/x2xio8hKrljY
/LTz6YxnKGhlmFxA7q4uwL29vHNUFp+i7w0dB1nQaHpBUbGGj6WK7pNOEnfemjp1
bDBzF+yr1paK8VELIetAo2d5+n6ZnhVIhSjceLbgUaFwXIDcG5lbCVFEoTE3H/CY
dPyqzPX5HNsMmaLqQEvTCxRoic0NsWPE7K9oma7WFTvA7pHnxdZT8GPC3gldM1tF
Z83PjD3QlW6/RVl8EXZ3p9n1jEm/woJ5oIk3JBweGxBbCdczgwJ7LrcHFRgTLsUp
/IN5acQqYVdsYjHP1g/c7w9pIFh4+cBlJiKzMiVqL7ocPI3WLxdeX/MhNP4HN7d1
esnbX2rYMO3KYBzbY12oR/P1TBQS/OTgoH0BrunjCvxpnPsRyYVe/UXLk4bClnmM
ZCaym7A6lzINQ1PWLgAKuP3KANW0aY9boSf5M97Ly9KKy7iyuXJTXTB88CTS22DX
7fdcby0E3+8f44Tzp2FddnjQ/dJRIpK34M2/m3sekoOvV90SaHOjF4BURh5S2a43
2xRJFS7W02MO++6i8dvZi1mVlveMW82CDUV7QYWWfmns5fzx1p6h7ZRDOtsLcGF2
Mu4LU1p04CrL/i4F6zrFPcBMMWsQWZoeqGcifR1bpmX/VjeKyeBYSqZmT2y5OSsE
lL2t1GD1co1WqTKF52XLLi3IKfArwLq1MbxWmE+cJjBlHlCHg2VuEzYRYHX95Ego
HE0vocmnGzugUQy/5dORB3KOfBqXAALjOUDQXgtkJLY1sMwPpmq6Jv53e6act8gz
JqkYV4oTTP0XQLuIwztwGQZZVWFQV1wZ7Tg1U9OAq2awgmhjvNwhs407mG/HOaGe
Zqq+Nw4nuStj7jFhs1NtVAp3ox90bXthvlwYUiNKgH3q21WnuIWkpKVwibdg/9bg
FPEF1qll3J6/3Qbv1YKngc+3RfjgnlTX4eOtCuVfS5Bq53f96/DB0HMOXdWs8KN7
xFJ9HL4DvBSm8fCjXmxla1yECJHIm7Ag9Z106ogIinxUbNsWuSTeuHVk+dRqrgdy
Xm6NT4AljSrvgt5T3h4QIXknfYg7T/0qRmGrSD/L9br3few916np0ohYtIEbaFUk
trMVRlm8w4wyHfIyi3t4Bm4HtYarnwDJ2jJ3x9J08RvboruTD3xCw9AsW+dhCpcd
yazEa97iukamdqLAlf4qvLKpCu8V1iUeFzSqLgkhMnrbD28++vXyiWRL4XPut9hK
63U81PzcZdjHkTglUa3+v4YXr+eyAi1Fz8St7+bsB7UYETs3UTGx9E/CzHFNcPSj
1rfaK87XotPCJWEcLPCE0UmqUbBavdeGcst2LkmThCrMyDHYJThZvaMDm1+vYVvx
+7NvqaIUVAiBwXORWQoAzT+CUK+OdFuZA3jSaLe7GiQ91y/tBwru+1dBJITF1KKX
62PmvtVRv3THu9+Ip0Ei2tIVdfWR+WIJY09z8jjyS3qIj711DzPB2/mgWgBz5aZe
4JtkAQ+uuWXtkEArl2RsVhl2uWLgbyWN1XUaB82X3pM9Kg+o/CiygT4/hQ/y/f1s
tUdUZzZT8u2/XS3TJini7Jdk5RKVNOZVvit06/05PQf2Q52NRkwebxtccvbQqpne
PZbjAsgOS8g9uSDIEbzZw/rmatrzwT7ZAnQ15VV8ehlY4pWieldFFe5ANNwXWq/a
uy9vWXv98rG21rwrzETBrWLHlL+CEpagmBgdh/2cgBevThC7c0IstZmil3GkVAL7
cOaomTovXcUqL1fwqE5DQ17Sc539f0L/k3IMo9klR7m1E8eEAK5VaBHBeb352T3G
xtDJAN5nt4ADVIgb4n1Pw2znG5+J5dca5y9WC4hc/2WJbbQ5jWle0BCS5ah5UKdu
ZwQvXjVNEMOUJZ8mH/I/kXbk+Hs5k18BLoGvmBx7Oesq5nbtDIc+P+9UpdEniiJv
SIKLG8lWnfa03BVBKsfi9rBHxKDpnPaDxwD0T5JDFQgMZFiC5TqkHdygk1ckZNxX
Qf/3vQvPsHSgf6Xyp9KpRgfQWxok3ZkGvR8+P07DmdVLhAysv5SsvWuV/6+Zo6he
GF5C7mP/WK+K1KHFdPobvATJnVztmE6lDEl0yRUJNTTicSCYFP+Gli94ew8IvFts
EzZv4Lv5jkvGfsB7KS2gtmy9NxhZAz6+apbLw9uskFU1iQ3Js+MAj9bl4451X2Zm
MeT27ve2vi17k2KpXg0L61U91DMukU/PBD3EtlZt0+qF0BXCW0Bmtu/Hn0rzp8wR
quUnl+08t5HthiP2TGur4oeWgz293OHDxS+8rnXih4DZTnrCL1GBobITKBuPB2+D
rAU4wCJlcYsE0A9huPZzLYG3q0nIK7PWE5GBGb2mZ1rs/jh2bwjuqex1fePxfwTW
ZI7WopjXf7UI8dVvLLwPCGSyu01dDXeCzFC8iuUdVik8eXLFxHCgzQ7y32r9vHWY
sOosgDdAYaw0vSyHOs19gIYxTU7iInDwJtUxDPVGpsgMdCIjNuOEyIbySEw4VHpC
iIWmV8ZNtmhOmvKQ1PtihOApRCLcUZyJi72b47FlYYQa3NW+ijKxpubJlSkZzq24
ZoH9Zu/fA98DCmTYWdZ/CS7gvGxYitM3EobF7NGHT90Peuml/EeWwR8YFgWD9End
prugIZJhc1II615A4WhDV/zMIm4zFsCr+NDER4IEdlXi69CYjGsYYy5WElJk6WV+
4tSJU2BwUChwaACeG4MYZCqqsk0pOKRl7rAI/5k89IIMbHVD6WgT16icsw32USFB
AdlNE4S4wOFOuOfFLvhM0w1iSMI4xNKXLJPijmBFZb39wh0UlWOsoe808ffk52/d
gh0/wo0O0N8I8W16gmphhm9CZJIDVdMIL8g4d+4lchT16TYVLZo3FgMCKVQm7i39
zmMAbonShCPn1lmo3+GEZGDV0kVzo7M0a4WdchuS3K3I06XnExmPwLjZR1YsFlyl
WoKMPnl8QI+Y/SYmbKl3FCoZz8iElmOmJ9Fw/obzt+En20LQGBgEGDTAstiODg4j
bzjK+55xZCgoZF2EeGIkaNQty0dPNMDU5lVPwbc0sTBwfKIiuzRvj44he8VgczJ/
4IrVIX00shgN2v6t2cICnqwFuhvnhe1mubqRwDgF9+W0Pqe2jejwTU/20ouEkmnf
7ybvfblG6+OymfgshFdKvn6yJbwNMiAjuZjM4nmDA2cux7kDr2R0lmTHWanQ+hju
2V8strU/UUHLQPihr5GJeqGQG4HSkLAeOCbGbTYCsuhJRORUtBsju4FmtmPjK8g2
duPlkXzKU+DhvihZXepgQ5D9cnYjhBdg4fFjZAnlld802mTXqdoINBnbrGWyQ2K3
NEQiDQym37QVWNLLRkAvX0GdU00caLNA4r0RLF3GKeFRqK07vmUI8zeL4AVYn13q
AjhBmhWNcNRQ9TjnK+/qRjMHG1fcfoBMSRwvokKjjBayKRYx56AeHC4zx31vDNbp
WVe20JaVWjCeoeEVOZ5xCq5gQjjCKdiSFoq83HKOXyl7gJUbqWfyg4w2lBt/0M44
RA3kfjfyWskUDDFfTyKKJOZBF7oNbrmJWY06MQK9T+i1vvGmw3h/gTEA0cLlYcWT
xWeSUoqcv3zdUzFmuXbFXnL+knmnfREHwJZ0tQk5wxL4hoEUGxPqCB5k2nG7hj7s
fy46clKaUGOAFGZA077aAqqna/b/4vzqLm/I1Eb9bUc5m8RAmh415+eaNnRCSG/u
OsRlvsrhFAQH6mfuULz8FyqLidQoJMGsSBx1XacgAQcyUm+2WlW9P2v2flLsBY1O
7fbZ/esQlDKSAroIpwMnIDhC3qAUnrfHpFiFjsIcstOx4zZt+AJbwoQewiB+Wovf
m3QBHRzY4erql/aSEvZYQSiTaJ7R4Osm+bur72NZzoVnVoWH2mcz7thdG9l1irxC
rYcZhyU3pQVwkF3/levNCJh63rLNyeg7WoZ0g3gig5MqVsN7zHQqOWl7s99IwzlP
gnPI3PJEikxtvWk8azu6/rns64z0SE5FZgE+RLBtmaDzKGJZ3pYAa2DkWWNhj5qb
OHlSNkI6YMuSK8JZJbvl3kurUVvEzbfZBcsAZfrUZe1Zq2gZRpxSAsMii0G7BCj9
Gy+51NL2EwSvFO2uXIWeEXGH22e/QL4pH9mc7/cNuFElZ5B9wbOD6OCv5fJhMPpw
p5tl1YWV8Vkk6vDvSINTZt4tDagKRu6pw96kvXynJp9M33oi8XF6KeGRUki93//i
wNErnj7aETjAjat4o4nT+1bMi8vkeue/8BzI8pbE1lhRNZfeineUamdxYKk6wO7/
BQ4l5VyQXNR9qhwzbEQruH03W42cADVQoZSZGXf4QEf5CACzOs79R7NPJeDneJpX
idxGNxLutZ7pGcsFJLPvLaqsKVkdngZakavociB8yKshA7htbzhmSQI5QrebYHSD
RF5jrVETiiW68MHJul463Dp9MqejspLxS/R8iquYqdGn7doe7Lp8WtJ36QZchQ+e
kP4CwsIXlSJ6H/xU6+OCxQNnpHNH22FIOthFJH9zU5GnK7GmZZKo96fbKCFgZ73S
zCflzAKWq3exsHvT4i5noLUipX1pRACM94aTmE+JvFK6jn7TFDdzwv8UzCmU8BAQ
U+hpGnLejz+NFQFk6h6uywBEzl5SyUIyvRyS/7PtBZMbIQmSoKkCMVtvxeSiBP3K
1ehPxSSo79zxlTNCUPA46xjA6P8IbxOCcLs5jS6EQnefLZOLKPI1CN2yKPoH6Fyk
FCqB4wA5uBr7/vbyrIrcim4tnaQidKL5IRkfTcDNqO0bjTNj+JO/023++/C4XmV7
ZnnIWHqoxnb6IXlOX/N1NzIG2eBPL/wFsQQ80h3ijryGq+Z9Y6FPQlnrn4N5b2qV
/sC4hS5NZerS2qcTccTsX7/xaje5utWXmD3q8SYWnCdv5mSGAEe4F9Mi2FPoz++V
tu0MlETkvGkL4u63B04S4vMUAA7oDAogASDKieMITj0ClHpz5U/5G+DO1Gn0eQEa
CZFAMx6jspHB82L3dM61p4YD6A4TWwEyG4TdMi6XBQcyvWF2Xlz6mPbITzhhebHK
jGHWWvqkUZ4kwD66/WPAbZ1TFLE1rYnHyRIASrHuA0URk+K+13iQS/Axq2MO0vUk
9mTBWfzLqZL5mi+RAS1CTxtbcP/Y3p80LkrAJpZt+GVEHZKVkUu4cufrUq82R8f9
27JHYyydux6Sq1lqZTQ9nZxMT4SnykY26WUdXrARyBAEX2bFBYrF2piYHIf8JWlC
dBHqet1anO7hmPHbdGeAXgXPGfSaeX03HAzHL0om+n0RQ5p25lJSJTGzwwR4a06+
VMYDp/tq6LZFe9eO8uBiucuqTTkZ1Egbi1fjnCmehyZAUQYVY273dxyAiuUXamS1
UrgnDN8i9MuWC9bumEM8b0aIb6OxFMEyJfspdbDcJnOW1ui7IAfjokG9fH9d9k++
CKGHuakNhSyDbXK4KqFTgGIhYoL1HeRxUDlhi9kXSRkcfyo5+XrZdFPLJFvpZDKA
8nbJaIwZyz/ZyCoARYbhKWv/kfcWuTEarvukrxMeeJK2PFZjN9Au9e6nkyozDR/C
fPWHmMUCOt1xQk8w2pc94X+ZA9CDArm2nyYRdcPVgmP9YERmiBjVLUscZh47keDe
llnCwk2OCnuLll0ZzQbQ/vARUdEMZCcDPtZvozYdLTWJIqa5vnnMUsg0rn5Hm0f4
Z1L1Mqrxw0bZ6o7lA0iEbJ8nb1yNw1FLhyHQ3Sr+Plb/cybbPKtKElh3P6kj9exZ
04PO6BIx2USRrQqvjOUcHWlhJnFsXl0chbPHTVAriT5W1WUv94oKyN+oqQ3Fk1Xy
9m2JjAbbV0BYgiQhEq6nvEfVOh8j1sHK0v29qskxwrxHjeXcLac2K9jWsbytBxi5
rdLHi8+UV+jDovgocsJSUyhAiBUwxqVdvii6+1LrmbFrhgQg6H/SZbNcnadT6POL
gkipozP/Y+0uT4E5Rqi6F3Lod8Dnj9wSNO5hsIIJPlzc+7nqSz1MnUHMFrtrs96X
qyN5zczj77FutOrO3CWRDCzwh4ah82axfX49mkUC0rembcdWSq91j39S877v8u14
SVbtW/QFTgFgrfOp2guMwPzW1JB+czILMWJdjFc+3jAeBw9DhhR2peSTpAkjOkOV
quB3tkvQEuBHLu3DaLpUcxvXI8l26bbzr1pMk43Srofvbm3QW1OL4PiBNvfbGvWB
F/w6zWTczJmUXjjcla2JV1okEZM6jyC8hr9E8o2C6V23/r+gkYPqY+qZ8/016oD2
0W7B6rOa+b7GypechwXAGFLftQJNBU9kiIja3MY/i2zkUsT/mpIltBpJQb2JuUHp
fHI08i0OqOTnmMEO6XOR5VPe10cCm3LB7wMee58FVRjuEVMqR9MdBY7XQ3w3Or2V
77G1SL2qcyFlLvx/7l008fvGpLPxodPey7bP2kNJmvU9Fk8yLMFsHzMB0myfhOo4
OA4gp3SZGmgRe+k0iqcxnWxgobGYBgnRsWN6XyVXQwJtczXVGqQWXXn/XM8qokmQ
gHnAX6LfEaDyB7DiVFXEvC7FrlG3r1PRzEvDVd68jW97D1wkWXZ+wuMLNPRI1kQb
MicvWXHx4Pxa2HxVOZ0V8xL64iLPkqwyRibgj8pD5C6jIxj8wnL/fdXislk8DPxq
fpTMaFXTfe5xF2wCLPsI86TfkC538TRKc6H9/bhJhfUKWY9f5QlF3pukuJRqlXcL
rE+XlQSE7p61cBMZj1rES7G2ytuVhc2Ph+iVZnZT9FABweq83xOPgRnb4EW72USH
wCv4fjTzaiC0WF0YNyNqyfcv0K4W/8udn9gESi6IWtoJJBsEahIeGDDuDFKc0jes
lQ3djNIl6QbdGSgEBQlvFGqUJ4ji8DKc7ONQiHhipPGeWVNpGevSY7Q0Qix1+a7N
BZgvmmA5NuzYd5HiJhExnBUtPWAbmJzwG7Mr9mIMnjoRUZlUm85DQEq3Ni+negVd
Y1E58CGr/Kcw28uCbh8tkYXdNiCTSslKkPsyVu+TmCdFp5rGIWOU4rRd/QXs8+H3
eT9aVMzwPs4k5ZYmf2Ey637dU0gKQD1n6LmDMi8XPYWhUhASfcv5bBto+KRYlP8N
eDvYMNGS7DdzvrsqMwdDPxlAKC94+f37H48P5xh1O0Vz/thgl52rTbelDNNrIx2p
D+jJ91fzHi0pHBRmGj4Ipv85QXeBKQTHK5euG95JcJIHQ1Nv+FhvSH0UCelVPyeT
Ywo+6gCxaiSTKKUZuXDbIkA3DZtqhQTifG8L+G/3XK3PvP0ZO51Uv90ZsZQfuWN2
2xaVxiY73/CzyqoCskR4a7eztSAHVx4HagWx1uPHUUiX9lrDavQBT9g3N2Fub9w9
WgB6O1CjgEsZM3mytYGmNTmJajbbhySILgF4JY3GepL16rO4q6MwhGjSva4YZGgG
myRCPq3O44F3iUZNKfgITAsDriGqNpSAiQuiKvwAm45rl2M1cWfr2AdmyILbq3mv
iEgn37q/PSORzLe7GmlaIPuh9tOm47ToXoI2y2Yks+9BH9S82F+g6UEC9egJJnU5
VoJu2XXBUd0/ru28PRAIaMAs+FeKvTfyYd0eEg8aMlv7KnLeWG7KbmxYtwTL3Q/5
Jp39B5A+hPB4Pds0lt0am2bCs45brdVJYKwBxifT2K2azNET54Y4pmEe9NIVjIFH
5Oy7BTSnHYCrc0bnWyMuJ8hfF7wuxtvFp90bylhBwKGzx/TOX5cA8axhG1VeCllH
ivnpsCcOqsh+iNl/VRtbkqhRXT5ObpiNzTe3sJZ+OZGhS4liylNm1RDWy2ZIJeNN
6hEleB5d4QZFt4bDuoZwH0M6PahdZtd8dXf9+nNXV3FjZLK8m9lJxyNqvVDmOGgy
X+978o7X4aDlWm9ZVcQkzCkiPec38FTwh3Joh7q80mjnsuKRmzM2M0bBHQK2OlT+
D0Ki1bG912ttOgO3eiLXmE3kw84VarIELApSC3ObYjISMNMGYqBB5HdEoT59OAgL
sX0UXMch4r4BuG846agLoJuvoNiooobrCkK4jhtrB/lA2VxsliCj+DfSpVGmaGg9
pzPwn4gCHNcs612NXfZQdGxWXIYDrMDpJnv3zAdD4C7lEwkeviTbTrST4yppKIC1
EZPClBlMnzkfUia2hQddzzwgmUoQHj1bPx+y4GNIZftlSPl9aaOnoUDNP83MvCtj
YLaV/QzF2OAVYIvFfuq0Jzs3J6pL60kRa7y9hIpstID3SYby79/aH5NOZAhHWaUM
1uR4FlYJ4QiO4R9jpB4GhDamAJGQ7RPJfmj6OMnSTUNm/Itx/jok8fucT9NaNB0L
5Mgx47iX7QJqVCGeYVrkNoxOYdEQUuINObr3y4ZexBrj+GzSRX2mdD3gxGNtF2r5
dRKpc4ksP9DMmZRj8jieh7wBhaqraheQa6lIUNn+lUlifhXPFagXVMVUUkxhC/bx
mQulZUUA1tqUeghYvqrwNiv+WE0ezY4ve8dBYYnLJgEq1yE6m9hLECdzEYPj1gqJ
GWKnqCDF6Wnd1GKhJN7tdcomELc4r234IsThQVS+rGgKmp2p0BCBGkQnagnYo2bb
UBUdh5jgnVgSPyfRHSJafokgp5ZCnmXoebRjzvkLKwxiEy7N5kPh+3Nws+0Z+6Cc
fHlNHt6VuenVwspK5TtlXDsXFL2Dv0QrhfmTHFq98b1nE+9uLoEfXSYWzEIL7ul3
2IsrwzIOGHSJr1atIFdrt1JSsdWYsK+mlHxzu2Etg15Cy6a5Pv15dm+v6yED/Z1H
cVCfxd02rkMTjiyI+jIUgVOb6Y2r8OsY7GKVN+93Lo+fTRc7OKUMJBo1qL3aKW9v
2FSZna7nk1oYdtVwGmyg4XTMjSgRYysiRDjEuEjXYzHqyfk2Kp66Up0//iGcDxky
I/pr5MTdhv+IWO63zbdW30zm8E6phYeYPwmfySzv/lkPwxYy0i1UOICNM2IcaoW6
9lnBpQBbQSTlc58mEERDEC99de/hLX2W9ebyWisr6R4dW1U+V03OGygxfutABIaj
DxPGgLbxF+MHeFmdV9B/nZX77ZGfZDBnjmX1VLJd5XQdxafRXtE+X+DQsLV8REJj
FOKjF8EXjCEoQKPioWPRvP5sqvhFkwzQTC2oWiQVU6h41zRv3s+R41BQRvysZKzu
eqALpqPLvU7nrI88q5l7v/YXP6F000exb/n5IevRcaibFvM0Dt3kKBI8KXZoaEiA
99c8stOY1VD/x3mmeu4Ngl1yl7jd6jrenY3aeLyo/vntP5yZ76p5BOVnhgDSc7rz
yGC7/pwlGseFM2UZTL/qcFxiGs7SVWMh031W1pHnunrlHZO1kfEnM0lPuUdGBzmu
qk1XzgMCz+5O8QTBKNvbAbKZCYZMx+PrcIrUpP0VIXEXHLTLzY9ZQriyxTwKQGwc
tnduO1bblV9BIe0Lw2pbbDxLPwdzsab7ygpZ5oGjM5tO/dIsTzwTmXNWmadAxGeU
zoBEFS3lzEzyltuK2xwKisJiloL6+IlLDi+dXV1S/kwNVFyVevclgguGFTeBP8Qy
ZCC1ehlmKnJ0GPKHs/qgDhb9cnEPUHdIWH+db7JAKlowN11qhgONBygV5dj+sC97
Mg/KeSPzQQ9UzlT39yuzKP9qz0QQkS0HGy3T6ugn4TBEZOlh/pw74g9EcO64lt4A
bX7QJPZvGx/P4TZgzU3n+efCjzSn9N9vStHA6qjCcyyXqlBL7LRPJC7WZtwUWuuE
hVPi1sSf4qbaE+IVPApnB5sg1NR9mgJGkbctNFBe5PcuoxyGcr1lLjbpp4C6U32i
J7YV8emacX53g9n2ds2qKNFsrmuYRbenD+atJXJ3jbn1FmDfvlyTUm5fSamMdfxh
yF5PgGYGdTuByR0t2PLj/TEC4+ed8/cN0a5xZ6URcaIl0FRtFRPTcPZEay+JEVpE
JtKUrUc/DuszLyiGP+zEnXY/UfHuA4BRkMQ9RV7mWvUzE17vQGKmsz4URV4eUvDV
m3d4Z6P4sj0NHEZZqUEwCkCwpVskyJzgSNi8mGkWEizWfOLEefKABFr9hdzYE5cK
Wn47pJJcM/Z4g46/K/1TakRHpNCitYUY3XXyNbnAtJkWxCazvAMz4MSvAlOXvL0A
TsLnK9CCEB6SFiel3MzIzLpEvf+MufwKCOAsLXSboLNr1+0d7toucSiaZKwsWKZb
HiH/XduZYyk6+b1tfbVIRggG85r85s4+BvL6tgNQnvAuhvO8kHurh8oO3iGJDyy6
03+GYMRIpAqfOeBAq+XrM2Pg36ujc6kwsj2Q3nldqAY1zljCqXVUOYeYwUI0ZwC2
KQ/6pgONuC5VjqYdd9iZrMg2WERYuB3Y2W/7HN8VhtOhYEYGD6QO2QJz0kwVCfAC
9Bb2Enf0eLdOrKkSx9gSQuga9aJA1M8NdE/YNJ5Rv9WK4k07mOV6fYErWGDgLiOb
IdxWK0wh2rReEwJlSB2jf6keLOWd3Iz6lVIAUgGZTQ2cNdVx82Ot2SKUurwUWCmG
VkeocQwwMp9wSAJVdLvE/ctJh18VAJ9qwkefK9EAFoEvtz0MECC9uiOsmCNWMdWh
VB/SrE8pw2OJTz5tuD22thBRB93bWiBIbYTIMdubm+boDhr6iy6r7BLQ1G5wPSif
Fe/qHnxvk0W1ho24sZGxsiyM3usWHrwOZi/VbN6YrBnBKtIh85HH6nWCF08hwY7C
rsxz+3EqpxufBffXGX9BW81ss9GqJcgzBvJBt+gj64Q29XbcV2WLvN58IUyDfeEW
ngO8zmykQbtjRftqDxEO2COOkZHEcL1E6H/6FncC2QXbPykJ8QW+6KZ7EVrpXiC5
xNgDnrTBqY1E3u6mYH7nu8vFdWcF+Gq9v7OKIm94/+1Yencnexj0+VC7OV9Kywc7
eNpxPxHcT/YucfwJbw8DTUHE87ErnQEMIv7wbH1T0nQMg0W06mc1itetVVSwsN0j
KE1vq/G2JBpmn1pniOHGxvrofTDed9X5qXcehLCP2nrRADbu9xjIoEGsVby6d8Lt
152U0O5z2ZdiuU7Oq696pXIjU0d6gnB75jXpSOPLHqW5v8ZStif8ZO9/ra8oTN9B
zbKXFWpovDTn6Ksgc3A53jAx09oUB/bWqYz28UgYiuFtOmScymlCS7ILrCzhnsxb
FNCk4619KMuDI2gHbb+9UMkNMxuvCok2axZaWykIbPEhb7A4fAT2G5JDBrgofCbr
/C+x35MQ1qv1l7l2W1tKdqjynonv2xjz4RqF3pg1IuyQC/bmijQ5SbDBsBQFtWTF
z4hP6hvDsd7pyzoVrROaLFtJCmJGe1fXbPH8IrFPraHbVCvHtNGafmKUWH3ADfY+
EN33XsW89IhVyp4VZItypi9HSRDuiVFKVetD+26FeHPKs1r5QHBb+uoQolmiZpl9
6/7DeY67YzRP+TB6nj5iuvCI2GHXEMCNmhd5inPe+YXy9s0zbR9FHpsOCuyRsG+7
4le61xZz64jVEeUwMXruhEcOP2FVlRhQQywdzZnws3A7hPiDWOkIj0ICqwTPcT8j
UcoNTYfY1hmjotUCcxrFWbODnsoVbTrBX5Sb2nrebaIk88t61rJWyH1hm9r2G/4w
ULRbp1IXFufK9mY+CrvrdTpManTNmpXax6WBjH1koloStQcYimFRarw8TqLMr3dY
rjEOsH3dLRoiwSFdV/7mRbmhkmeVnLJEhM3hshAOQxARUPIPpj5dPyesuEvWU6w7
LH2YdQ/feaieNp2LoBE7uL9dZAlPiCLU0YWOfXgKQBXJoCGfsX14F8j20i5yrxma
D1Tdz1zd1GilBf67p5Yn8iOzxkpoF23wbhM/LSV8FRf/8OLIDRnjEwcSZvejBTeL
u3/xaJlHbIh/gRB6L7zMsx0Vc1mXE3DvuIRcAcc9dLrXb9GVNx8L/imkZf75T+9w
2mFITvudr9bhc55p9brhhnwSnmmsyMarGAx5mFI05J/hlzr80xL55necAZvYa3j4
emuT0NE4DZ0M7USYQ/n0+LyVs0corTpYicoCJUaDvd/Dr8taRMIBmbQkPVjEWCFY
NlVAgKZn5bim3qpTdhPLNJ3ivF3dkF5zW41G4o+4fFxRHaX9/OaGKV083/YPYuwj
ElT1G539Z6LFp32VBMM+ULSkz6SlFo8tI8XQ2A1dcYggRlTtCLofHC4lhlYfh2wK
fmNRgEGUn114mXcHs0RDp3A3Au0ScH7AgYnHflj6GmQ2501k0bfiuw4yZMw/UxES
fm7Q0p1IFbhhvC6wSX20DSM2ItEdj0LPHFKw1yEa3/S2Ryk1NaEIAmJIS/cttEvn
YDZQaTE5B0ADlR5UjR9b5Og+yNzi7GAaND+/i+hRQi65IclDKKdGOwjTP7ld8TlJ
SlQvtW0axDUKQGQfOPm43qWPvENFzWkxHI+DiAiVVGEQx9h/zxCEJLFihQARVdAZ
xNlko4Aj00ISdRwyZPvqaX6ffnQEVF3TY7QyE6bY/PZGMWe1dr1sp9yiZwLL4e/0
Qb9YnMnm1lJAQqIXdiHJxi8XJ7Ir2gKs9VOOpugb8U0S4SQAFbf/I2JIpkUlEhFv
Qvyme1xNy7P4LmXJXl/yBgV/k2Y3lBZ2IZ8xgfnvb1bekh20gNrKeIvQ10IJW07Q
6x9XjVw1VYcCg8mwwBKDcE05o7a589lVbtTickpR5TWnRJVfqyMKrUGlFof20hHR
Sm7jj+BGnkth44P6nu4SayLF2vUAOVKVesauc9JQJdvmUZL7JyhnhqO0R1Ko64GT
7i4cVi2Ztq0ILP6WWcGx0gjFPJXtm3I0eq4LDqKA37rbCxL+va1cjtCeuuPjRD7M
IVmabUy9Vjpmm8OzfbeqdohQgRE9frAxQPKdhTLF+yqTP1wG5+Swtty5cMXfSvG5
fEF9vv8IQnzESMpwWBeHX5PkkGTiQrH8Iqcl40iwuQn+EVQvIIu5ezUJkEXIUYeD
dNLwHetOTMiAdZpB5qcQW1dT3W/ZFheNi21h3JXpEqG7HFyfQcLSWxyLmC8zcGUB
3dKGVUvTbgw9np86fSwTzegyQ3xFGjnDxupndcvlPYSjGV8Cwwz1MLCXtr7gfDTf
EzFRJb7NwDTIXIljef0k37HMGg5JPxBwX9/9i0NemMUOKBqR30vxD46dA35VzScN
+JjLl7V94NcDnaeSh58L9IXBfRwT2cEzg6SBx+fluAUZCxf3j7wP5+lIFY6WVqbl
ZV811AHgnyzjmqeT4AhnT6S6D5ryI2uXY9n6eG6pKtC5uW7L6itrj7kxSenrDZmr
atTmq9fuzAPaJFQuAz2FLNno0S3+r4wlvrQb9k5RtQ/9AokqmXf523GZ3xMy/G+M
clfzGZSYrzUMG8l/SJMlQUeiboElJxMVXk/hCyABvmvvpBW8eSqb6Hww/wnvaGW5
q+YILDOb6D3Grma8dpKTR7jbTPyQHoPXui7Fb+NATooUsLCZf0X89TF4j2/1O6ho
2XCrK3CfUPnkofXz0Zco88QjICi7pl2nDz+q5hmECcTUuARdFNLYNTp3S0lJ81lj
2KRh+e5UsmNHT7BwWzUWUVft0P0fhsfrIb/KWWv5hWkZ8R6HmtNgl7IrR+GETRdg
EMwzam2gj7GqS0bZJyBSinD2dYU3yKJ6LBeXoQtUA14Pn6hsSWljf/lKA4ZgROdK
bU+9Vpx9LUhEw2gs6JxAohoLcdB5WMGtREmr8dgNeegPOwoEsOxfMG2debT5Kz+a
EVSjf7Ts+FEWQ7rPvEUiJ2xIMNQOaAiIjMk4jEGi4ORjChA2Yzkj/w432rhhnnhf
oOulspQfaRVEY6tKVmWsspPtMcYiJr+4Ko1RB20EQtUbSnt9XDcwo6/PKWYTDeIH
Kdl95eSWO33PCXJNPOK0oFpHERg5hQ49uAvsFA0kh8Gz9TGRHuWdR9V0dfWS9EmQ
wZrgSk2jyiNZA69X6ZhHWIWLOU4+IwkZrDdCpd/pIGf/dcBvuTLj1qf7uWk5MoxD
w39ClrFB3QLAd/NqSF+hlBZC0go41m50J+3ADl3IpKnvBhgs0XXdkqNpNAoUf21n
nLvM/r6TQZ+htlKSsU7iazYuDJ+HY1nTHCjqb5bY3LjYNObdU5PiH7CwJA81AgWP
QsXvu1n4bdEKYqqXgruDfs3OeJh+LWxAA8SRwxK0rntvjsNQsClup6r3WFQ09rpl
nVm6rdqfMWRgIIe1a6ukysTkwKGpm+p3ouEHSBbrXP/z7wuINe7XYHvfbJhtd5gI
wPGVn+2C4R8s1BWla6aYpwQLwy07XgUjvYRPC6MYNKfVsiQIc0u4G7VGQ1vW3kfT
9KUCQkvYM4NYbos4ouwcmnvcSQEWgQRrMl87Qr07jcp7k/di6oyQ1xC6MrM8+g0g
V+AbiJggQ47tDYAvH4dxDQDjN3PK5qTBJroUeB7eud9khWnDWMMX++dm/wOuW9Rj
2vciqj4d2H2c7HgLF7nznXLZvPErgp7ivyRsTPx0U8T/bYWjvdzFPuUJI3PxBaBM
WFnjjuGNpk2unvMKsUl9uU6E0JLJZ+UBTSNs670OqSIw1LrosNS96i7tnU8CY4OD
wSUuCLE0agbdHc4+bBuIRPFKLx+3uZM7RaTJRnn97dgk68IU3TEL9SpLAjxvfPVr
D3C6Zb7vd/kNIKdV5Kr8wu8fnCYUJKjpodTrNZdnyuUDeslDpf84UYCkEG5/iJUc
f60+XS+MteWabUDhPMEFkqjsFSKr8m5mlNjBLKkGOcXmRPUQBKkHzUM0ivtrF1h0
Azl5cJfzt7LSoSzNg7C5GPJEpb+awM9k+Tqe1qeAWOtXwhvpfN+KPwBGVZUTQiFR
T1IUcpe3Vhy5eQ3V/P+U2CIaPv5kP7mK4Z8zQJl0Wuo75mvpCFMbcD1AVYUtzipa
y8TAYPiq70BhgBdyx95s+5qMrIAExR5APZg9kNRNbJ0G1ArTX9eHAd40lZayF4d6
llL5bHD8QbRnMQn8iHrSAwv7yZSowYgXYoY/jqb8X6ka/byOn7O0XQE2Xw+fpTfe
fIM4FicwFK+HUNsbJ7pobXdvJ508lNZaw1NngDXJm6wLBMfCyMZKe7bxBEZXlqdm
wXQAJjkiI/3HLJ13wNUscend0/RUpN8qVuHJUYtEHNb++/b6xI2yX99Aa/UIJfcM
n+8QjymJgzQK5hewcNZ95hVq2Md3O2SMgG9GB2NX+Lu8WJLbVf7JCMW8I+AUvQaW
1pp6IV8rqYT2v2QXWicvAwAt/VY+PXzMfW6gVyErcZXLVY6ELnbQPLHlFoOQbmvY
R6LTisA7Z7jB5VCJVmeCKNnFZWYQBbzJsfERTrZWIrIN/DaRKvv0kc+5iUVgzC5M
/5T94YhNUkX0YpFkkuvnPaNhbsyN1UB7cVIAM+s40E8GnMo2izD5GkzWZRJzWPxg
WQWVN5r7kfJIVATYxXzS0Gp0gZNYBhf9o9fHyvSdcpjL8JsDEei+ArzpE2HENUGU
Rb6c1aZ4D9BBOQQj6JSCGPJ/xhnTkcB9dA8lQIBWMwYrZjSPY+aPY9F3RJqzzd1A
bmOLSIrVR7aHv3abbqtqTX4thOWiNB8xOeGCNYR+gzjDaYhCt3DMx82zaOmwG5hV
oBmcrgSRfNjiFNbMEVu33eZFOeaOiRnP1Ub6et1TrtMud295uVG15VE0fLa76Jes
sMNy4eUn6j0L5IG5xwKE7hSnSfvKlmTpsjrvFfHYLgD5r6rleMN94AQcNeCweBXp
9t1xB35qlXjPVoqmsEAe5YMNK2lYa2f3qhA05L/axo61dHlpGdADj3Fr+NkR9t9M
waABD9Ulmq/9ySBp7XmO7AA4ozlT4m3aj8ICLjjElpizqrkQ0PwoIGC8kohn9Eo5
pVKQEDIgs/yoDfQdZhewY7/9rRfiKMn+ZZsTfmP+hjz5Q/vMNmk7+ljnqaQq4alp
gZSsywvGcU4isIRq2oleOQpqri2pEKMjrdOu3UIglyLRBrwY0/sikIAzMZf4asbx
JnwA+jT03IF6Q9CKAX04DpaFKCb1vMlYaq6ZxPJfMkdInpXXDYh9b3ODwUqLxJHd
qtjhRjX8/xwFQw5afuO4GbCKYYVlRLr7V8H9UcUJG+H9htFAYVH3PwJouoe0JuFX
h3WA5/n78xITlaRUaJQl4wcCRQQWkHLhi6lSJ1o2e9ewO4aQ1VmR7rg1Da92VuV4
wC2p9xCbuBUjyCdRLVFfUBRpfp4Zyaqcv3eYzASyyclYaG2Skg9uZu8k1k27s9ek
svLut//Wunuf5nNZuJ8hTLAtMU37cDzI5No8mmbicfpHQnZkoYdSZwq7ncFMMz7h
4N2vuFp3L24gXk04yOY3gKDhXY+LQiWBisLQ08pLvULjkmkU7XhB0M7tLzn35zKm
oIjn6wuqhgvg0ebpZzkw8WGUXf6maoWpgy9AbbHMNdbpHAcHvOqMQDeY0BuImE6p
pFmofA7WnwYoeXLZZuo6D7oeK/RFeYw6gJ4AjmlY1ZgWBTLdPTdNNy1m/lYmgWuN
YfE+ENIvVsE0tLZOr0QkvM8ijbP/cqtgYYZXilOYyy1166+zU9O9N1NMEwzH/Qjf
BwpsE7WSv77VEo0bspl68ZovsW/vCfHh0EeIUG2mk3CdO85JWFa/+5fpi0w3hiHO
IVai0kho18OB1E3rwCPYkqu9Xmq8qUTamweiE2mbn2Fut6lL04pL3Tu+j/UFezqX
x1RLw84STTdXGjTJgLXS5FlW4m10q+NXDpBInkWKdvDr5m0Q7xjJsRvyd6PP30Lq
oOP0B9pYMkba1AJStTp3TrTmH12A5y07w4ej1O8IgHbC5L95SwPJbZL385ZVYRNn
oLsxH/sqS+lbosjc1d9RWFUj4abQcbs9C+CXV7ufsoAHf5+3qjrmg79katNVe9t9
zhwIx0GBBTcOIUMpexSW8E/AzgiVBoRgzfO9+b5yTEKW5lI/GieGvHhdAGbIEpP0
XddVUADPRJigeBVvMpCXF4aHK816Rpw+PvErLSH2+PwFgy/OUK6my/rshuio+/J4
tPddQ8Xn7my2JVPabx6W+dleCgxY6qulsy/X7myBAJXPS+CKRzKL+AXDBA4XSo5R
mqkZRxvcK6ENfVrMCxqux59rt5esKVJD19oplYZomW/4kIw8NVi4M7ElPv+FRfnk
R+tlBwlGSNkekH39DNRjrJyRCwxOVNjFz0KE7Xocy9HHIrIbbRF4/0HdTqGuXvci
NQ9hsVzg5ofdtf7BUdQAy5ykhttPxzwDvx0H3b/amQThwANGFnGSRj5Q/HufGsYx
b9PaVFHSiXBi+k7+YvoFJ0RCCvmrJQCs433Oz9XI3Yn59K6cmb+ANoeXKZZDE8iW
PJBPH1CMAyhNWBS9vqtEh1mzc13nltHMB2Qw2c7ZYkpkJHLWNd7eVpAhwa2qY3Dn
GQedXHgjm5b4JGhdKRKqJkWVKLVDpbJqQ2wBN5KSrolAX+kaHWZEzaY/fB5cSSzo
7S6uAnlioPzBvtwteu2xR3QTzRLJVAwm57RaeMonEZN6AI8+mHAsDQ5MDC00Sov0
mejHSWXj9x+beub3mWdg4/0iPSYcccCLHuA77RBVKF4CCdoHveYKsSfFeIpM6jNF
MBhbZVG2/q4Vykf4L3fbJhavTcHJUWGFehbPYpgPwLNghJO3H5lVV5p7jqmb559/
/AgLgbZIf+8ZzFrlINFqnV6bBQLt4fi0BseMtPjneHdIwrPkC9tmmrSM9lTdTnWC
uxAZ4DkcVbRwJnnLWd7eoRHfOFj+ua6sXi+rs9WK7WMu0AjmsF1uhnfydORAaHE4
ERAjpEzrXJEpPGfcoxBFlQzYiTKaDS3WUFC6VyIpAk7FJ7FHPwGWl9B9qcnM/whO
pGxk+2uP9pCvMThHut2E4QSF6SWBKkTH70br+ZROaXea9dpujZL9FMBcJWAj+xca
VgXlgauNj5jxSjgi3kebC7q7+4yF36O2M/eckFhU7F0WPyYSDUF9T+c0rmzyEy5U
NM/54yfdEbIYn1oPBluoCLSkepzF8/s/Mqklm40jjjNIDRexVMROotGYKcNbQJAb
BWWO3hjgR9314UNBWoeCN6AAHn3WloqTHzeEcSPKcacTTP+mFqq+uqyo7z3KRFmp
+Akz8GGbT8dzq5WNY6B1kdxwoNQarByMnaClga9h3GHHCBWaBwHwS4PJj1Cjyjvn
NugxAgbHLW+FXUq97nzBdF13lHtfoNfKPmeAPQM4xtvHZIc/83j6gX4ta7DCoqa7
Y22Pco3HqFll3nGHtXfqxUdOnoeorHd8MVa+DSvHCaWNjjcbQ63yOib9PTnJueGa
9YT4MEheZ7S4V5PaM/ghPV5D6Ak0TkylY+jznh9GMO9R3uMyY7YVnjQ0W9NkLtPz
hrpaC47hSZJDYS9m2hMRPIp7dNMRqpDNUzM2BDVNb/94+xRBbHg1+crUqTzXl6Wr
0AMN3frzExAUP4Q4/t892PTQWqQBL9N2/ZAnH1h3FH2IIptmcRsShXdM8MRTJzw1
EEWrYonL8hUEU487Ny0Q4qGo4OoS7MoPzk4geNQS9kvv+YZR1dyTEMXbWRthEsrE
bAVDxyqI1rnQCwP/ufqFHIMJCY7W5rqirq8U8EC2uJter2lwnebPnh0bKH9WmF0B
2Os3ijPPyQO5nzcdPpdwzVWFbNrbDcvVTbogA+SSkBnyW+ea6/k9xzXT+z2MJeq1
ZayKWkgJaaFpdDlknOuja84dBT23WvtHwVXFHSrlDL/MRKsUrtGWF05j4J9Q+i3D
1C/K1dumqBvIanfYquCszVzFyXbDrw1fgDwkFGofdZmzUJp8UVwUAMmp1ENWT2NT
R2WbFmxsR2Aw0BatK81sAxszcm9XbkzO+21Eljfu3MzO9wKDeKtytJ9d9gmgND/Z
olIAHNLLyXtZAk9bo1/jcLQyaS8Rvrns5vhOBIFWV7ZU3QMZ3wXp6ssOstpoQzJm
bvZNx79DUpx9dez3aTE85MmCNaKRaAqzO9F1L6lnzx26RGIMORf39OTS9BdNFmmG
dkW3q6MGQZl3zj+lZDuDj+YOujHo5mGIYyXnaTsu6A+gpfPhSGljXrcA84MpUzzi
UsCQfVEpRS9X+235Pg7M81vtLOjjtTUxos86j+GNQ5rw2lw55ld/wBnSlraA9Cty
jZvOPJSHe3xWSAwtsEZvzTe6bBxlnmwOOcxHGoF+kd9GFcfSUhu8EqpxW9zb3brq
L9Gidsa6tyTYur1Eu9xd0i2cgtzgowd/ENue+H8hu423ksSSgygypfCpBqw7cyK0
NirgfKDUs6fsQ7y9SPwPy5erZYAIrAp5/qdeyY+jwS6+JWP6DxwqklAf+SGfsXnq
dpSF+0YDpyVkXGzxCNQBIWMvRNanVAjiM25GJ+g03a0Cl1Wb5hJcZUB6oR5picDt
YLtLjRcq11Q7Q5M3TGsyUcsMxEDkPSwNX3zRMTIKM+HtFEJa5XOHBwCdjJtL0eqA
Ol9JUSGSpZzmY15u2RssCcztppXSaN/kTHXG3wss+NjcgUAzFfuCui80YdoEjkCg
Insx2Nxvd7SNtnx3wct3IGk0AFDGkG1f3h5eSVVUyiigJUbXehbXA49KTRNuiDK0
zLYSave6ZLJV7s/+MA3I8O5ThmEm4VeFiwQTU5yPj2i08/b4CGaqHPxD7mjBIpDt
g9g4mhFrHBCiLPgs2t8GQzMSQCi7ztn2DbwlhigLu1nMkGxSri3fvK55LNmD46ja
s9j2XTHL7lfzvwlqTpxpK9MvQN4mND/VCi06QVhqfIP2zpSqtnvSNdLzSafCyeut
SHZKCQIobGoFeIVAPM4ujzauW95RAcmb6LW3rBKVbnU/Fzk/zvHNWMC1f/s5Ntep
IHWlOqjwargEGZlO1pHzwRL2lzH8kWhJKesnZHdJ/eeeidybye48QxDn0CQZ4inh
XGtZO76rHNZ4/FZnFinlFPupriB91imKFG+IaB2BCOPFGMb+dh+1T1vFm+kFoAo0
9m/zgyn7LO/j+TR+v6oi7AXguYGdtF6MxrpZjd+DI6KYOitSkp8uZNz6koe72p/n
kh2V+t49iFY4Szj+zOcHeE1Nrdz1z2Amgge8xu4u3Ufb5Qqiw89ixTIBma34nLC2
K1KpIAK34Eeh4WZA7rqzg4b6oesWv9GXGsiDcIA11rxYuv0QPWb0YXBDep54kZhd
kPvn4a7NPpwqDRWlWj82ii/a2odHM2FnFH7q9lYZKOxY01J0+H1YQxnY5Klsu5Nc
ZsqqvF0tmOkiC8Hp14BJVAhLkA7oVOkajkK7S1RKtgihhqLDbLAI5pKijKtLPSBD
sevtJszCm0K7POHseG4CLnIowHQ/PLuARTQHbqeUZKsRH75v9Elm4R0rykVEGKEx
7ArukZvPDSGCPUIIoJ2xn2k8LyPvGsQYVxZBk65swysjnLuiD9K0fIXeVEHNvRXb
Aa3E5uRy1Q8cvEQTAR3GrJtlhNhH406BJXde21/iF/nVb9tETo2WouTyK4VSUghC
j7FHzaeY3M7kWg4Rn2Xf0M+n5blnxVrfbnyovmAQSy7s2O310BeRvROHomwej2gN
IbCGU9eCsOzQC8wiphKI82t6Sq95II9m82MrBK2unNLh0+2r4lMT4JTMAgyH9Wo/
o2OrRn7z9qZcYZMspSrmlb6Dlq/KjGuKQLVHhIpJoL/hBGNahyuH39eEz2FgQBny
LERtuHZr7wvJMPKdfdZXqJnwI0tPmryO5v1WfqzBtdpjUxrkJgmxS7/+rRBcurZ0
jgXyQ5ZuqKdXK8hoJqWvPswz1FOGPMH4a+4Wj0G1uhysvddQVbCKlDgo1gCeuNRQ
39nMWsvXjqkovqAE/vStP2xiqgOrdZsCZgOP1Ru7FmFppsozpVF7JCrUrFlrDX4e
fxbK10LI7XTOyzTPZWv0Ei3/kqkC6JHbW7snD+JwkEuWY8gNlzyPSweLXNf8R6w8
hLEnud2/WSRophTbvi+xnpiV2grUGPHLUAG9s0XPl9dPRTXYEKfkDMrQhFjR7CpW
v2WIntgrpclTgd9j2R3Q/nvzp/QUY2lIj2OY6TlqmkeXmcp3FNH/T6jMyRCxjUM9
DwXfaU9XgRf5Cbyhzsho8qVxWyte2itHcFjiPHxh7Wp/U3Ie08EHOY2r/MHqiYwK
NzUWPtVWZlvXxK+J/RoHWTS/9i/k8hVjuooEAbuOT3OB0HTHMRPCNfTGjXPRx4fu
IAhMPzLe7OhP7yhRMdIdkRF+iG/xSyaJpzdWisgHAYfjLXFvc8MRNr1XIFuRaGOQ
tGLU0AudtgM0+HkiOmw2if68Ap3Vq8r73/ElTowUDoF9sPcDZaiYuK5iGe+oEpWd
Za1sa3AHoQ0SJM0ieAwGQttG84j8Th4lWmSodYBbF5ajz6YmxqlPAPeegxmv6wDM
2EHTmpCRmMkQhyszbGtmtktbc7h3pX4cC5JC9+QIkE2d2X2w20tjlCDpGY7ckSfz
AmbARQgraw1eo4SI+r2qRE/tKo9fRzIjmeSUFYv4jMk94622jw4r71MNWEhGFJrR
BedUatLuib3J2npkot2q55pjL3cGHOm53NyURy78kMp4cb38uZ6eYMD2I5vJwAG5
uTgTs9au5DT+8uGZc2dXrnLP4LGmbZ/nEhZrh1cUmNJsgExDlv/jNpCenQ5fnXvv
8jSNHkhDHwXXPb8AaK+tn3EX6QU5lGN5USZhIc0tFg3MXQcuPL6W3gNiy7XKJc+S
Yanwylq6kVPirckqYLSwcVUfhuvG8PWgkHzVVfHozxFKOSpHOUShT6Gl53M/AYqM
NRpti+yj40fvS18fVuuzq4LUxxFnyEQDK/KcoKbs1ktnUwjrX9sgecsrWJeThpGV
irr5Jg++HmFn8TbjxIx1hIJl1maxes4sOf1ym38ORjGE6U7vXz5gnMZrv9gUnnng
1jGzZm3rnwRHUCbE20IqrfA6WC4oyCZc671KIvWJpyNwPJUKLOvx9eVHIuA+gVpz
AWJBKJvZZGX6TQD34+RI12M+ZQZGgB59WRWdVqciBwQDyMAFjX470q+fgyvPn0uZ
6TFe9L3Rdq/q3MUQ1Zbyy+bkrLiqBh+4PIsVCTFmiU4HIm5B4VWH+l8mfIfKaK3x
bapOBFBQUUlqjJdHXtG/dQWtMU62YOM0EESjearRIxEx9VyIlBduOYko1bP10Qs1
SX4hDsEbVJ/kHlLQQlqtwIt91ADxhEHPLpaMC6/aYSbqmRfKqfoWMemvmV+hKC+k
HpwwpuEExLx009yIevCR61ttugQ8T5n94wXoj4yPL6+bReyBXXGzxC8xemcD4csY
UTXLrckBmmNHt7DIomvbAraLmn8UmdlLH7B0Thut6ilzMMekBnZjIc4aY3u2tv5a
CxiV9gzjb4gi69w1pvBscLahwflIrPtbG5mEKJc91A5nVAyVE590GWI1XuJlNsjJ
fsL7fOLH2z0kDYDOnm2ROI1OjiDzGhRW0aC98NCQrvNJU2EXqXNbn6Op4VGlTSVd
0rvTXJi4xo9BLWhCxLAKfozgSp8ZMP2h/jrt9qxf3PyzhOJ9yh33mqxa1xT7LElN
z4BBY2e7GIMkgFF/XRU7j7IP5st6jp3uz09jhg+8cFR/D9yaOAHWCCuS8n9FxnGL
UkIPsX3Uv7kkOeTb4XrYm++xbRqS1+ujuloS9K22DdVIn6DmH0WijYnZB0xT2FGv
uGLfAuPzs2JOS1fOC1K7hkPFepOBnxbv0UKe0GHq0VwotEYSaOip8ILBkBM8lNij
4QjJRE4HeQdDGP9xuMoOSOtDuRcTYVk6TGMH1vrMLJDQV6k3HkzO9n1MjufD2a4t
+LozCk1WJWm4k58Wv2uHo7/qQymQfTGaqaqvdAVsxurCw1WFp2MGlQx7AXy5gQqa
4YW3P4BKbNqWJq4oscQ9cffOASGdzlB9k3fMm+pbTmR/RjBd0/rDgzONho+uqKhA
N4c4oKuLq/CxewT+2phDS2udD5r3ExS3+yEAaue6xD0F0AJCh6yek2pQ+Nzg8qTF
z/e+vueP7gTS8FeE3J830XBGkA1fC+0nVjgSRxzt2GSUtemJSFv1sHvDphvPHuot
zJhP462Nr9rdwTkoGX49B/dCHGu1QDIlT/GhdDqLgFEPypAz1kbJohxiE6l0oilj
usLhbwUIgaynSc5JsTtUL1V5ZSHZIdGDXKRZAehOkFF8JcBfEzBoEaUcOOY0Gq0o
8FDoQQRDahr2Q/JaTAcwvTIh+aeK4WPmrse+Iqr8rHzaYal68zLMSVFI/nKE42oX
U2TfDSgHfCoW+1Xt8eNArl6RAxXM6x/LCCP+FPTtEz9WdpIaviwjo9F8T2gXJjz9
jKNXoonbPwRanJN/tRIwsoerRsIVoNyhKjDuTps5chawun5W0Z4PuPKelF7f4aO2
Jazn9sNJ2NNM5ud07XvrJK9JuDG7/AoY3oEtKC8IUqGvba7+GQ3xPlp2ikMSfRPe
mzlNTT1yeJyNcH/htyvjdvNRJprEG7A4UeGQQCPMlsuHkCjwV2Yb4/+UDa4LraBw
Vak+oZBncQ8Ul6UUWt6wUxkp3Gu1ew7H075VaQN4zWEN3jMVPLASOGW5qHyhgqiU
W+iuUNSR5nDsmnKb5wqEExQDWuBIEwU5Elgfo9qaJ1ROxV4k5wv5IQkHObPoNRSy
QC0HTPKSUTqM49eekbChLzscaDOJinYRy3LchGrQSk9jmXiSx3CHbDU+jct2ThvZ
VQ9bJnH9n94dpQNvv7d365lvE8cHKvoGbuEo3mCK4HK8oukOHzWxdPAPKqB+kle0
omYM0VJ4vGG0OP86A7pR7L3fIohQjIMH8N0U845xVD177+/jXgGm4nVsxfZ9bqHp
+JcK5blw+RpziHcii2A6+vpyOuRLZEcxDYYO7gUirsmvS6ZYJoiOCQUpHfLouFjP
GtfPQRqb+fRcoK6SLncMEutzMKM/0rxZoN6/vmOtx/7pTvBCWlW0afkzGKIk9ZQM
KsPLk0SP496vSt+wwJWyCcoxWWjYyKfuYKbwy+KS5NWgbEcwfdyrzsZ8eEWPcb7h
JfJ+tv1m6roISXvFOnXDFx3iCzkS8NUDqMva0NVV2XUGNtjz2qp9n1Z0Ktwugtg3
SDfO3GFm0+KtENvu0XmNgUp8YfKdVuCJhafdSx9Vuf0mpfdRtk0WcNNzdCHQ48hT
XTRuY1qDr5fo08upLd91FUeggClDXBSaX7w+RsYhqwTJla7HWyrDnryzRCPQjVrP
6CFhYUXDhk43yEvDnQ6TAff/smZDPoI9vAaEDXD+JIpBTkSL31JruTZ50Fngv2Ls
KZ4LEnybgNcS/nEvCU2M/DPns6AQiKhEJR7aItKScHBDRmIngiK6QD8hov7Vb9wc
sag+jC2fkR5A7GM0/OKE3y/o1OEtUDKuux0PdwWjc68TT3IsOHxvOsX62BBJ+ayQ
NTz4p3f8AQmk0virHTDyA/H++s40maVID6OAWBeysVPBlT6UChtHfURoY1L9b/Xz
u84kwjiJ76RAhh9E8DyeABfq4+DPMGjVWGQTBfXkkIKhBC+5TXDDP1RCHFrkshKy
UZ3BYhr8L7j/E80fQgtr6DT+XPAC5aXfR6nyZhmkzudGiG/Ya1EAHlQXs+cn6sUt
KAP8eM4kb16Wucjq+lQ8iT1jvXE0/pKJxxfA5ZJOJ4ugLVyCUk1ch7/AwjpXrq5c
2vWlJAqgCiUXEpxO2xQWAYEYLd3S5pVgdF54UcR9vpxakkiPPZccYFjmyim1lVG0
xaD1azUHhJ2odd/YaFTQ8wZdge6Gw8nqkdADgTT4u2KfOFynzppoIvDd5RewRB+j
hiy/yFeiAMqYPhg5XO8/9SHoyD7/1fsiFv16VjFCKtq2K2a5g4spjTEKOCLR3bjw
qJz/bOrs2UdcTY0qvLdTMzUkHRmmn0+8VCKRYzUcN6+loFqOxzAfNIcniwHLM3gS
+ESV6uTtnR1mXP7qs5wFbaqC3W01zgR69NY/qvmOhpgbA/ysW6jWTGjmyPsqToeU
m/Eyb06eRBANsR7zVFz9c+vt8jRlxnw77D77ZtuMjujkZowbOwJCU4Mma2WGAkA7
g/oMNAbzcSapJJeKvMwW967c3l09J698OqoW4b9+4Uv1n0Gp4VZynFS7dWu03Idi
1TckkMa5r86KNQvOsONqzL7wZgRYE8B3R88XfYMhXiWgDh/BP3wmFxvRWa9zHVH1
MG3d6UePzXOSmLxcKLim1l4asMyz2Lw48whJ1Bd8viG+Zyxiwx+8TSv5kI+jmVdj
RRyllxvE7zryGx1q0kcGAh3OwBk+XX7RjTqYXphn0CRs0aKgONCFVKCLVcy9Y16c
wFBK/2/osCl3MW/ZAbGhnf1oa+mL4N0XO0DXonsBUyNqXDsmHyDYYYRZtFwa6pvL
uilzDKJi4rmsCCxwjUV/c6gHLG3Y8fBf72uBilSn9Mw4UoYnqFQw6SNnBB+iV6vc
p4236umrtAL+pO7LfHvn6Fc6WxPpjXJ3AcnidYT3R/0bSd9Eq+2g/VfhO/1houg3
gCvwgcz4FPUnM/8bCTpZXu3mwKQb2uxZl5JOoCJh69X302Iwz5ZKrlZDBASwCHnM
+69h2mjBtHej/hy+R3dApbyxx+FMHpur86/EqvAnQByh9pY7xEMgIEyAUJNy74bB
ZuYtP19d65TYjpBHWBZMAdnr84H4WKfeHfcbm4ky570j54A/2G+UPCmigCSO4dg+
T8EJB6t+uWGyCPJPPCBFLYBAcV/2cFJZXJJfW7q7KdAgdeYQ3ogAqyaQfMESEcQp
v+aodNYNg567TUUs7bHZtxxJ8a/RTFRqEBFhBEtwC/6ZlGIFHv6JDVudN9xGbeBN
kE7AEq9eVU/uDkeWHYX5Nt8cMXUlArOg/i1FVNr0t1xuqEw9Py+yH109K9YC7wFA
q2W/zMjM5nMcbV6X3xOCEsfOh/dWW36C+LBS8tPjBpBBxr3A9K/vuJBPpX9YOIvE
mthx21cMQL5EBjQ8/EaExerltPJWrnf7m5jMX/kc1DjZq9E3D4g12paGzeyjWqSC
xaO9jmWBPlRPx2jj8JO4SSwTyrf6qCDD6swqsi5B0pj+vQx83euGZ8Vbq1ZmAvIj
UMMIyndTlyfM2j59qtmSeqFFmEXPU5eevdZJgY7mDEIgGvqDwfTKR8x4lKQUmtvB
6RZsGDSEfY9IUBbm374EMvFPw2jEB4gGKyq5hrytsod05rPTNk0wz8guc0R3Lr39
ondQDZk+feoY5JVPzehOkit2fMoxw5AawaPtV4JzgAn+QLcteAnu+VeemAemzz5y
KHZYsuujQjQTqdWsBuNG5g5l503myAbnVyKU76tHJNmsKlH3E//rxZirjhw+NTRy
Bm9yAsbzMmkilXvk/bRVbg+CJ0zfdBVySOmBs9/8JymP/380FoudzHH3tQo4yTlb
iXdsAmE/Ep6zWlRJ83TxumJANbsMVtLVF/jP409yXaB6ZNELAqEqj07aNIgAvfqj
Zmpx4bYSPdpkMsBOOOEOrfMHtyq8FTBx8szw1B+YQB2fRP7tiyoMRpw0gpf3MeRW
wHWtvPtX0PhddOhQPEMVvyj1h/wA9KCgtmlIFGU40acYEQ83AZErlHCeP6sY+ECc
SghShA3oeitRnaP+NTgTXKr8eoRoKqXBoyKj2QEQ6AxvSX935BRL/BxiOq76Th0Y
QhyQwzuS5QbsqSCF0aIKHvwbYHlCRefCsSQWcAYA25Sox73ccWSBrexHX0EdekXV
jZF+vTLOLGDjjYCSXFW7uh8CgbL07q88D+hAeHDBnZHVE/gHVmHl/Yh51x9/lA2d
EqcnodRjuZ/rYs5MJibPxdLHvnww/Rudp0dJz1597KexRViAK32WM7wuKHxK9+Xh
4Bkaw4/J54cSdrdpGCjayixax7LLaJQ59P+tE6onMekPZ1m6UnjN/OS3YcGfu5Rt
9JADXA4Ruejs3vgmvtVWSkO6h+urEVhNUZzITIbOx5YXBuFm5HUGMA9gQBpNaqWW
RbtHiuGdnncNZzPAI7HAXlqD+neoJ2zuJpgnvenBTOmBkx2rJWzgeapKg+4q/Sjf
SuXQ7CBrHuJ8epQoORM4/bSLZxtsDN9VvIKTVP5ZeogqqyG+kKK+CqPyLTYt91ak
/ETM6KnrHPvVigPesvkVgwHknNIlM1uERGD+S1cEvQ/2ksmZPudWO3zyRZ5qW6sD
mJc6KZ4xOPGK0uXufE6oXAhQynabbXzIRoTJ2UZAQITmiGsoeVoa/IhiKW14gAAR
sVVXnE33uOjp2ewhEfd45L1GS+caSAuIXlaKEoILvJGa2HSW+pcfaF82peSXVwIq
6FCib9s9PLZStKSfXg5WkCHgmtMuSk3p+PkNMTfNKk2E6PdfDyE5ExDIkQFUQ9qP
dY/Dm7Kgh+olb1OblRhBfzR20Ovj21nPCHnuvsM6D8IMwa4i0yIlTwJKEVHK+A4H
Yus3aqJ8yLVAuoNqf4VrjU4eYVhOE36X598AdBZn6B4tV1vdgdo6Lmdl1F2rmyRj
Z62fxJPhunZFp3dkxHlag+XkphsZsM/FqCASrZuXQXrRZC1Is3JdDQPvzurjetjf
hHP19aNS24Wo8rbRpKBRrF7bprIsiCxGWOUneqcYKWl3LB4vRTCjGTxmEj0WZmQb
0uQ+LY8ShRHsEM+wPgTxkvmWIbw683awieEJc7RtMHEliwXuWw0omxA+R5grgUJm
ASznl1Yd5qs2/lggiky2dnnREHRtIIA0e2/W8JpJZtbQUP97SalgBElgZ6y45oxD
CdIbL0bJJozVjikyUHC0CxOOmyj2M7rD2X1ZStD63ZxyWMqwXjGHFRxh7QLsyOVF
0FDuEBGZsl3jYUXNAT+RtbLnIMaeUa/tZ5Q4qcv3sNhPFgERmpkmwg7xtxL34y4J
Yl1nicOtj4Zn8iQXyIzo3jhCUWcc6wBRT0Psl8rXb39TifKHX8y1qup7WzjjLxSK
0KdwJp1f3F25h129icnlyBJy1JhcNSaEGdBCJlt93mXDAXHqkOfeTjYWeZ8vcSil
GZanYCn5k8cFVfBLMflrGHxBUBvapPZNebjPs7Tfm8fQgs7HUDgAjMyaeCGZsXCO
6tL788yDtvJFUTjk/x4NBAoDfmBKzzUSg6PxiDk9+f8inQ4rWaho1h0IgqTnHELS
kngYdom/aUibWrlkH7uoI77MpuHf7tmCD7xU60oeA6AzSmCe1uGXB9rumaMoTi0C
UEZTXfHk5QwpyM19q2e9hElxthbWXx8u6BfgWFniNSI/8vPLshA94s1JhydVDXfU
EcjWPtEQFBDEx/q3VgUWENupXKXJnsHNRW2EDpECvAMmvkeUw93DUk//j0U2BOKh
g2vmGiP+EhxtXtK6K+de9oM0P0cH4vlMVSBkqXgLh0w9zOPvpMkIyf1KtklQRpEL
QVKwW3GGvTsfGdcBGBLKvBLNqpLK4+1510tKSVOwlJBWoi7A6UEAXC0jvhtYI1RC
oaK/pmwb/1YSiALRzh9AhSYW6Bfl+mnAWXo26gSThhprRVk2CVaPZAkmxFEUV5eR
yWAR1T9kyskQ9cgLtIf0fSzMyUnukV3erWVsjcEGKJbIYA70WBUu/oODeFV/FIN3
Bf4F4c4HO8Vx6Dfei6rbv8XfjoLAzhBl7Zgv6H3DTE+wgN4B9bcpa0I+m6y8OGIo
K0GMjCpJpNuS+Fq2Oh1nWIcWRux9jMR2txId46Kl5dukKQBKXIoYxATU6sZxLfD2
8GpJwtYtbdr+GHev0NxZbozIqzzfYRXxIDngVIftFG6ys0EWCjfi1gaF/hKgAq/4
BXBPWcznedB8aPB9XVKVNd7Zwr/s6Rbd/WLBeWIK224ZAgtRagJkrIURHeKZf1mo
S6h/iWh6WCzoH+Vx5CsnJfeTy2OD6SW7hc+KQOyTR/ZYTXXLN7j0ftV1hDiUar46
Ktgru9oYEO0xT/fI+Ak+Mlql47ohhk2/j7IDpq8OixNZ9DUea600Y4yPV/gvwmIr
6/TY9ey0U00Cc+V+ne1YqAPF3eEfog86VBn0KS/2OZPYMmp63pGEP4BkTmtG1Hig
neAjU9+H/u/nUFhbNgHMMNsXd/vEs0TWLVFwQxsPVP/5+nKF5t47TX1Q704eHAz9
qBlAPSqR8QePzjwrkQjxuvfN31XTFmtTcLYPsGvv+tNYXiThD3nmULhP7plXFDVC
g+1M+iiqupH/zDx556uQ96AFZZ7jrV8ooyFdknYuL3ZKf+8GNuHov7DAcwN6PJp/
kaZYbZ167xT9ULe6HkaGPHZwUMC9fv5B4qAaYTck0CpEsitHxos0i3hI47YxpKeD
cTvrVBxoAChSiL2jGjYiAnIy6kLJjdYQsP8pz481a7/2odnYg8dfgMgFM3LZZsLD
dOwo60PBpJUDJAKWP47pOduN3QGsBYGYHdXhUvMRkJIkZkAPH+Hh7dfJd0KaItB+
oy/PNvmOqsqS4oVS0iKRwvqdRtF2Zb1nXB8s8ts0STXpya1atnSnKzPm0TpSDJnB
SJ1+DHxbHyPfpkNflmop38SM7fuERIhZA7Ra13FHWha6iBkba+3VNoAJ840d6aBH
wzAYzP/ZLlzSjGWHzpqlDyb3xAowY1JLOjArdU0ShhhW9tZR7jP4QSYyB6EtFLaR
RbnbU1b0Js2eiBSMgjoRMWvpLlNREBsAHu7n/tC97x2rC5l1hZ7UfULzc7bHhLco
QHAuVOsEpYJfMswzI8MRuiEk3HnxTyhgWQPAJInMm0OVKFwTtZMoa1v+fD8P5CCW
aaj7+gf95kqhDv+/QzB+rHG000qNH0vw/rjyCchIF+HcEBBynyU1zAyUBfQNiKle
XECgcLTxMHM7kKLiDqRKhc/bwgAyxLL7htp6wPfpEzHX7ZLqYKrJ2pYHvYOIHZi1
b9B4LD3hqQOFSKHh/evd1X7o+y+SvLduDxgEWfxkQISjty7fNT3QQkFQLnFG2ae4
l9iMLnaXeYxv326ijRPxEq2wB9j49Ll96KXo1L1zZNEQyxoWibZ7b3A/V76Vbre/
qhvCwyAExbckFO4R5JDumM/iBRl7MNQDXSVnmcItpIO9CIboEkHr3IOUaRgu0ZzP
NGbyWwib5AWsf5WjZydsEH2J2EQImvUJ838tskKO3QxAixRXPWH4FXePgLizIom/
kcmFmBSNe4FIPd15mWVq5G/G0zIrZ71XSCVIapQ9DSWMirN/4SIh3+dyvbh7pZG0
56XriMfvj0GxpnhdsPsz0fDuyxcEsWjz2a0/HBNDlhNDkBVB97KC03Q4wxVgjJO9
s/paL6x0qpQwXYRgExIiMmZv3V6a3CRe0dq7z5xbuUy9IiiCzZ3g2PXGmqGaTXFr
ey5rka95ahJdm3S3f57ltgccZbitftqECvgb10fT2+ta/hrXyRZ50JcGR1BQc7XB
gjXn4/WgMbQRMs+Fk9dNuB+IAqk4XdpOc/kTc1iktttuYwuhCvtF7pjEYbfzMUvG
zxCB5cdq3dMBeOUxgMT0GbG61B0UPeW0m9g6nOgv5sAz1yYLC0NDFIvSFT2nG7Zj
4/4JigYMaFrFLAuQlwtSb47VzGAxL+9FmqU8GT/Kkhwbw/hgWem7OKU46qD29lta
YH5zd/dur4oRUSV3LDxrujMD0Roc+5ci9nSH9YepVPRy3V65eSFByQdFSRB8wSmI
+OliYQlUxznYzLb3FxzOhaDxDIK0Tp0Gl/je1yPRVKjMGdX4wxdmrkIfxWaFSWxY
JFVcjC1APB7pCksanQ+xQ8enXmTbXWMBIRklilRHCdu2lflEU9ZaHaIN6FCki4Dk
JKsO+ABVRGBF1pPEdEMs7RCrsFoAN08+QFy48edM3kJpsANG7VGqx++xDs3+I8V6
hkXwvEIigYt/m7HooCJ4TZiSgWemyurxq5OHHpGPWFx0QVi90oZ6kdpLlDqw71UD
Bu1MJ2l9YgfvP7LuLWJB45fVKFykCZSzdNB4Ko2BQnDgnPJ3bwXUYxcW1auSLzvi
RgRW9FByyZ9Dyilki7E0SjvmZDYoWd+GB862j4lKR4bwjQu6WDrRbIIi1BwhhRgu
O+bt8j1otCp1BIqxszCrGaCXXLEbA1Jp6eL3UQfc6CvE/+2sj2qN519hReP51v0E
6aNGsEi4FpinNFnwTUO/UtFxdG82qAT44gEsFWVjZAHEIcIheRzg+ruGbqYmWkQO
Bef0LBCoVJfgSceHoEczu7YYbPLSqM3R+M7IDbYke4YFglHeyg2dtI8JDH3d4vai
G31/2GiREPoot4Mt4Y6U8JkgLdaiRaYXzoFL35K+Kqvf42VUiBpPt5QOSY3o7jEJ
U28yd79uLZFNdfrIsGK1QDcEHiJzhZDYFUrzPxXObv15tI4pI2PmDBe+LdrDhDj9
/T/6N3Ldc9BiziB/fxN3PCytDFlPZ9bDRFAXOrecNs5gwz+fGtAEWAhjX8/8VUj/
F2gAvD0BHluZxKr66Hx6ZwLFfMhaBqVm0YxFI6m8O1i8ZeMoZSv8jy2iXbTr/lH0
JvTRNOAO93Msn1B0ipAdDYTE21FiLj57cmTB3RBEM6EGHAOtaMTJVij6OYoOfq4+
GakPffaO9qlqYvCG7YICj82BImTEQNc+MzA0UwTzgtqZKF3MMjz4LEwOvC1Fw82m
7z1cd53sYyoJ3kOI/036TkoS0A6sBxVhU9TXgdYZrJZaPUiUrs/PEuivcb/zoI/r
4trvk5vZeTDvgb6oSGYsjZdv0AGYNLOz1bZ6JwDSPqv5r2B7lkU8X97PRo+FKGE2
brlFl/G+2PICAjkynpSI76DlEFaor7cVsHK2EG2Z8iWnaKniInzJnMJSeq+5QdML
aI4yT728TAec97RmmGF34SgmHeGSu2z64lcH0+/I9cgULW+PFUYx2+Edr7u9KSOW
uWwB/bgaRdxNNo16BvdOmSODjs7fPTIuR75BRAnqtWRFm3HRcgck5ihEK1iVP6TN
PHNEjyRPJ2tsDxEvqlmsnWFs2F1UcT1qACdJ8xWMBewxMwBd9hdJaY0lruQghklM
zs1NV1gRNBTSjbC0ssaoRg2BTlCf0NiOppL1rUQb9pTGoJkvtasE47HyPyaKs/mX
Cj/Q6v9BVU1uID/y3fFd70X5QrCGM0iauUIvBD7CL2SsXrAAerSnZ/Y5/owR9ltS
7/mmoaIaDDW1h2Hv/sQ3ohQ8H7ADlirlMs5Ml6mBNkRMsjvHVEu3OPpNncTSSHJI
X6RE11qCcrcuo7acgqn4DApCsTEkS+Ns40fpws8wSeg/LN0/1+3bmPgOtudpen3Y
Bnq9K4CSqRi5gk58+dAuONFU783KJq7KNmmn3Cqi04Fy3BtcqW8wBMPdQccTzLTw
ZfGutHdEucUmApzwUMvi0lWrNn9Gwa4HG+s92EfVr4Ixmg+Ve+bxan6ukX22UdSp
5JcxaDsTodNJslV/Mxjp9xLbV//3RrFuq/YymDo+mCmuyCOVwRboSa7IKhHjM2ms
VeovVDqvxOfnhzLCqzkawBG9tvj/aTPHZRgSGK1bPULcR3gpaye3VFguAn5zeb3y
jYDKXKhE5FEA6oW9/sbnUgjLVIEOXryc+q3SKh0jDzUy8dQH/0UU+3lL1wXcrJmk
M+fsYbYm232w85yflRlV6oaLH0PE6Xxp0CwE3bvfXYzdWdOd5pIUcd/tFVqYYMVD
Gl/OgdURgYkyHUkvO75TJ/FJellM3LJT3QQ9z/nIEkoLszam0DwPDfPyk6MkIMoz
mNUBG3lOQQWd958G6lHY/vu3Nu6Y1GMe24gYx4zJFzXvb0xm/NGCYuybqDqCHgX1
iTv76erJow6d30QGNWPEL4lRN6sgxgJGit09/MF0r7DvBu8W9HFCtPF8LygutiM/
30qYwcjjcEMeTAMYemPuTeoobVj9JHdBnhu0gFejPVgBmwPSiQH8jUAstx4c1GLZ
A8/Gvh4taRzWc2eBIRMCd5fuTGCqcIbqdcSmbB0uaPyaZ9zebwNcontTWVWk3mAO
BUlxThMgTBKymBOeiC8xIvsphsVltjPHgw06oPK55rH/4qbtaMuW3hEpL53tAXSO
THZ/umkhcjnaQ/SWkllaD2HfLUEtGNrynQm4QgiuF+VIwXujQFFhaJuMC0kSPUw+
FU6AMpNBWKhGYBSfYyTKPt7Dv8rtKvAd93dEf0Ks5bx4iOexteVG+aj3mOd5h3bs
/VtEZh3BwsyNd7VgCqXZCvqXBcgzBD4kRKr7ahQIiTS+krfgcTqTHlT332/oX2G7
EwQ0CFz9fSObzuoM2Gkrg6/m+bSnost/yyP90LO0To7KWiR6vr39rZGBvJ2Z8m+H
GJcGMacbNPtZzM9e1iyCkUQqStz1dbuq9We5twpqgoL6AfEDADkyzOVVClFdciM6
Yz56Dz7v+fr1MCLFy7aJQWG2iFMH+A1EUa6pNthpNEt7hQNNS3tKisjb5aOEhk4X
r9sm/qGwlkOaEz38QRFCoTWdPm6yNPoVALqb1Iqf7o44mR6tM2OEyAtr2ukxrF7K
A40T7CbMi9uGtCX9cuvPpEHNiD1XoWJzojnM0Gcn4SkEoGgfgpbE+b+PGqxk8bEn
J2Kqc19NguoRfmrLUKFI9W6FcEiv04HRwRCT5Y5kFQ080/Knu0Mr4Ftw/A8hLNIv
hevCtuExmIY1ipM7Uupd8fBAek5hp9NPOB2TC5iIMBRAVyjeL8Eb5Kh5iNlyVzur
lX+NigNjiBmEgRmXmfjQfwACwijBKQTfEYtcXqVrPH8jhP+KO8p8amXBEcehwpux
g8TUETFmmVTZIPdyCb1c+YptpkZt9vwWJhwWnz/CcGC5Nti7R9RjGDc/JQiOuJPx
axUyMaByoNDr1Mw7BjcDmR/msRy99bLq9FJkhK2CFjEA2wqdDAWR/9nGWYIJQg5m
wGLtKa4sgWFZ0/9Fk9YHzP6MgwjNvmRtjEYQQ+xEkM3jFO8zI0rfPVjZqdH+mRxR
WXA9p06loJshzOX0yGQyiYvB9W66bmyJpFNgXN6p+U9JaYGCebF8bolY9UlTth4g
ifI2s/7rNUcXhW7/oH2lvkh31pyO1dB5JojoDSWKybCPPw4Qb1HQhEC/48Ntza7e
b5mWte8Kb6ynqHQwmAM+GUNvo7ebZSeTNSmDeiFHNfGhMh93ab4igPtYtw7z4V67
5NkV3UB+78P5GekhEvf8c88JHjsDYaH5Eok3b/L6no5oIfsh/QqJKLZTsu9BBLHb
dnjXpC6h7qqtNDzc8fnEXa2sPDj1F/ccyR77MqQbs+IXnXbhmAzlPsFl/a/wZTbv
uDOZfDjNKrDdOMCjvnXR2sdMpGld243yjG+9rvvBmytovEczodZZd46mZSjdL4Xl
wjwg1Tto9rN7AGaml3AkcmctB0zmfI3jdiOh2laC+YGtRgfp2ImM+KWDSHGM0cJt
xtih2vGW6b+y8PoHzhrc9aAQPmUUemCIrDu99cdmXBavSvkhQ+BdjlalMIBPjTmB
pRPUHMMWQgHUNFWw4Bw3do5gudqUh0kMUlzAUzkQkE45BHTOOwlnvg2NnA+nYHqk
dZATSS5rKSBrexNtmulYvBhYBg7vkHz/hjntkiBkeNlA/M3cBAqUqIrM+FpFGq+t
LprU+szfEw+f3AJb+snVtsRH+DSv593PbQxNAtaYNtXQxlBUEZVlDpHa8B05zs+3
5kRSDT7UAiVLxCNeh4kV3KL9iKutM23oqVNWlQwsqBuY94u6ygqJZO++Kg+2wwMp
XO9OUIuKwE4LKnuILUWTRyWFBJZA4xK5TGgMfGWispe2uqlYDfisme996s/narLK
IQhLE0HQv2SbThSQiidGrzx3zPHF2puJuNvV/BWBbotfl1pv9qysQxIPfTyrp8Vp
uZ52P+IV9NaPJBjm/sp3p4ufsMYh9R4ycW9s7WcgVARSJkmB+oSyEfpOGRqUPCB3
pLKoGWI/KsQ6uSft5N+BoBd58j50RAzXfdtk046/ugA6e5brWTMEGeuI/jZdP4ay
O6uPA5+DvXSL/XAthdKo65jM6sTkwIQAS9I1ZyynBJa5UC13Z1yeeBu9Q5U/CcG5
HwaDgiGxECYERJRsngeJhPBr53CeKIbqmaKAR7FzcF/g3JeLEJsU092mvxEXDD5j
21wS+8sOPZ/T6y3Vs0IQt/06dxqPsfT9PL3eJW2zNPR7p8AetOcW4m4A+ocf8Css
2iMKJ9h30Grfbhq1DZ2k5dQz7rm0xzsszaHklRG+bo1zr45ZPA+a6woNmj1oLqoX
JPsTN/ajHteVnLeDO+R/ii+XC18S3Oj7UkmTnJtQfyMkHIl4N2Txraxau/QQr8LM
XLYJwMIDS1ZZPMVikh/Si07splUPtiUrd5rrfBfBcQ76wznKoxpTJFQYoyF4J+/p
fjx6kpKPeCBN9yc3UIPPb9hHEZ3ui1AXT3zBJDn4ukb4qVgr9VHinUTRvmCIWkee
WHYPnlqSxFIQyG+alDKN7svaysOglHnOk3rSYFGlJ3Q3mmPuRKLkqG5JsXiyfv3Z
2KwGXWLNAFJbAV4gBHgNCxVkpH94kJwb5amnPzjBkU7ZC393MGT6t4ffPMbX+7+5
wSsNttQzqvgm6BvZCDodZGIES5XnHZ2rkft4oqiU644zZ8zsUOtduYjCUNinUobQ
RLmHi0rf158BUUHkO6XtRWreOTo6AYQ4W9bMsSjPUuvH81LQE6FqXR38LybsEkJ7
se3dAQBfX+dhtjSk8KPgsh4QeZFlKkQTITvI4fp6zz18JaiQP0d477aMApqunfx8
iLPN2qLsETDI6l0aOF9NOOyNB3hHABcBBLlTPeUlhK9Vf+JQRm+gdiYOnSMYz2ur
UrAZsWzaWlNPabWZ3IVyBWZSVG8m8qQTEj/wnpmWnjfw0CCk1wHnCaExK5JyWM31
p2OpfHLlM3AW4TRjo1IZSlj7ADARxoWybJP/W7WKOBJH2MVRZFC9g+TDVPnUPxix
KqQ7hUD0lz9LhKRm6tlSO6Q08M7FEbWbexblNByhoGMK2A/j7yod9J95oeWRbhAc
dmSgpqeyYCHB93tvxluVyvv6C1pLPKyUTgq4Zx5jddW+qmxyIFDWsYqeDDGiLoo5
ocMxPADSluxWdrURjsKOLdOvOYOH6NwrAOIogwCNre1YRTNIl8y5ytxHjuK/guGQ
TL2k8mFoSflwYxItRUu/Xcc5TQ0ycp/8L21bRQc9iqZtYs0atxDqxjn40RpGi3aT
tGxdCoLs37iy5QXW1jRypXru1/yDQhEjELln81Rorjxse7Rhl0YR9MDdSvYxr68H
NJDnd/1CZurkzFr0CEB2S59fFyfKteFbMf6NXw/xD9FasrcaPyri3NbW2RyJHQ8U
IgJ/TVd72cEbHGtYUWWXFc6rYvafY9v7xgHk0WmykGuYUVc6Dgz6Oa75AWCChGd0
ZEgTt1bLkcepdMAjTkoGLbkWIxxUlO1vG7abijgm77k/HUqp0qD84bxuR75/DO20
wlg4XLy9MTr4jU9ahUsNahMBczQZQfu0wcuDi0yuPzJuOtl4r9/NyKe+R07sRpg7
51eMytJ1QRflUdtJoBqEQG/SBJRqVWSIHqQtEcNTnRvPjDeN8bZYArvp+N0plBdq
yGmmLkPPs+9WBBk6L9M+TRKbz1uZohDiVog9K0rflisz15hG1xL79V3VthZV80ZP
mk8gyGW2zFmlhO9aeo8dWCP0T39zLwVYIiaoEBm+oQlfkt7tK/TrCa5Gts/ue3rs
6yzUaBRxEGIclhtmEoVcaXc7q8UzpuNMEywlaIH75rVTs2Z9Y2p8P3TjlX64Rzfz
qbMOTAs7IW0j8xrstpV9U7Ax+TSrQe8YrGjIKxAoYBxQwKEhafSm8jOEHZ5WA022
A0/wPoJoM0RutG8+utDwvjIX0Nivj4dJ+n6UjLDTY+DF7Qo0DD1XmXMaHrTydtGi
vTrBktPzAeUDaUEWayFH8k4bpFGjWstlWHLBJjsrAH8plWpEXi15GEqE/NGoS9uu
G3xmMLORmZnQa8PYkn+oN5+l7T4ufCFULb9iOgokQ3To06fNh4ZgKUqUdaOgmEjv
eH6lu8URPUASrO8dYKih8bVb/Qc3c/XTL9mIjF9m00IWNxD0r/gaQiL6iHn7t2bt
2IaROhZ+JhT3zFkvb+/rZeeVRE5HA45EWHlP1vTKqDlBIqZFu380xYk9gDdazBRD
dYPZ6RmwM7lrBvORWnF6Z1b8vJWZaa1ITq4BZPSSduoUvfGApyzhYjwbuFK6Z+lg
YN1/viYiF+RhphmN9BiFQlJUQTKmlpPo+MtmwhHpUZd6BOOBhbTzevT2R3dqMzE4
JmmTL6rGueruo0n6HDbGPXSZmBOtY5g96EWhvNrglgbYv17PxVtw7yVTbKzXgl+q
cVbRI57W3hMsOMbe8dsyZ+4tD8q09K1XsJSJQ4/9eWKnaXgRn67HmHI4MRzCna+k
+a8Z0b9tuemXyobfCliulABkZuDmA5TI9NC0Ou0UENO5JwTKqy6O1ZKycp3tX4yI
ZVp0M3V0mB6srR14Iuadz9HhT30fTUni9vUEr3up/sFnTV+zIMJM1qN6yRBuyzCd
IXVs7w/uX9/ECmWeA8FVx0D3ZQS/JHouAehpkaMPzKLvCU3sQHTRejfCVPBo04UK
+vo+Z1U8u27UjCEzq56vyQ0Pcx0ZE1Qn/0QT8ULNpdrxzSLSSD5MTmMwDX8cIwJu
CFnNLcq+gCIvvF3629clvjEIOwLKbSRYtLH0UrwP2k+zSmB6Wqa58EOMFmp4vH6Q
R7b3s/7T8JpBMgMMHCvX0UEmT5Umx/Gr4IXa3UHLiliBfdoGdnUTg7KAXs8bhtEj
0edSqbdAIwvUTIxTZvdNI5zOuB4I3xpR/PLPlrjI8eI1lu8yT3UfdJQk4ikxCG3u
hkWryciXd4vSfBYbUuOtnrhhEG72+yJgKrCi7NZDyvt+dgV4UG8jUgE3zXTHU80j
MCCxy98pz8Qg9wXczSPjvrqb0JAkZr3mYuttnQ+wJIXkD/rt7NI0cSXMrxohlILR
jA1Dj83NQXhwRrMSRfgc/eAVTm3//tli8vedrrATnexOw4kE+0yq74JGkGcXpWdP
bhlDQ5jD8mXwV1oKmb2z+/SCA8HRvk6EiQ5lK4hToyLGoBqEMhlHr/tAu1rHUNuL
qqUdA1CJMcUU750/SmRntHulgCRZXUfcZ1b7lOW2Jn5Izkw2Gsl/o3EraPXJfRoi
qli4vz7TSDQqhZ3PIGvdF0x6h376HTRK6auuedCnT8myFv/Uw4qS6vhXSRiMzb0z
LFPSaoZTKXvAH5CnXgMShqMaau4NbUnVwsOjjpJKNiHxLvgDefM/DGJWYUR6ivHI
ouu0jiIjYJmeIXkhTTWfdNDezUh1gCO/7vqKhKIpcyuohVoPuCLRZtAQVddbYanG
fbJRjXAA1AVz4C+ynE5rf8itu49XDM3mfaP0eDfQO63vtpDg6rdKJCPGnTVGGskv
t2L/d0WJpTZo0QH4MtAlQHrPu8/DfkC7Vr9RyVwE9tW1cYzvPBP0JqYOdCXWEsQW
90Qw91VHL9C8VgZRIniyEZ+yaFMgQkymORiUxc0OIcsWycE6nw9vVhXhkYJBmgLq
x1J2xDPfnRuW8TOLar34RXCVe3CQGPjGUsfYLJNySHzXUSjUuCe5vyIUKxzN1MNd
3Iz3vSMdWQKPw2cjHiIg4ZXyQptD7XbfdtkDbrgtiSEJGKYZSEnRNgbxBTGtufR+
n/t67fGkXtYBSz1WZ0ziVB3owwh4KBijLARxRtpyaoTnpnDJKYbMOoKURkbkFK7B
Qh8wf+tyOpW+/JC/VdhFpKxI2RXElIgnm2izY9+2sasyO6+tgiZ5pp7orrJRFJ8x
mo/O90592J4naDAdZnGKxepLRVAWcHPaAyqJg7NtTOaaRkKnpZeDaeqyoOm/d+KT
s4dq5TZNsP9vzjt5Rck9jW22zBUTGKSPfSV8bxNHCAjmv/9+8pXjst5uPvLPNpei
jLQocLqgcPjEDr9NvN6IinFSTurxHReIPVG2MFrgpVW7PczDbX22szWhBK/cUH+l
UYfWxZa7vi3UcIg58fj3q2bXgPHo95kV71A9Yrivo6UX8ZXknyI0wiCUO1YVFcZx
BsI0YbB/RBS5jTQ21isbQAyjZkvzXm21kAw62QPc67wBAAsX37Ir3a1F2CeCTF/W
9mmdUi/WRzyQMSM/wb6U7Abq2mxUW4XyZZQ2vEWvmfYEMHcYpALCKyLUX5I43SMV
xjP9p8eqon+Q5EGteCGXFexw2jHntsJlpIUlzk7TETm1oHzoK3Iw9wDlQOCy2Jmy
lhptTzPwF9/w9U2U9DmyHob86zb8sgiCjpTIbvY9nCyKN25C6EPJoIzwPvjf97OA
dYoxLOBRqHO2WWwPDKGAxsGBz32o3dqBcSfOPW2RnlWvImdIlHWXPTwViKZqATCE
x0uxNpRuF3v/WaebMviw4Y/ZIGGykbw8/pWMTcUAQoWA5MDaHnPfR745ir37CPd6
uLb00pdhaWHNf+aloo3KXHpHwTbvhXYHYGiEfi/zx8fAqyYU8CYqOuPAj7yrIGlg
ZZ7cMsN29kU1JNcBfKPOBcPKcryu6/a+puBGopY4PWilUTDz9Za7lTX5Av8riLf9
Wh/1OX4ttnPB5JQxqNo5lfLRaCht9G0eLOL9MZooy6/t9Cyvlu7CeXpDIsJRl591
rAbQOIU3kTSsepP3lfXIg9Z2dAdUzN3xb2aBjcwPU+dAgWwdCP9b7Ieg9yzMNoH+
3LUeq+Lc/bVuZZkwMeoJK9U7j61sNyGYxzwGAcflznJnjKK+9XAMDZf1vwLKeHT0
w6g2TjRefgfPxrmWGkhmnRJQgCkY5YM4rHyANmPth8ggEor8l44zi0Um6uz1HX8D
BKzVsrimPST/zqemkUu9ruGa0dViiaOJ0ZpQyb4gxW9c2jMaUcXQhRxQMi2h2GxZ
jSMTrZcD4p2Oc+GHpkXDU7Cml3LBjPSyQLo6tqcdB5V+CKgiMC7RjiQiR8C4wyfG
5Vuh4NCzBhsh4vd+w7Rf8p4XEScLYhN+bs8CYP4iUlidd5j9SheoUEjk+P0u1TAS
//T5hsE67g8Be07+tQ0O6vkLASpsKcq57whYkbyLUMxeKp+yJ546FHS2mYexChHn
Douo+vf5gu9p9u2I8LM2g6u+fP2jmLfw3l1NeFHdDuV+YnCn1FxW5AM6WE5hwCX5
UEgXU+XppbWvbqP/6+7jffW9XEGfxrfcH4RVgi3nsiv+o8I8NKJ3xTU76E9TL8St
mKJynpE8FhjBe32oqBxtPntn0yrq2ZMwfTfIQWshWolJBAKWY555DdULNnVfuvwR
cxv0f+CsSDu1Wx3DpWfunhY9Ko81ze9Wy0xvzNLzVxkdMsB4AaAZ76h9mxMqq96y
GiVrlOozpTFkXEEcvNM4iAimoL8JgrjzvBmAAZwvQv4dDXqGRkAY2XQ1oLvn526+
XzVD1qnDkMOJNLGStOe/u9hAnKzQ0gkzQF4mAG3tEVnAncjfnvg8/LBQ3+rd5zO8
GjZ8rzS+R3t8OOeRn/ZkBs7C1coLLv1/brntflP2FiHIJwcegfD6Qvn4Im10Ai2M
E1KA9dviFNGO2klhJKqXrEfBhWfJIj/WsrRwC9xwTOip6ZJ/Vy05bFwXnHGtu/yA
KQg5Ey3FtiEQFUKWE8St8bgeUP+25gZO0jUG7xVd3v1Tpt15Y4mxkTO6oKuQDqZc
f/ygXGSxrjwfDhaN7S3VDXGIkY03gyOPM9QQPbuyKt1Kwrj6CUGq3wH+ZXeHnOcL
6bWGzxG5I+C3m/SEadPjHQvMj9xSLWVl9ViYB27W1Ddaxb5Z9GBF+vPCDVmQUuzS
oamIgXcetsc1xq8Wmh08Fk4E0g4RC1Izy9x1aP5vSrR16e28nFNZ3j1IQZ3bdInT
kxbU71a1UVsDe2GPcgdZg4Os4Y49bmRs7/DSOqhBhl+zmN1dUO49hzlSjRCXTejy
H2LzAQjkeC5ePkzD/fMPtDCh1xuzxsXTKGwRH1YfYNS1V1WgI75EgMMEjwAlv6p2
CBdNNp1yNm+a5wkbnoL8Bc0RHu3JjWipOXoj8aLKj7Z79FdhWJhFCG7DJFKu9LdH
gRUxSYHfvTW1Lv0jvgL9HyIwzxpMTjgFjlknftNDn86v42UngkLdvCQHRYf7iEI3
+ZrnOtNG5yIOkjAwKD3mRjsIgMJ9dYU1NF/Meix9J8turJwGGCvQBxJcu/DS86gf
ZLjZaU5WNIFK8VTiN+jUljvt7e2PZAWJwdXTqlr2L9rEwgqxb6T5sBxAawfOu6ei
Yx4DHzijYhvVjPydH+x0HNe3T7VxjvmW16BQTKq/VpYyU/dnkNTra6q3VTJ0kZKX
FiWMy4iEtM9PvE5sH0XoSeL/UJr/pfLPbeLaWHhz+oAej/S5FaNM7lQ5Ewocowk+
P1fqbNZdHvrSin333YFnxXv1LewLtN37i+XXQPkDHR4ITX93+Ufev/gH9+8htTuz
aZAFy40LPhtUTL36Kmz1KwEpV5/0i3XD0dJV5d11KeXaJeec1yrOp7xxKq1DpedP
CQHBS4EYRT6ypIKxlk1m6YsNVUMp8Bf6c0j4P2RPvhKknXbkGJBblGErUT/9uzHM
wOCchmOddLfUAOJDdLMFpSauvDY2Ew8iU8BSnf+UzIcdO8XXoNXdprK+9HOgs07V
GILJTjUNf8KjZooqUyDGilBvj3aD1fvXBUH2+qyBZDSb4JEuuh16lYmbMLjklPGy
dOA6n9Y+aDap5MUDc2p1BmX306SenmyyXZvTUf4o4Mq0flgerrFeSd2XFXPw2JlY
7hdTcnIxggZaoYb7S5BEtpuA8D1KRHLR+m6/n3kNH+8NM/S11yXgJ+jImVilbHNW
gO5lsUrQmpJqk9U5J2Q26+VxPud5lrLpcyg85LqitFWAK9/24kSirlAK9sr1ar9p
F6K8enmekmfkfq6B6354lTP4h9JwQHakcpW0e2vivzRFM0GgP4d3nthIRQPqDFqi
iqE4ReIpAv7OeNYqiuT4qYTtrgkUJ+90nJrxQo2VAZAjzbigtDm9mF2bl1tf50uM
nmjJAdnrlOQecE4kL1cEnN/iP5TEhV/jzKiyHWt/E9jezpP054XKqYbVDNXoHqF7
mfnDRfOAqVO6DvMpZkZfUbX4MTJA7/Kg8duXmHDTG/N+dJ1WM2atQRSncMY6c/pX
0OERa3OdHuhd/dPmmXTHchPu7NAhpNuWujoXUcRHjXVYvVvfhxYK3RdYUJkQBPrc
R4Fi3lGCd4miOZYF1UUnDcz3GyOYwzWruNP45wIi4rOIXU0dLZ0cQNhu26sCY4DN
+/GatoRHbgXxyCXU2j13VQx9fcnMz+aLUnLDD0QUUqU08iFni2np/DBON06jmoQX
+tnMjoiLBbRit0BBi8sfNrnoKVCPoLS5+1F3hS6XxpI5RSK9IlSUXFmp6C0wqXeT
RoG1HTdObWGP/KKMiTzSAsO93ASxwJbg1gPs+C4nBVzsC+LhhK5TnK0c435o6sRp
LDXl4IIpTNVu1ENKylQiqmaxclIWccOtLXapAfGNlWS9NaSmStg8Bx3ZvGx6jB8e
px4nRCO+WKiYOtlxcojUAvg9mHpnqTN3fU5OIiWMjW3eqfhrZ15ML7ycI8dxwX5r
MAETmi7chNrSbdNN9Uo3QpwiL809Wxu+tP+IsHp6pBphNd+/F80Bswv2xKo4gUnt
hzcx5Bdm95hpO1OC/sg96o/A9q/Y/GkmzJ84h8wOOjdtlktzj8LIeM1umfVVyxyC
2vKTG/xxn23zSYKMqB/RCeCSO/YxlnA46RlkAroqFVC1jFza4sC3KfbiZl67OGbo
yxNXux3yj72i8lnezHkHSGAsCFA1TLGn3raeUYRqBirgoDipKXzmhjB2g2xki6SG
f0oyTWV306feb3TERY6lOKMYAmE14TsACPTJVZtqc8anIX78QqiQe0A37ThHculE
ABFlnoVCX51y4nsTvCmbBtRlNhuItUtVvwxkwMOjSrLpgiovamIsBUvHmN8lW9SW
F+F8T8lPzIqxJJ7R9QgBK2JM4ONSSzMsY+Q8d7lVroFo9+arSwLQPOrNtIvdSRrn
r99rHyGcN8quVZ62oP9Jy3nGb7nyfIiAzlGVXMfmmh7+otLvY1mED1Iic/tJdqeF
ILMY2VQSr7w9wk54fNK2i588LfGj095VXYLhXKWi8zx3Q70EVz+L3EKe7yLvPkUT
6rthjd1Z/O7ukz42D6n0dn6+QrxTvCK17AUyxJsApq3Sw2EVCXJfFkBOq31VCJPm
h3o6oYptm3sy169sR2BscIdYY1JOMa00ThUopSblhAge5ritNY2fU3vVtzqbwvh7
NQ7J1RNYEVLHNHO98cA2SdjVWvAXYJ1Y2yivbgBdjuu5cD8zPrDfNxenFzUmpJIy
6uFg0nTlmVjyGOBOtpFBQ2JrA4vfwlFHqwrARnjID6g14+98VX8K31r5Vr29bDgJ
sCWkCiBgse+wHZ1ZL46AHxZroFUuKCC5iR4tXpG8jOW/T66kpI5uUFRXUfoLOcN2
pTupQVvMX7vk4L+flrhk+IMi7dAavbYbrVO/c29ctv9aaari2JB4preUC2tGH1/r
3CP2P2tQC4zI9H5uMYFUlBg19Zle+yaxFz2/mV+yGeNk2STHzG0a1fOvorWvp2Xh
EsmBsastN1/jAsZ90n2DiEmIAAa7w2WRk+vdwVCQOtncfsr90OM7y6/ZlJsZRsNU
V2ajoYVSGtBpW22Z0jfBv5W9VBFFTQJtiaLi8H9xFwBTEq0CNHUp0TDWQfjcLbhY
QGO0VVdcGV38QTdLJaGiowLC2PEqw9jPPmQZ15HiMyVFANMhoRMbsiYc/2dTSp9U
q+aUWPvJ3/SKaz7kuDiDRmDgqknD2u+8N/1XUO06ZZcKV6ZuMOK5OE14hh8utfzt
7+RncMKBH29nPuQjhlssWqpN/IrBpudwdrFAS+lKFQNNLBZaN9LzNt2xY43ThDEL
Ga4SNs2BxrFlhctJRGUHCPs41xQvtEY7WMPJwB5h8t7hd8J59u5P3z7ajGJt7Cls
UZKCt1Qblke2OYOK9Szko2az/OJjexHOnGfXEULsBhcQkOhxBPD7YSA+Xmp2zUul
8w+/o2nw8quuCl6SwlwxkvZsMK6cF2swZ/jUNcVkFbS0JgBmp0Iokm5nVhQAEBRE
2D8zAw0Mwjdt8j3Nzj0na+YfxgfrRmOTB9MXGZjaCejP8p9j3o/FqM7Npmyew/ma
3mySFbNYkCGVbQJj1dYQYCzhdym1slwRBAEsnkqWbfM5bzV4oU9hLtSXtpkEy+vL
WUrDzW3pvkwhaW4o8Dk4rXfNf8cJ69YmVjLPhdWYv8bfibDPnrK5ogB2ADI3Y5B2
64KK1WqkqN1a9mC8CZl10Ue2Ln4Q6oeVqiFWLaPpkkCEqapz86kWG0y2tz6R/Zjh
YXrQYNTlfF2YcFdO65q7x2p/hEl990gL+er9jTBgnovMaHAn2IhESnXnHhYXmGxz
JftLcPcYo1JwOFyqdm93KUbEwRyIEKrIuEaXg52lwkGuWPl5dPGW/8zl+S6jW7Ce
iCvUXYdhduDMnQXFcZ9mx+OU9lzTwTPTDdBnbzzoBa66i3hfPrhXNf3zyzvkUTTO
eLovZkWHNQHiTo4K6LDgW7Q4Gigi6KFRyyliiHGfiPjP9UQRs5fXLEuz2l/Fbewr
TDhjwlPBfUTRCqVHskV7gCQVYTYNKfzdvL4V++WpErgqNiECV2paNGGs0hc4sp1M
A0/S6EH10AkPmnut8bTDoBRZ1PuDnlWKex35Yk9mB/xk88vVDV5uG59z8OruNiGF
vjxvalPRmUum+P+WQsdfuYwt3jkQF8N/EwBl+IP1j0hpga4+9Mi02LvjRgasbDPS
pn1GR604NOekeh22fKHSh7mYfa8dugpXY9L96K3Maszl+2N0Njj19IfmoU5mjOJN
ON1LgnCsOWQtCqVk3R3rOwfWr0z+bpyadLAowaDW84wDoDno8xkeLmJTUdX0NP4o
qAlBcoLXnfR8gPZLqTlH/MJVyECQ21jNVBo5d0ZxRoVIZIfJZH7ENwRo2SrbW1As
gRT6dG9uoD9EWj9vvl0SCGnDiJtP94MhsQRJ55dm9GKNhxriGfGHGIm5RKvXKOr4
B8QhDJYxZVPUfnR+WfPGr1AkVspNh/394ahVYqj14/gzV+NqdyBNWB5K2WxKhWkB
DkkX2t2fIGk2tdjzBwl4CFfyaIoWv4GOo3RF3HHJQ+InsH1IizW6w5QaoJRX75FE
PEeLO4pvK9PcJi2bzhU+xaz44kJgzDV4AuQrXB5UEUyuoBv4tf7hcOPV7PF3C6+w
MR4x0JR1lGia6wTDT2R++/+7BgA++aMocRuXVLJ02Nm2vGzcwzcpXVg1eCGOBRav
FXA6KaAP22Q9vwK7gdzRXi8pskau9F5MK9N3JeW8vpcpe9rohDnRwKQd5B8/H8Xo
qgSBMMj/8Fc9cxqB+yypFz6I8ZLETTcDVhNkXa+onKVrW14I3Ig7eCWYZS23F+4I
oFeBTfLmfHj25/vQgyK2CwD/22P+ZX9Ue+w4v/A+f3nGRpa4+iksGf78HALkHX3u
1Ch3K/WcGF7l4Ix6mlhM/HrBexbAY66UuwMMIPR8eKkfUOdu9sFW7ETUBk8JB8y3
ma/CVXJv3swiGL8AR7D43uYrgRkO6fWh5uWhsTsHiSr0D8XlEgPtrXI316Pyj9lZ
ee+9LJmbmbsv0lCNamAk3Qgpga9SxE7uhQ+nVn/xhridRSdgGgKZgXnD5bNhm/UU
3aaqikOOggLbcPHQukECikDIidpi+NcxigKOvr1Wdx32p7Tna9nsQCRVdzsepe7L
WHcKqPk00I8pVZArusdkf/GoKyz2JrTifAeOxBdqTlkG5nGrOdcFzpoWGWvLlL52
KYHbmQWkaHeQCNX9TOBFWwx3/woI2/7qEAXJz0sFD8I/yvb2FAXbAQhCewKgqbvI
Nc4H4W/6Jgtu6UpdrWs0bTcP4ggrOoWCWRiUEZkKvJMuufStlB2gz/qWHjT6fTXp
iYGoIxwTOyjd+OVjgxtudvaiUW1Yl9RSUeCmgr6DP5HSHn1TTEn29OUHANqOyjBm
iBGwAAV25cFTqupFxTc1dtdN8sDnTfv7XDX6BeL6ftH/pUoqMAGCRVTUWy8PINy/
ti8LfqtzDGyGm761PFr92H84/S5+5mOIwcfLyjOmwt2wrw5yUNIPMbsOzy/Fy9V6
hvwunIzdOnDFbk1UeEXTEgCX8AV1JzoGs/5cRS2PxalFHMF8Mc0QOPn8K6w0Na7/
CFGN/tRYabk8uYuqtA6oZj2hhjjnyA2Qrxt3NiH+7lUCclfGPgNxC+/FjUOnzavX
Ju3+hX2dc+s2vsNgp1nJZTxYCYNBcMoGn4ASvkQ/wmfw3RXTaMbTwV7FG1hTRlIS
eN3odvLqDGG1MTWu6/WSvrWZpJKmgu5SogpLHiYKbdas2PTwOZ0DV0QYIkcCEWsj
p0aALmv7zKEg8kbSiiRY2U8MW6sq6FvLjZIujzt80NAQ9fM9D/tI0iaUojPd1f9V
6cZ47ETVUlBmoQzjKWDxPndQpGyS/mxwy1i9Lyu4fKNpKCuRiP0uKZgzAfdYIF7E
X+dfc04ui5fwc9qJbxIP2OF5Xtsd3nzplutGnnL4/Q9hPhXYLUxw0YzaYAk1jJpr
gjF6Y8wn0qecUO70Tpe1i/SDybh3uYWHSSrFyQE5VURjXahbWtDQHOaCEPYeNSqK
fAKUb+p+MzPw45QNZagI5V3agvJ8QAhqt6yt0BzhiyQ1ZWekSKJtoQqamV+liEXC
iLYfEuDNaTKmfLd3Ct5D3a3idse+kvgJciO298glwnnMLVRUDypjqMGQ/sskbMYQ
sIM7DGWu6NtMcnMsluQ7oMRJv46xqyJkBhKgGrlgsr9D3UpMhxrEvSryHg7VarHq
rbXI0+z0KzkygJTrr7AIt/Bi5qHuwUzN90u6DZgPWDgV+x0pPj0iUDxJYEFKnl7a
8aeWBDLbYMHtp5bNZVZI15pml4/nME19q9aMsUHnPImRu0hHwOf1XlnnJdUbKrRn
Cxue/XpSdk+oRd3glPoR7DRGjN3P+ZLkr8BqwiU9ldGawUZLufsOGklExyi/KH/m
x8yRGGz8FpKl7krN+EVY/RX6Paalte3mmraf7yJ4Cfhsp1Lte24iDOz3LecZTFq+
T0vm9RmmlredMzCHC7sbCrGXiPgKnZDH5amOQ3YucCI++clENAD6K5iSep1wEvmO
1pV6OTJp1DkGsoT45tbfERew0acLqqkJjrLbT4/9IZl/23Znf12qU7EyrjbP/biS
CIs2Fa/qkUgLBndcPWOAohYzpZM4QjXefQ0ePMS1qWZdqHCgESvSca3Zol/hrgGF
cDrl+a71VhaZ7bO2fV+HvFtrju0piKOm9cWhMo09G4ysO/ElGTf+06Sw7QMJ9rCq
qM30hNNPk58KO0EnkMpxl4olu9tWb3aOb1B2tki7C1XQ2c9ioNPvRQ4iH0Q6+jMv
Lp7cNtrZKthsNI6TZ1GEPD2WxDKg6YvgHJenCzPo65XGVYqdJVo9QyA+s6RlFZzo
0NSj/XdtxN91tVY/0+zhVaJGndT6ZZg/0IfdePWUu3yf3OVdYo/5H0l8FLgI8cDM
MwiBF5mvqxFRNYaSBSGKtp5LBYsb191jqjKQ50F24KuOCYr7RV/QiVzUkvgB/2+E
igRp8+//cpr6UONzKGpVAUoZskzX4KWIuRg7a0z9pvrrKDb3/JUV7Ykdnh7SQQlX
4OF+Cd8lmJ8s9S1Qmq1KbwcYrfYF9/d85rPfpF4drYvu7tGMsqvuX6yRXrjIh+GF
JVs/4dflGmYoCsW99uL7fnTN2rnzgDr4D6hhBl0XZ2f5MFzE7cFqIzw2r3jzQIQo
C6UgiY/H+hiJ3qRKANEIYUWpecHloWJEnN0W37TwVPkqqUpGL6f7+KNWkrbs6e+h
7HXX0sUejQWfVr+Wi+Lu70qx8n8A5lhoFeqS1CYpZ+qG4iNzCaqkiM9DYuSkwoxY
5BRCH3pboeYun9Z7VCZB/z4KQttchlh3cWO+ibgzj+7s+ttdeRZkT8pvu+wvnVNF
b+NI39oh8qin6258JUCvYVX0DmOua5X4Gh//Ds0ta3yiqUcO8V/XR18unReQV1TW
7BTak0Hgi0+UIM8by1AmSCbw/NK86VKStB9nHDDv81/bo94Jn0Rsr3y+2mR9DqTe
onlIl6Gm2QFcvzPoQS+UlG1/sbhUsHKy8TGM2ZknC8EBAX9jCvjXnz/XZvxMJN+1
k/nUqSOnUXe42cIaDSmxTbtYIh8PUIbOkvPQzyriL0fXBSp6UWk8FAfaI3lQszQ5
PoOzOVKtYxoZH0UTPfUHPx15/EbgS0VDB4GKMznvY34M6XjhEMP5y386Db61uDm+
mN7PMuAFpTZdyWfuP0LyrUh9eLfmmAPPc+687uufc7o+1b7SpcYxqunWsBPueVV6
Flha4gaNcFSeI08hmYbTI2Y64m7GoJQNMgMwphiksfLY3orlkfQdNf29XW4NlIlS
Jmcv9r70hDtbznJ/LxgRNaE/7mxSq00+PkWZAxRuEfTj6oZjf9AH9dhjEH/vw7QV
rLN8Vm4GkvkrQ5gqECPfharpPk3JiD3SR85TtbgqajPyo183K1QSqJp47GGUrr0s
zq3rfqRRD9XuWV/vAlhMcx9PWioKTUjy2Mkzg0k/xdNAg1b7zUCVMzd00WiSg0RN
rIaOYA0PflEjlH/XgjrQ3pg83pKuhK4Sr19EbjbZt19EvQOrU3mzUHCJm1IpA6VQ
8MHrcRjwnfMwgdQmqQ5FFMvcSZJxd3MKLuxOE0cuVOsj0YBGBnYg1C4SogFQYuQY
v8KNd8FpujuKEII1K7qQ7K/2H7zqEX4UjoLi3RCa3WNFO87GXVelTJAej+uWBw+s
Z9fzBRqWuJ2fWZaSrEPGeYl3Vd+Zz+xLjN1S9Fw0Glqh43O/mJrpnrXDvB+vteXb
JjUO/oqFO4B+pMebm43kO6RNv+EsEa/N6ZFht5uNCmO/nEhXexV0zLNC75ArqKIo
msccJ7QlgbdyEKvpxPLbpTxT7aa7aGybKJG7bdRX2mp9ONul4GNvOM1lXIE0Vzis
37ML3l/4QgjmLvKjDjTVP5rwS+qzWGsKljoZfj/+B0Oc0I4nKBzITErBA9X52rXY
7HeaYTZxAWfRtQ63Kbnsu0IdZQisG/M04bmTvhp5Hxne5nI9d2iPxboON6ZTGTAu
yo612esiubhKc1btm/Sef1L5Cdf3m0QGn7EpmP+OUNNvxfBbx/lx8rlqWEA1GBex
pLQic8HIO+1agsUc3ER4Xkbu2Zu9Cxk672Q1SVPi9CQRPA4uqA5jYVMkEk3J/EIL
sGjTjtviqvINVlEmSfk8o5NFZepGYjZXNlTje/0Vkq/zod74ztxNwuUZcYOmpnLq
GgBiCLOHPBsLtoGVMhR3zfW9sYddl7KfiNnCfCL6he4wHLBILVqm0a4uUJzp5yCu
gbDsjNZCnmVo4dWnHqpaLyEDiq6m+UEqYKysebWAyEVDJTq3r4SdP+6a6umUd8Ov
BsrXbl2i6XtHJFhYzo+JcMkLKz9jQEffoTXfRvK42C0Ta4z7C34IZOFqNijFQswm
e0w6woaDgsdsldkvnXOkLK4QBOezOV8YJwck7p9Lr7Z7G5BD91h6v0o0Q2ZsmEvf
obG3ejunaPHZR1GOt9r4wAJhBrPsumav+QYYLMcv7/dSSrUCgyHqZKmssrIsG2fh
PDpETUyT3Eysxy7uJ7ZrPlBKYiUAHLUuZ7lyOPbDtlkhHRu63aakcQ5XPgZ4OApd
kyrZ1/ZqNQIyfJoMLMXwong7Or68NrjbE0E8GAtTX4JxWDzcLviy/p3LZxTrmBgP
1PpMT2nZRRtZRKQppSk6muoBTbEtfi/p38NZf/sHQ6jR+WMRvZED55+SKkCdcbJU
5U2z5LBEe/5FoREW6NnBOe5K3gV35Oh+4FFxYNrtfBjUXgbco1gZelK9RQvuFMNt
CIrOWS8lCyDBsOHZQynvUVuxsdeWgnKmdEFl6knYFp+KMJBbUT/EtFh3DTP3wGrb
VyGXqMEzKwNmyEakaOfDWG+sn+mThk+9qZJOzxWtiAv/9vEXBcic7ZzmTdbKoHYi
J4vtqf1/l1KRyKopP3gzQQ+xI5C0raLkMipLwR6/gZXZW5/WjDg/bkaGFnEtr2Wt
e1+I8TFdyeKw8ouiW8DcbQDJM56dvBjcoVrOTlwNXpuVW0DWX8Eq+SokYu7lzk4a
c1/LP/SWM44WTAySUJ/fJYBDo7aBt8XENAzVyQPeUJdKH8fbMLTLORtlAqFVG5nv
B2c9jqvDhfSDeW5mTdQnKoQAG933G3tr8sIzRRYHZE/NKVlbVbLUKTRN+XO95djx
whTAFKjAgxf1nalqPg06NAysrNVKuVOeVhIVsADolrOgkzYcDWr2BgIJgtEnqC3t
NL3MkGxXpgb1cdwx405xOpzxZ4FIFHtQ6fqcIHQGmd6tLYrqUOKuGIMEwqFJu5XA
IuizXZecIVy6vCaU04NoGPaOu+p9fr/Ey5BzgSn/N0uaaSX9MJ3LWlenRvVtWBNS
34BszYcHu18w5w08ksZrAh384i5nPPji6eVuPVejTAc4bAbRToDwP22ZX4kB/CkN
JEimSoD18/bCMGqKFPhl76wdYdCclhUlCPlx5S+4S0P68D4ipjzh5NWaA/jGC6gA
2BBgvLNeXtMML9LSjJRD+rZYwcQdEw/VGihETqVbeAnKGP4Sb8gEuEyu9Vic1mBh
vYEeDiv/PevrTA05szAe3kJMvUhI6dA8oLDhSySRyPjrKzElHbYWcK66vVkD4ZBd
NIdEbJmZAyxHNwv6zUDgSfnebfAvYVLfOcSKk/obBYWPy8XcBk1P5dYW1URbkF8p
DsrdLpe5MGXdxivpFELHWQI87jSY5TSfFhRIOjvMPLe66/RbHRPCrxsVkFn5uY4Y
oI3ejf2CMFzuAWMxLLIC2Puh0jYCUHHbuvjmfDf1yzTOxesfcWLvnh2CzPYqJwvB
WTJhYjN47v9+L0aIaH6N6soyKt2L+qIEN0I1uasA+1/b7q2BMi5sgqmL9myZikjo
AbxNkj4jDuP+W9L31EBawLr2oyihBKrPfxP5fqhdIp38v2vEOzyd0JKwU/iZHZev
bV3x3JHKoW4rEGbil9lnykAEmRz/SbAYdVcMayyM6huOvUerpPDL/W9UNOUGj4Dt
9rM+2x4kbXFEFRdGEtJGxh9rRPJLLQ5p+15Q8H48+PMtuDtlt+b0w4C+i3sFwHFi
f1tZQejtoJhwkgGO2Sjl0m3KdbLo9LpW26oGFpsTA38Uo+AKd0lTWAWbPyXSARzT
ZO68wzl4tgE1Kvhos0DDL3gA2l7bqWMQgLzfT9vXuTMfP86UWWQt8RvxJj48xthC
mJgPiSLqawQS3vltS5dg7BZ9MTcLeZTJtUw8+qLAtYPpC/QcMalJpfCl7YrTGqr+
BVib/VtKs7BRtc1VWnSgWIfqyogC5at1et9ss+ONy4vZ0f/oF+OXZ9/XtqR21deB
VZ+Vjqbi1U4r35OTUeKY/KFQuI4I+hsiYN+BScfwoE+dF/85xWiRtMUb8AdTf43q
2kGHPzxZa8YiNA1srr0HTvQOwRr30TlTiEYgdhPmFsaNB1M0FJW3qZLIpDlLNu7z
0ue075prNJlHPJZ+ZFOCztE7UjBd4HwUy4kVVc7h+aC04K94JZT8y/qCAT4Y6JlR
kHoOVe2mVAUfStQuHw+2xPnPyMiELdZ5Wynzzf+PJn1FzgZya8LGSY0Dg9haRhNj
K64z0/QlHUp6ylNQB663F53WhiXFsct1hBeRNLarfdHF9LYrv+gzDuNZ5V7TeLI7
rh080vIHQFByjDonfkJsAUnnzZQsKB0DPSxiNWsqFXaIehlSF3ZwVUsTV5dx/foT
sEOx8dTScGN7XHZdmQIlfY39vXAbGyfSsijb32pUXX2mJ+UoJY743RgglTNL3ERg
vEGwABBNpxvqzNUKJxmE6d2oBzywrB7swaTCpBmqXs4nZvYfQlph/7EnPDqmslc5
FFFNTir+k4V6v0oqlGVRiDgRwp2Wvydb5XNz1VOPWfGBJaimFgXk+FhmbgG8ZJt+
eTWviQ20x99nNOb74c8hK/+4YOqO5xBLzuOyRu7+wunW6INfz7g31vWeYKo97ib0
bU/QtffLfZ81pxE//I4mi08kON5PxaxkjZ/Loz/jMly4GgpUaXpJYMB+QPHxEKYQ
pwTM+AfhAyb8co8zWtJCFDhJmq3RxvPyK7x3MjgZq+Fu86axjD3xviligJ451xLx
aqKiFcSe6E1H7lok3M0Zebam1SwWWsPMYR1qgrXGRo/aoL1I/phpT0AGU62hvliv
B6smkYdVEEnnr4t5M413N/TrJq0AUYFLcmR7COfCsoTviNx/d7z31ELPJ1GRrfJ0
FqGGutXLM4W86O98Xu/+vC5tmSbSPzLp8sHFlm4FSSSzo93DnEFHotoI8lke5w7u
yY9lz0vECpfzS874k6o6OMEMDQEOEBokveaV0b3en4o9r3sAhojvj0I11gij6aYp
l4D8gnVN0L7A/AOyx4992CQaxrdzpy4vrUrmhTeF5hlTVqqg07/G5yXG4WSdLBLB
4oEz/kazSsAnKgWQOwT6kWyjWbHyCbSQkiKJFXzCQx5vYZd5yp8QS2IV03QeNBWd
1jsgfAXGcQpK95twYF6IIpvyttuunlQoDRzqXSJHTR6O+XTfZQkr0e4xjdoGYRay
hBV/EXQ3jZfvkQLckMyRd8FTSPQZYN5EvXzGniRBep5IB1ojywPhdgfRM6tvjOWd
EXLcIhPRcRdedEeamcoK5JLMxNd2gibOJjGP/MhrO4nyugfjE0fwVm5qfCDM5S0U
O+1jB5NqpMVhW4DJLp660hTlGpc4u1APFlS8vi6qIjx2CJRoUJJnNI5mq2nwa+jz
FNLTjdOxSCLj3gZA6FchSZzzR4RF+vjKGLR5sV+uep06DaLZliZf4EK05JHAnE1I
uzxtQO6NKsypBUqnGYdcyDE/YJu1rbb5Oy6kp7wTkWCMIvJIJy/bK4bqahimJu8G
pgGi6lbl8hdIXRUVzgsCll9s+J8eH2ZJ+82y29GKKcKTfV+k3YMs7InQSMUi5yYd
jcmPYlmhzanTRUV2H0GewrspyR6NxyVqrD8N/6V7GZWi+f6wX6rfeYAcpvFHoalL
X8arlXM60xy1v5osP/NUKP95Tg+dD/JYrGmXb6Yw/7EXLO1YG0BcGW9Hqg27ycaH
Q+hgKjddSH51krwkvM/4c80BFUaVBQ6w4YZ2FWHUDZ4JSyszLB7/86gx6t1XjEwZ
AEOOicUlDzLqZcFuPqU6SCRnO9jWsQrz6fc40Pyi347v6Gehd3zbTJIEcQgmXSEk
pkt1DYNHQfcEk0CmJ5sLNhHhGrmXAzrIyroknY6fn+RiI669QhP6VYDHvggWPKJJ
8L2aF7EIDV8c6UcVSwXh8LhxPj3b6zmkfFTn1KBMVcWT/v01Io9bgFtxIZFGNjXy
Zeu7oTaERI6eE+lvn2Qdm/QHybV1SyAMC7MxtSgbPIv9Y5eH+6IYlsB16s20CRxi
l4oGl32830Qtco+MIprZC98SjVjqg8OXLyVT28tc/WUQfCaoVE/QgZPTNbgVZLij
31bmpB5o7nCYZ6uW1NfUTI+6cx7XirGRhZMFUmBKj2xhyM0ScUM1uOl6MSTO1w8D
jFidaA8WYNh+XAXSZpBeSP0l/clzhff8kuVAfR0qmbN/efT7qi79+WqU00E8Kton
WjdKdWz4kCMYAUdk4STWwbwIcFzmhI2e9Ijp7sBV+wFVyMbpruCKo7OQ4FVbuxOe
ZTBZ2yGcHn8cEeCr3u1Zt87mZOKPe8SFEdqV/glbH59sr7B5D7WMkzni9RN+2GX8
z2Zmvo5+4xCBu5qZsU7LJCzRd0Ml073XpYCmURCpUDicu9EQ2HQqiaUJXmeBuEos
OpfMMdIXZFwHbVODe4y/Emxj8dl6S2RrIT0s3duBMGh1gWvSG7mSYlFN8w1T78Io
/PeVCeulsZgaqPNweTcJAbf8W1gJblJEs6f+P2RPYppmVpOjwXwLS23XFy/+5ScM
Uq7BVej/Vhd/oNS3RV5fplA9+hQ3qiRpD0r8B7r7mZAt3E7+nW2UXRiFf/tShEkA
ZMumwo8HAxzX+0LEgBS3Zf4XPFwuYN50g8nLBV11Hc9XE9SsQtEYCZ9LZKS7vQkV
BRIBTGnRdrN3PXN1BJ75ckZ1JmERy1tuSiGoJH0hh6MRIFm/YuJB+Q7f/wICDSbg
Z9OXKSEju4fGeDnIh0ZUYvRwjYIN8ihsjCSIkNPXYkzBhsVlfV1HMpIT1/MOk/sp
pKZZKbmaI1713hD1t87/IezeCXjBqgc0UURWS1V3W+AHyU3WCoiUKzQIGqK0/Fte
FW6hrexbCO1aJE2+zznCOEUFCafr0/9qR4RUcUNu3JKDxr4pJ8AdfdPqUB2bi7FA
dSYZ5czv9meF46fe5f103huSSD8IE5vVrQv0Jtjdw5WsNp6a7pgXppZjdrY4u7TM
v4oq4SGRfAkgfl6RKHjNJE+Zg0YyhlpfvJOlzEkyl58APYqu9AMmxZ5faSL/KhmZ
YzmDrxfDDiJORcERf4dN8lWUhRoBeZWz443SGMW9BItPg2TOEWSqXjeFiv+tLILc
VF2LqK8HuXJIk6S9Yno4egENBJprvDVkEaRj3tvqsF3iQzzhiiw03hwOoWo9EWpi
t/FtziseuJPtli3BlTPFhJd2ZVKOaSDf/N0svAIRnID02LesuwP5pKE0LdjrzJ9Z
Ewlso5oAbY9Fq9zeN1xBeOk678F67oYgcVrTv3DY8OS1MqG2j/iE4pX1CXNij49C
OKtrIDqGvONU3EnM9S6XEjomLPB7xDLCqnbmH2HgC3FP5mt9pyQO3+gk/9yk1+UN
sf7o4TqEomM5cCI7rhSALZnbm7ALOScbX9baZURxrjPkNlTALctBKacswFi8N8aE
hN4R/WNuhc9RcfZn/kC2zGLXtH4vGEY0HfWYOmoaC27Jf2HbV3Lgb7XBu8t3r+I1
VeTUTzluel5IidOjJcpl7aU6I0jWUKYzsHaXTCyl1/qJMP5lbxZRMTGe4czE6cTi
/5ESR5bR3+PqO+90eiwMiUSAI1tYkisuDqHOuYhO2ma1EccDeM9SXUKcQzdCRhZC
FewKbCn6mzWb/uJdmxerYcJ+fhPJdjT+BSKL7ldn97Bkr3IsTpP/RtjPSRLUiuSO
ceWQHZ9tue6toO2b1Di0bYQnoUKu/5TVr+sTsoAG8JD2fmhK2BbVWzfOuz81Kd/T
LxS0W9LqM0a87gvb0Z242k9sXjbJps6S0B0hKalWErtO0nD1HtWRTUDaI8vT0IuP
5VBGcZ+8dnPYC04pWHRRoVW0ye7Xn+aSSQDQZfdTubEcep+KC7yebNQAu/NwYk9W
m/2+191R37FKHSviwSQ/UOef+aIeol8KnJS/pmS0WsQHFS8/YjjZgx79xEMkSndi
kGrXDHPudbIas1s/DjDSG7dxCKZKpiGmHMqaJz6qDeoh4E8kGf/VPnrXsdUh3u0Y
0jpuGXfvDzgSBlLdtzWUEfbjxMxGtVnL23c5P5CHFeIgDQGC/LwO1FUCI8Av6q28
BcaTFsDzCe8x3uHfZtAxWKX4MW5UBy/E7sdHVa8Yb3qwoVrQMfDjMkGjMKdko3yT
H17r3iPCGV9ucGfNLQN0mQA4yGbH68bUtCfQN457feQMXyGz44beSUPGSQyfFWbv
Q4tMNkIY+AYRfF3xpJyTkULh51O6mip67xNGspv01oebdxsRqDHOutC9nrEgM7U8
EUzbRAwqwLPZ/40e4R8/UoaDPos4XR5r8LalyRFXMI4xeOnrR5G//Aj6O/u0KMWV
7ZhLNx/5MSQhMnM2KpW4ipUyBMjSpcaosTJTfhEl1U5WOlnBSohdtHfTjHY9M+xo
wmqKrNZFFgxZZiOVo3iLyOYNpqGWHEKbbuObqFh+QNKWA3LNPQLQZS2FMelaVgBL
UWVBfqesAJShQM2R3EGp/H4jkW0uWDN1Irv8VCX43sxWzTf1xxqawYKxQa6CncHZ
ibwdat966YDE0CxnuBb4wbIGotBdtNfETcgNuuucPDDHsmAzONg4v3hgUQiZTANt
wlHx0yD9rnbQN0miUb2Ip6+50gSvAvdwed03gLhsIDA9cHnNM+uTlOZYHcKPHS6Y
9I7vu9EFcYqt+Is9MP4UxiWnv4RDghGcf/vYYUK+htElBnehPTlJUqBMFNTzCF7P
4nssaCTgCuxXUgp0+YDNHk+5hY7OaBC4JV7dwYpXcB8wOiFi7ewQlPKsxyFm1AH+
crKg3z1fbOHp+vaq24zMFiPg2N2vKYShz6NqT8MMal9t8cYMIPUmMNQXfqvMQ1US
fgSrcnl9EeRrMAUuWiXLoGLFYMZqh0JoUwJka/ETDSv7kKGF72y3Zndm2WNRIwZe
RsUI+r7Yn/sde89XrMvgXFygsUdhNqyWIKm9A3erdgGiPhTQSSelRQ2GVolO0y1W
PTMNrQw5OX9C9poCxKG4kyjfOHTV8Vg18XENW94GYTsA/QbfTbzX0vt1kRaBp5el
58CR6oDR+zEDTCSm8RDLakcp8c1AFi7XCl5fq/0br3Sw5wjNMUVmhhwWKr910E2r
5DKxB2QCc6rVFSAd22hSjzZ6t7Z8+i3c3Ws0GzWAfXNQVSEoZa5NmYibHmhRkics
gajPyjcQQQWdM83mNq7ELU6Ru3NgezsyY/992K0masNyt5Uenu9V7A4Tzj22igNo
71bieeYYmvfBSb+9v7SCYLUbL9K0loDO0pCTLeBHLWuh/oyWr4r0TlmCCBBxKcnx
6KklV79/ZlL+rNgaNkvw7e5d4qsBzuepiNZt9tIPgNX2sqkTkuAzfyQ0HfOHieQP
RNnyaw1OcYX/8WmLf/6bq7doocvniLrQ07rku3mVhs46r9/63SuujUdpcnz914KG
6idXesi/O425gGMjOO4Ica0g0JskbVgrde8TvUv4jTMTcvMZ16MplUKapctl8bgL
vPXY5fIwr+7mijxk8++JIa4RtRGOobfrbO9wBiBlcDvHo+frfr70BwAXwG2BRAKy
dn/82F52azJOlD6I4O4TogWPtgUaL+cnKZXje6SsmVNCmjbuIyXN9ZbCKm/UstAA
AI1kA4Ey53PSBTSuK4B/QYgfYGpjfLz4CZKlM4GkdjBfQRoq3f3T16AmQL29RC0c
eFHurra23+euxPCghj2vG71XsNm9og04RM0jcyKYpNkNRCS7oAP0vCiTTes+vUT9
znplQnLf8KSk33ylI79rlOcxNsVsIHG2n2u284zA4w4OHfhE5Ay6ziDpXmuoP2Wj
RsBmmnV7GlZXDktj6tuv2c85fw7eRlBZbvhDbXoGtwa2v6oYq0rsOjYWsLzc0T1u
mHFqMrNc0Z2AGlSl1bKbwkiYyw453U1zp9Dw8uR6wT7av8S4ozilsKglpcU1fGCc
OeMnI1TROoTAJAcdNYuQtkq8vj1gX/BHq7wH973TESuPK7MKN6RKB7JSqMhMSg8i
ozY766l4CSemc6lcGTFCqnK3bDYS6dPWMBvDMaToJcpl9R+nW71JYHVWyJxE9/Hl
FGqbdETg4MZ60l+wuDzqFU3eFOAMfj+ymGG2phX2HLH7kJSvwAOiWX7s2tdSLcH7
a+WnU4IM4pSweErmynGHXyOS2UW5mAPRsowbMNCA8FdreApMRTTzjjETkzp6yunp
l5EEiVI2mmim+HFAl9pwTsdjd1na0YA5GMt+EwF+/rxmQtdnG2idq3EoNQJXhdl+
DVjP7p5KKiDeVxAR4cO+ZS9/bj6sWYSawVhxwa8GvdUJ04MenEEGanjRn+b/fPCV
6tKB1dJfTXm4T6WIdh54BgQ4vbaiZDVDPVAXbJ2bm4EJlpdbKCSSsY2houhdH7gH
0WznkMWYxPFIjeZ5gltyJ3KNjX7OlqbbNbuVf1qhCkTuP4adFc3ZxiR80Rc875iZ
fwq07V5J4a7X+JhLQfB+kW5oZION4+FedsJryD3GCb9+RxgVuIfvwmW2g7ujCA8/
Y0aQDK82XmFFRuKpDMU0vcO3iOv98b8T82oQNGJZBbh9XN29E1H7x2FdNtvuCzsY
xQ9mr7/xD39ICyB9xO87psqEWqUIKSVYsqWTyJ+wepvTzwlrbZoqPRgD466RRveD
kqETUVFI+JMWWIuefaGxxj3FVSX7gMihb1/GOMCNvsphA+VtVN+b5yafmDY4wS23
905S8iTyj3TbchKUlSQeBTe9IkRIoEvT5yHSPqQRyZeNX8CG7CKR7oFTKNVu9W//
wJvYm4gIBBB6W3uQHY1C6aHLq93Ql/4nCkXHkoklkCJuOrNJLdZUz7ZwSgUEpYcc
T+Y+wSWXkJ535/vqjk377g0uLIJS+74YUQEYOwn+QQjDJFeHgEsK5/YaLRkk7/E0
9xtr8BGySkl074dsYBjO3n7EWRNT16FaYLV6gkq3jmTaEHxopeUWvw2WxHLVcau+
HDrgJu+kpkSUyNYqArnD0Acl0+CU+P3/EULuwlACq6DXhrpvsWOxCMAf4S1HeS99
9iTuqbqPKdxZYQcKbOEYpQWWR9AC5BaqBIlPj/21rqfIx3yYCH88Y+nSrfJpi5H4
SCCrb9kzUdG0MYQMc6TIDoTeRkZJhbb0z+1uwlLGkhFjlMAiXA5jZ+Pax68X7ZqR
ikzzKn0K8dDUHjPjQXPkvb2xIhOXhpMZHbYv1+lY+za73ur3suU8c6jn6+qfW6aH
Zm6k24r77kxoHWWdwZGKLwhHgvE4ZRmpbbElgJURqlr4SLZ0Qht9Iyd4i1fIQ6HV
sZA7oMZdhPG1bSblnfS91XdGzgxcJv/fIKmRXfwD+L0sNBOXdmaY/hxoC8sGJ9Y9
izC+QTTxdNgj1Au55+9jT0uI2aSsgz5wiTgfhHnHTkAZP2OZ3BaO05NlQZtgFcTP
/V57FunECLPsh021gATxSqnp0n44AezLrR+NuEpn50+xjt4L5T9HCqWiWuy94ALM
6JX44NvKFIXFfaf5vFmpxLzouh1xgXbhOxl7S8dlxomb78s9zJy8MMPQNdfVVoJo
eW34EMhgZdxdZEzWXtmwp42dNl1QpJJIWao2d2ys6KwD1OzJV69bZdsGUKcW+cgf
juY3VAluJ+gKC6ZAxBNiVzhCqwwsCiee2d0pkX1Q/lII+6xq5jpkju+vGQJoNqQg
RiFQuZ41VnQzOjqIvq6nlfNv2oqdVsxcCf2/55P1ZoSqgk8smEg4qG5by6DjX19j
9o7sGryw3N9jjp5ZrMvAWFrVizars1U2KpBkjDwVWCGOyWRla1PEOFfbzusJjiCr
7bcq0Ko8qn/UJ1Qwj7nq+4/rW/wY3/yfKDEXgIrCyEpTcmYojWfU4v3P6PhcwQwI
0cLvjsGgK/RUa1DfAV++1Y7VwrTgGTmt1rhH27N3i8m6VtJV+5NxuRR9r/q05auu
CWaw9FU/p64O4mN5e7KWVA3wJNO507XrUJKmMu6nMHjv5MFlh+LCNa/YlG6f2nwZ
rL2lmqGYdS8Kd33ANVCkZqt+iofkPu1ReQ6C+dXdOyEkvo5dp80bQtQ8lG1CC6SO
GFxyFQgviEnir9KgT6bUgkI7sGLHCcDQPrfcbLCZ6HjITFvPpTd6izIrYi5ssM8j
/b27mbbgUHTrKtIl+5G6OBUtRTMbtswTH7EvbRQKjXIeO3BrG/dxOkJOUTOu6zpQ
suF51QRnUYY1cNj6CfMSlnXCrTL74pnr/uf2ctY7dmHDbyqomzHT8nMb6w+839O8
+2/+kE+13wOvlNh8m6WxjLt65dC+uOZgTRBJfnzUm9kvu92IdaC7WEEdEiFlJXvr
4ysV+Bl0wl7pkb0KSi475v+BRyf4HyEA4PKXxKMMDBpi5gEXI77GzZRx1TmhiBaI
BwvzrlQcWKWqpvMdvgoAJ3FpOfPfPTMqf8S/7bhH6pAFk4wR5WCES7uA4/Z4hAne
OZyXEzaf8jWhvDz1ZFnWgQpsE8CaZgjNbJbdAXBYOsozfp7Wwx92cEUqchzwglPd
2UvqIvIETIP+YVRH6G4uv+ayOdItLJ3X7zWW0n4eUxOmshd4bkDZPNxUGjdHYjnC
DW1ThHWCz40r3BukmWsk1dNI+TiuAFSFJdter0pPQpJZU8Jmve/jtG3QkvYRkAq9
vsKVIXMS6hXeYik1MZdDrafJ6qrnP96bUSdvcPBcj6jLDt0IQTzhQhopZFW1SKfV
DRWNollc+GHV3USYjh+8e8U9twpN19oiF9SyQ2bmIBgH6i+6pQAC4FcbmgedQJNy
BJeTDbNENo8tdOMZIKEDENVVC5tr435XV5WMi0fHm85YbElxYiySHGzo+oX0vS/C
leUvuLbv5jTh9UFwjWgDwWmyZ1KE02oO7EJB3vCI0Gx5tn1EICDUJqbQ1Ldx6ueM
fAcetyvy3Vmilo4qgYYXoVxSJF0k1kAIBvYr+QJKm2kxgERyUwwRDv0h26Or16UU
T3JCedkodiO8cLZ9jRaKO15uFLxRLCJCFlRV8Hrdw46RtpLELAFTSYwqvUZgWTeD
bRfNmAfLh2BdOF1hxpWkVxHw5LV/fc3aSgXt9pQ0zd3ji1i3sUAdIiMbH6T7X6Bb
urBkzD9/n+NxEcNDMCXUcd26Zij1CmJFqtX3N9EBHtW8nvqCUoh81F/9rHeFjfcg
kU9EiOZIb/a0/9vhXYE/UuNQehlXiZ2Gs1oiz29Y71nEJNbYRkwsiGGa1N2l0K+I
OopU1URWCtWFbnvVrQg+iFzJ9Y4V76ldhD6tY+rYlc4OP0/AX3lmdgNdJnYN2cbE
ZCC8aJkZtzzIflw3hC2GeKG4OhkpHNlnlHAMMdezUGMBQwKSuhUcytVrCAPk/HNU
YYRXGBaGWKxT4M9kkXc4Q2duKY5YiHXd77aHrGPpJm0FXeI3ZiK0HRE2Z73FrkXf
7LsoDvjJL683D7yaprqYEDTZVa2Wy8jkhSY3gfEtoOlFJIxenKkUCIrIXWnGr7qb
HkF3LDKuqplKVyWs7Ct8NHq9CT4LBDrPEGdhQqRnI5JGNfRMe0HGCwP2ZMSJFN/o
j5K/JlkAaw9KuVRKPyk4pJJEKqPcYSxTZrXiQrHx0haw1Sn1IEuS9JpB8/HFlrv7
C6mr1nqqA/U12CguRj+kp7blhvwYTjnFHaqLIJOUhu2fnycKpfMTz2Fv52HqZlsg
KIPuslzAHYMsi0HkPFYsn9QX4I5TCXsH9e4uOWIFdc7JstF/lqzOH8qIOf7bwZ+p
+bp22/9hWo8dA6hvwpPyST90dtFd+ELc/y4YRNakcVEIU6kG9P5Td9zHuCLHwtuS
Oo1uC25j5OvkfSyxnFVoPG3c9XhAnGYeVCslZlicsA9EiVAdJVwWgeaDLu14LzQ4
JPQzVBHI0s/kjko8PTfIIPfe6H6QBdXu9Di1wB6xJGJskxbfxL0TE8yEFIElvHUR
oCeBuvUc9a3XXsYubCX16OGPeSttBNL5wdr9ld+feX32sVdsnpzg1Tpq3wRSM/7R
cowX3b1KOGvMYuOf/nxnOvaRZ5cRCq+bfWdmbfoJxQo1qfuVxXmET3SzpYJc8ZNy
1XzU6HDOpoGFWBA2NHP3FI1zBYK+YdgF/crfWO0Iwuvsb4kCb2uiLE50xjsCozc0
+xhWvqhqc0Pu6G3EVhkE2cb0GVgHRQaOJJz9ko5AffQ+DWNPAAzSZ4G6OWBqqUkv
n8LZlCw/p1u8qHI3XFMfz2lpsz7cRXhJUEb/vqyYYLr7EQlZ24uo0j5ZcEV7xDBt
YNd0Z/ux/HKQqxF9O5As064d5rTr8d9byTH692rpVNihP/vmhiPk05pieXZJ7IjW
p6Xu6SZ8ZUmp2K4seG4f3aQYm6jtsn/xEJw86jqEKNOt6t5oj6iZC6xiOiLLj15z
dvRR6cYzg31IdH001k6lxqsweu8tB7rvJLEqxB7lm37Wy91j5zEhlB1w6lMlKyeT
NEE1L9O8/E4M0MVAmaGZ1yOHZLD04s0DM8rHjvJG4QHGO+PfQv0z5RN+WKgssbcF
wXwRzNAs/eoVpA2tZDYLM+tW+424ajUkeXciwf89aA1s/cyBX2QtgwrvThu8+2jW
yXR59NCBVmzXACE8MuKROQbcmzscn1WO6zMNBQDJGbMfqU+JSrTZJmJ3iu9EFwKG
gvy32qOgCOtw06zeZU9GlJoi0lnItmbapsxPTpt/BN8s7/Sxw01zCoTs8Ld0XMlh
owdRi5fPeb1kGEHQ2WTABhQgVEaJ5gT8oh1Kdtr+kAbSWzeTsK1lFwaki/8txUfu
vW0RLIa4ZVRC13oD0B12ywjRZhM/OqK1EgwAmoOdcDfC1lGksoQ7j4ai+mBcUizm
T3YCOVeepeWoqp9fOZTYgaqXg5VQtem/a/qbEqNDgy3cmB7ylqQ/wtKYxSJcpD/G
t8OD+1lH1E3wjbtJlJco5JbFxRDthhYZx0u1iFD7hmcYjuLXygMfrcWLQqGeBwfD
28Xs7W0E9pfMEcg2U5I4g5622GJVJVwwkXA3TY21pyFoz+cRzDj7HL5BjlrSO1EK
cg9VrTqaR2bORO8P9wmGvg/Nfub9hPa6t1by/bZbs+u4tPabrJ9FmwRQUOtf8tNL
7wMMgvnM2tBouUb7pW8dSYWPrAG2btjO9mvevmsHIL3ADhBP8qygqntQe+/7aYQd
uo33HywLPfCbdXdHu2iN1pa0czyJ34T/rl8tJetEXsdhtKs0XwCNdTG4JG6x5gf7
LotBDYMN8DSpBgOu+6+hVE7EIBes67BKdtJa6jEP5kk/df/NZT1eN6FiVVGLjtdK
rZMHF8OwusyKUHU8nktrodeuwYRqXoPdvSy0fwHc8mXpmB02vqZJo7qpet27o5gz
yeVQ9wkJ5Mmm+HP+k0wI/TuO7il+CF6M/ALtDhgTdBdfxAUtltHFxQsQBh/Eqiy8
e3Dz08ogy/GrvfUKCz8jysPVgYOYeYMC5xWgCRlOFZmw+zk2EXFr96lmcyVo42NE
5vsHWQuBb8ZWXf4fikYZAU9Cdt0ZM4CVVT7Iqy2/2gFXZG8dszIeXb/rM1LzR5SW
s81pZNfy0MdL+M04x9lLwZZmDocjBBBVTnv5mLdj1pXUcHMuUYWK/ZVUXBZ7CzcA
tnhA020Y9IMbQLx+rdc16clPjF73Ax2DfiOpDjWW1BSswERkF4GnoQTWko/o/u+0
mhKIKuJHxphecwnPXWaXo6BhhT2mTceammTB3Wxgvs87iQulVrTgxCY/MgVl38Bn
511t4IvKsCSsdeWumWVC5CQ4m+9ZpnBoLshk3h0w4bY2ZhAwxFpKYWMi0rOJYSXo
oakfQgHoJxrkP7yLQAo31KcPZTA8KsruW0ZMi18FNENCD1Fx/3e3VJDPhmF5OfvQ
ZMa+UKLhy+3g2wdAr21LfcQEdiamgZhc/g1ANjTg/xoIBlnWNXHK5tPbK48l1oio
NJ1Rg2JVZAKyU9nwgxDb3cNGAk5Gsh2yMpN83bqkDlHC5bcFg8phx2M0tr5pkbNA
XWJcbgnD/7OH1vMoL59nNVKPiR8qMUYiEyB5p+l7N6wJ4Nd6Mkll+4SUOWQpu7eh
b0tOzji19fP5MSgC029xd0nd7pVjqWX8yMZB6wtPaETpbY3MZzFv1IwFQ09y6Z3m
vwDG9qClVGgHvI7qzeenJqGvHVOjxEqqX+js1LZvTZZ+qdFkUmx5jsNmjMvVJGN/
cPFpP71oJwZ1rycUSrWG6/UlFJzChDGF4kdohoaBOH9jkTzUH6pUjFH7dCxwblFj
nwPGHk6XHADa3ixSSPzwq9CePBBSAUNMXqye61fhVcNyLD32uQDi2QDMa0qkPJnM
2aFPfnoa6PO2aLNPm75bv/goXoVG0U4kH5dF+/whor6BZwLqZwb1USLL8GdmyJ33
ZQB9XPP9OsysahUi7wunI879zLVxlbvwc+Syw5g03mTrwCAh1HxeQ7v0fMuY/TIN
aUU+tv3ms+IpnHe4KEO81k/c9ntrY3fmbWiHsa7+6UMPQpbCWxkHnXG3isoF+Zqp
co0TALwSs/zQaDt6SHToxWVP14H/uYAb3+7+jCGDeqYAmA6OjlQqzRGyjoernFmT
f/UCOyKQdTyue3eCX2qZJ2mwjM7nODt9CnGCX1tnAnrnJv4PpyBcG4sjKk9hI7HW
NH+IVrCz+gg7QuzAlu+tv1938ByygdlbNNNf+rqtSFvS2+V8rZFX6pdL012gl/JY
/E31FWxTmmW6+DeCEW4Fa4GHnDSTVI0YksJ9MXGuZ+Fjw687hBpmLa84hiOMGqxU
evQzBpAX+vBQhiDnJbVPxA0Rs/F7gZXjXmT24ND8e2RnQtK7J12v7r49hikpTu7L
S/mQRUu5hp0Gpkdvz1xSGiE/VbjjL3w4vdE8d+9fLMXQDRBceDCjVTzP3nk/sgsU
E19J8oTa/eDiIJbwWNsqM4UAtwsdB3swf26wx2hi1pFg83hSUew7HCYXWZJ99ZVI
dBDpd9mimLEdoxbCnxE7CUd6vfXBzwdwdssS7b3j70uaulHPUKlcPr899fl1aKWN
21Qn5Y+0+iG8I5HdiP3/GxwozXJ5+4dk7kbfnNSok41TexEZXozp59duNT/eIjl2
b7BBBfNOMaJu2c/ZjTqP115VuLGGeBzLbq70og6tDjv692OimzDIQxXjL6hw/AO2
zR8xVYTCJnjzb66z9x5WTbAFVC/WPyM3lw+2IG2ehNh31rcwAJ4cIZsnWXtbsaOU
cpr4ga9M9nh3i0FvOxXbq5mmufhlpqCTA1Aw8cP5aTj9GhTE4uILJgJOoV18rRZG
fX/epoanIR/UemmE8NS3UGbO8FbLFw07OiEBJpVbMiJLzoHgEEhG9v4zpE2b+kfj
CHbKBmg76PRti1yyV6x5S8P2d6FUvG0PNQaW5pc2vq6meELn8MZNSq4t8RCbfuov
2OcoWHrAOa2AIZSJqh/n9ofv1tkJ1SejGJlZsLmH45+rJfTzYznhposo5ikzpQLx
eZdVGSo4XR0h+/JyTG43dCa303g/S5NfFRGTYl7nvmILXarWbD3Mo2/mx61GwGeD
CUBQBKZl8M4h6dfdZxgQW722oXYRaI0FdbPVpmuBONyAc1ePrMPhnhtq6AdcsWWx
R89vv607eYRzPkYvJQuhYan9vswUy4mTmrkc87Qkvx7iJGbNfBzwhpE+2kHmC/VO
DP1SbedeoPy+ybSzOhFZtdlpa3Mf7OPw9qjFFQCjpmAVuHxmfKDGRz0RQSVROJOK
agYE7WO+kP++w2QapJxp2uu0TNu3Xcvbs3uCz/tb2Syk2JG7yTC0SqF0r9GfcZMo
Tu/DXcdZ8I1fJQ/jeZBguVr/YSeasAwDEVLGPj2kXkIWCux7DmbfEbDGrzpjYfwm
F2LVazU2xUDJlhBahzlioH3isQLMUWZP1L+RYfBGZuJAN0mH7ylKSON5jmTp9WBz
6ovfLCEq7lKuwDm7XVsjAUO7ngfR3eDW4upAwP5+kvcND3aFW8ap1lDud07QoZuQ
2FG7b+DtKgcsTekdzXPfbuiA6CSSlZBAF2fhI+Ir27FF+zLukb4OTz9RgF8K+JMw
mY5ZnZwQ+HTVNrIZtQbsGy96HkqVAKJK0lWFna3r6Kj6FVYlXvQQ20fCLWmKuWAR
H9QG7DlpNJWe/AC6mpBNkIrwy07yl5yHlicLzlHcUXv2Qw/doG12gSo8Ngu+QGjD
9yZPgWNwVTAhNv/F8g1RtMV/WwPpoTL5AwBdHr1hHRIY9k4G6D0JblZfUOhLkurG
Cw0BBjNoG8wgTqyUS62vwTUbRACIBuEbZwzz0xH7YRwHtPrJrXiEvjf8Yw7jZ9Vb
GYeepRepg839L3xi1VTYWTzqJhT1MQaJQnj2iQG1SBCrCBGVEzvpOxDLJM1e205p
YzKK9nz75jcViuPseJveR90sGqQPMUAFKuYjfXusC5RAJojrnl7FBkd7C7QnUdv9
62BQTVWnZHdeTZRNTndpzehBnip74EaZQUWMSIcg0O6MWJbBYSUb87ajtA4lLg0s
FTTJjRYHBitP0zd6p1ujaiSMsPtH7kPDqxLQ6TUT38xZwRxkRFcSFqKswi8Wbrw7
jni936H59zgBB9OUWm0AoW0YYO7kDj8wT77e/0HTkGBlr8WEfn3iEbrAj+/KlvEU
mQVa0o1z/CtkCah8syEmK6X1eXbyTL1M3LeJ1WKuwhWHC+4kgiE8BQ7numRZ8LXA
pf/lnG/EzAcOfcqBqd9MH8buoSJ5n6mGd4L77qIS+0SvUoQ9cR8EiA7LKbOBx7fF
AEGYHkDe5BcVQ2xtGGS3NIBsoXc1Ll+YRaUwQyuPPC1scvK9kfPjuAuX/edrW3jp
1BbMATo3eyL1M0xCddN9Bw/1LscW/NcV1d331vvrd/iJlttTjfdaadUhtnyt1ZOC
eGDsCS4yn+nOispzN6OHpdbtlCmoXE2ObNpcrAFayQOz8sSDxC7or4YcdkH9fi6G
Q277MCtC+l4fvPCpnlG9C0l48nPE+XI83qg/klh0MKxyhegtbm86GI6DlNREtlH/
ZWTknn1s3pSK8a3/WptHYwxJxUQX5CitO/ht86Jb1WEmomDDmqczwsTaifHoeSFG
vZrBamPsLmd+mTFWnbJ/5m+eJIkr67uGHCJaXp1METmvaI1SvbqvxSORCwDmyOWD
m2+QVAKaYwGnWvckmpyaY7WN9ZaLnx6JSFL8vhOdKBaRhugDDEAqwef/B1LIx/2l
r4FwT64iYjofY5PPYt2gSMzmVZvLHF61fUj++IJCTPwkm37lrYAu8NLsgm3HULGU
FnoQcwz2V0rQjWrp1O/NHk936ny+K1zVIQYAxZeajXYfhqBDgGlc8Vsk36BCv+tP
YhRmKpo9R7r45ORMNleQJi9mAYDW8p2r0giAzhmXkbONfBhUjD2nLAiADWI1uxMN
2OT6yexMujtPgNGj2AWWfOyMrgG8qoUt2vd4eKWthzKUrw4Su43+HDIRC2RG4pyr
eM38D0m5qTFPFBjPCmh1lzFIZ4Y7Mmkt7NJrifXtsN/9Ut01K6XL4BsnT2AE+u3X
fuyfzjC3cwM2VE4X5Ncn5G24H0AVSFUEY3iZjm4R7oSlbN3uQAniaW9hWm7OenBR
ErDsLQAUlXoe24Kwou430LmTU3S0QWbSk7ERd1QPI1a45HDg/BZCRuoDVeQbFlt6
WbXgAwWQIYApvh8Tsyzp9lx0QCFfY+Lvqpx7gjV8B200pDlOvlCbD1vXCZHU/ZkE
hcf3Rq3xaR27siaFxEu84DnK7037kl6vIS7a/UO3DNHa6dnc9K1ZKjq4iusXge5q
fHVdkVyiCkBNpqReUZiFqBeJ5La3qrloE3N6je1pkR6Xw7raOpZIddYyfspqKcdm
PNtZqKCMKhf9TEWQsOeNIaUFaL75dvB7zrtmNWyS+a2tV0T9a9NG68pn6QR11lfF
wjs5JzTGbxVPyxx0VZOcnRiI+D4x1X5dboy1kOzmsIH2g8N+GNe7vc9iYQVH/4oD
34omC+DPeklse+suBpLOPqHgjXI1EtO8/XmRLN6qNa/6sWzg9OlP1LbUQ8Qf2x7O
m7crLclbUGw3HjsrldFCDg/6suBLbC6cU1hGWQEjJQxz44io1381ES/GOESTnOmG
SC4TMb8QIKhplsSj0SlnLW0iC5tw/sFzJ1jsA+EKG8RgS8CSR+EB2R3zo0C6P2Jr
W+Taf9w6BY+AihR+48ciX/d24c+0//bkLdp/yDKlSl4k2tStC0sknl3mlz4PBYA1
I0RONkPN1bJZhL7r26CvU9avYTZhTDSRiszHhHM9HURg1Lf6gIzW075huPhWdWiy
XYOa4ABvt+dhtDeVMB/CwF3e7wBDPjhoR0jJc01Ew3IN3sjC3UhBmm1jLpbcsK9t
aCPI1nTT9Gk23T8EdJZO+PX4ilX3/Bz94noDURYsxNweviH7rVcePboRaq2YhVjK
riPrOvnTIS3AD4JzgzKmxTrG5N2ytmYxBPkzPjJaUptJyuju3yzRsDUl+LpKNMA1
SX+f/17QplFQhqDRpLPc+tnau9a4w7xhq6q0mcMfZ9hDvm9gz7hj+fzvB8agkvkn
URcPqnr410ftFgH7niChMUVNUTywNzWZbeJOtysI7oZ7INxFGfOaQGXjeh7smYcB
PJl+4UFyfFPluWzeC4WKEE9ge6C/m7K/ic/y/1O954Lrd8am1HwM93cPJ9sA28nF
o/tQDs+EOeKyHJBF78ZAAMSEET6Pocn/wwoEczdc3Lytb8A/TYt3MVbMnkDwAxZ6
egxIOBTIyCd8lYvl+RSW0/935TdHHuSG4Oc26rBFPqpn41IHoqsEPKUxIPzRkMQb
TDDpTuiZQiwdQZNkITsl9j5UYK1w6u9wCMe+o1jcMGaDOvGSjFW0K06GraARR5P1
Nsv8ShOpKfuDdZwrb6zn98+dAUYJlAweTGlUfn7dBhR5G5nm0REPltxLfZ4ET3K4
/xa6XLo9A7r3xYYGytHAuK0Bn72p3Y2x5Goo9RHfytB1uT4xjkxV7RjwOxbhsdoE
oNhURzIcE0IQcLWdRn/fWY49GB+8Ug5olbj04NpJOLjydlWxC3ms3LYLvL94BV40
FthqKZ5SmGLmNmTLnTxZX2CxUnIpJKmzkB6GtMA2T5/wtYafaV5XCo//xugsis+y
eoBs479u1C3MmX0axbAJfahox6KAj9UZRUOH7FUg3fnKgc0Uyn4PVdQ+6ntesd/6
8izitGZiEoXosrFKNt8wKolwpOT4WFF7eKgAcuUcvH18day8gAshEdVv9y+Z85Zh
p+jmXaUwEQxOzt7Ybr3qYjlGUexiOT9c8I1pEhFb4Qrd0dJgfw/rMOOrGFW8Gk7n
llg9VpU4sxCJc5O32DKBY1gfYflb4Dd93BzIiNnZj3oImkPnqFpjIxlD8mGoowt2
wdfFnGTcL92kUOkdS0sGgWAQLgZKQPjjfhospzb8rN8UdJDoRTYguysq22Fj9S6K
vWExGonVyNS81yN07AloE8q966NwDJZg7huK3jzpRMmOAGpwbiIIwssQguCuCweh
c6DJz4AzBPQn47vlZq/5Fiohlw6//Pr4nrpL4kl41Yf3f9lzLKVC6fVtTMpdITWx
qGcDEENCjmm441vAGGszUvTTZS87QN1gi7CiK+Z5pRw+tYWJqF5kQrzJNE6uV3kS
eF+gNJCkuLCzjaJcE+Mv4iqU7qFXtUpmX6dH0ObtaRYcxT9PLVr6yt0c9NYoPrm9
rHMTu4Nd9pmycypv0XWFCQXy24DjeJPYm1xAVY4efqEDGJ7kmJIn9LRyXN1mIDtq
g1Enri4URU7FhmfWN1EgY7jb0MDhO07V0WjOUR5t86fJGi4t7a0ZpaO2o85zp0y1
WGzgN6JevbdsXw/FHpqOeC5OfYERadiJWxz4vwYeoFzZ8r5xsZ6Gx9TJ5ZZx+Q+P
odDknRhQJ3/ZrQoNxFwTPoPa6rJ8hYwlOZhe5fUvDGWfoIHkvxfLJ9yKht5MHmDU
khRMLhb5G2qTXD/gF0IMBenG0DvmT5I8hnf6Y8vBFXqdemayCQr4L24J6V4x2NZM
Gv3fQFR+KRt/piLKvEpNDLu90+n/0TQ3kbE7UwuVz/al56JUbMXHlC4C7V452Hq2
OGqCD7hzhBUvbGLTO17gWQutifga//J2trYmfFOveJgHJbtSShcVZFpoj+vLKDnd
7vPRJhuSjRbtz2+Q06GRXfpB3ypwYEJexFX8oEaRSAXg+coxXp/7aoq6FXodVWCS
/GGd3x+gxl6J8ABPd/inFtoiHo4ml86f+B/aEPc5hAPEddjgc0IQ/wmAEzTAEnkP
cPaQrcisP9xqvuqYQz8niI12hVWAQKgo05KXmbjTvzvZyc6RErj9gF9SLAxvD1nk
GUEbN/dutiYYmXrifMgvKktuaAfDo5FzqT3dgJ/nv9E+kDYMNLDgaI7SF+ijv7PK
3i8x5m0UaEhYGstztluFtoKJSUyfbdcjHNv8RTs4ai08Ut9yoOzVIJtObWU1osmM
ttZ1YAYukt3LWS08wGTCD1q45C6m1LG1VnE8JWKv3JcYYVefGnZAwM0YL/deRtiy
QqN/nQVU2B8LoAWZMKCLRV1OfaVVV7/yaC1/R3bzecqXxVx3W7NoupXz5yvTm+r3
kujPySgBgY+Cy5aCt5ikoWj2TKtxsqIaHMukdsJJ2eq+zMPmsUHRr/8wOTsgikY8
e9uOmi5pqu9jqZ4KQJFunjnNJOL9zcQwS0grAWhBsrE3kjnIUI3KGviD+CPHhLds
dj7DsxLR0s/jVffPEpuFYxgCU+k4aBTfk4pzdo3TNlo3mOpgHfxmSHih6lrf4aAg
gg60Y5fpo+lj+wBdkmp++klHGAzy/amodq0ow53X4uwoAotwLys2urTZVTbVdSN3
sT2jJ/nPWOgbhWFlKobN2LR1C7aoKYZnTUcqnyoV2lbGi5TjoLx/5UYmeJuh5cLW
jgVtixysGsJE4yB7pFcBNJ1HDMpHuebDLuOVSncrnq8Z6R96+cdDxisqyFHXVGOk
iqCk0iS80Lkt3/2hCkdSdSpDBIzFMOkvOAIku4qUhN0hgogl0k0hiIyiRgff37KU
MRPC2SjL6ip6/jHUaFSORL4dfb6FNxIH/hyUBfuyLaMKn+QgEKm8rqv7olcqGWjZ
XRlE+N24Zl7592xEhvgTgjyghZZU7DpqF+6VqZ9b+Z5ANBAq/G4w7SWW9l/SJJsh
lSNWcCEo2HkIwPvPO3Yp71CiQxbT9ABKpA9rBzY8BkHu/jD1ghDtfjZ1axqW+jg6
+LpfuKfAHZoeALJ7KfcJjSw8p04cVVtR08eyg87itWiE/psrnV3HlxqGrF0LaqwP
i8LFT5aeKkRs3937bJaDjMSIwyALlIXfDBQPmHvW/dqUKcJqnWSNVfZi7rIDhu+H
caE6DGgxQhC1/wF/Hy7i4Y73pd1AgM2nrwHcSUfimVwhUnWNWsvv6ofzA/TnuN6g
kuSEzoOjhd/us2STzinxV2l8LnjxE175p44OKEAf2Nwv4J5gQo88bOUQAGSPrgS/
MczxEC0qrwYjXn7xulb8w5RcOP5eaOPWpVuXslLS3cRagq5Nw/6qZv4cJUsgQK24
WUhFaZM8YgDsVgZKBD+h5IB8TibenJMphG48K2RJgOWdeBMQivsZhIIKxFUrtnGo
wUnH/6ocIkJGPCeIcfh4J06jbtg9Gy7CBj/QK+baNxeYVwjWRumm2yejVubNJupa
LTMZuEQlFnp/UOBA1cBTZsYdvqDttR0Wv+DsRCP/pAoQd3ARNXcldzKVAo1Mvr84
aHGRcNeinnjMEKIaanKjVCIE5uK6dp2g9TCPezuvEe2AJAtE/x5Ju0hsxXsrGpo3
UJ/zVwD0bIR3AJSdQUpM1ycLt8nwNXCizJtXfow4CM/W4btBFzBCm/yNP4032cx/
1A9XkAFjGvEEmmcAtDKsCBUFhp+NwF0mXwaVVQLM2vaUdNeOqEhvuQC/vOAvUPGC
+P2lqDeT9puulWOz8lajb/v+r2NDMHh9myfoftYXk86Z08X9WymprnOvm+0ahleW
kf3NlJNoG6Ibq/dsBmIsQ2X5rMcaUsTXPUmr5FxDQ9ysEpSrmm1lt+A1yCo26brt
bIat3/dOlH+EmW7sEZBH4XaKmTsyNX+oYMlqoNtLlNMi54cnVt7XdgjOljr3IVl+
fhjvoJFaU2FIlBUhry9LpbOFy22k1ygUme2icDFvE/DqIpb9m+kPNUMr+JFsbUeW
PCb+nMkpUN6GoYg0RhI8+M59dkBvseAG31BGXidCLYu+GuQt+anL6E4uXKmuEpd5
kB5rKuA1K/JZKYwliTn+pByc2EdWCkcC/ELUUB4LA7EZd2GNEDPyWd8UvULowgQV
TAzYtSqWTlTAm53UTQThhrT3mgSmzV1FKJyiUQKdKW7MLaJDURotuhxTyKAkc9eR
8cyXpQqIZ53r0mU+GKL0nY6S59M67RsdqegHrEVFwcsplpaK1VaT8ByQ8k7zquE2
XvUy5lmcpHyWD7coCnwP/EXA/JVew8FR38iGAYxNOX5eN3GwSeL80FE6jLtIw7zi
iH8NDFT1HG8uKaozRnB+r/DvIAAt1rYeEdXJlUzh6H3f+AF2PLQwOloRDk7kkDqX
2DZiLjPC492gBf4jl8YOH9jV7WFbMm/NyenUolo5BW4PJ5t78b2Es1xLJi9ijxJP
G1FC+D/RVN4FfR+lTTqUo2oDMiSTNdtkgDh621FC8NRPWkSAIqpP8GkF9NMyJgOK
NPPHPPN80avvZuHCZic5Iqxp0R11iyBd71fFnCKvaKgTSPCmws6kZTffrLqWbbWV
5eyrLRCD1zss1FDu8V90Y+5J3XJrCVZ91LhTC9l3FPQU64p8s9U9vkhxSCKJmheS
oPsv4OOcxzRW0tuNr6y/9beHKF4c3YcYD+LPnSJJzUV7zsdf28Y+cH+tk5ooQl+h
gWtzxyOlPKEKSE/1Kc8eVJJBZMRcP3tO9hUnFCLXoVk5Z2DT1d8LpWaiS8ISOIKp
Z72dbOgmLCyrMzQqFHkdDmOfc/ehKXvuqHUWzGKslX2B93NflkLG0gZBcTSyD2Nl
zGLK8Too3syepgniCIUw16QL23Vzz4BgKFula7HVKYJlnxvjZ0cCzuv3G8kn+1Zt
1v84sXtUxQluJHxUDbK7BqJ6Up491AhhfA5EEXIEYGNWX0kgtmfV+Bf8HGJK0DK5
TgzHCPF3qpkItdjyBPg//yA0Lj15egvqTJ8sync/CcIzrzFOymhDlWKYyhAfPyxY
ZEywVS5BnWSMm9kAdc1pE/nwncUPdxKwwgtDTSeDxmmZWAy15lGBvZChqTqkr+dX
lAA1rynffw+Snvn8Xw+5E/m1NFQ4J8dvgHZlXHOIhWUNGyoYFLxEav0uyAUhSiLf
YirwL9ixfUF3pK9A55efH5xGX6v+b1hGqt4igxY1jDFIkcMYGtARiMI9INlGWVTt
5MqN2KqrIn7DnEmNYa6CJpm/omO+bX0We6ICJcwGUIetgdYtQLkIHycCvCMoQEMf
3rmgpK9K/YBBIVfSyc4Tu+bRIhTp3KDhKvsnyjWNXvgb6MkBiCzSKuNeVi1LuSJm
uHP8lulihYhD/JjdVr+EH7qRUJHRTSh849G0nxxo1V4rPqw4G4YoXzymjI6vLdUU
aF/DoYDCuebIleEObp18JCwS8/IA/g8nhXUFnTmTrhb6dgqYLSxN8jBqqyrpWhI4
2uIZN4GN8hq4y2Pxr70rmv8rGwCQsTPQ9ZrIz1GEkmlbQ9ELM3Bpxur5mUJCzKa7
1UjR+B4ftxkMx+nuCn9q33Wdv/AfbRIuOdG/1SRFj885sJfEYfSL+DIiJTMqbOky
sbWApkiS5U9IPlO4Th8XH9I+CznBbFfp/9Z4/PoAvLHjqZdlaS2okL77PMHdsNrT
rohebXP4LYm7jNpfHiNP8pYfRPiTkyXb3lZqGAmE0kZi8km+VOehcXXMovTqxbAb
ZJ+Hnz4zfNQzcAotA8pPNKxrYlIwCxm+k+FbZ4Q8IVm3QwRH6JXGCpYGesxrseKs
JBkko/ZbBa1TtUmJOZYkBUmIgoStiBL3L94KtIZSymoC8grDCGMTat7BWiOuwrUq
wipoNUqUl4I7I6Adg+ZzdWggZFrv32J9+/SjsmdonqhntLcbOf4b1EDzxuE7fjel
rWDJSlX+vVOM59/AhMmIWxCU+0YDJcUcPFI+IBPP1wsb1OXepo97Pvw1xGZvPxIJ
Qe64R/UvKcMHldP8iPmHQ/K87SbTNkYUSL//ljy4ygH1RKPorgbyGtWzrNzr/au+
P8gHf51TtKifdpTWdvK26ApEjlK4C4wewO1YCJ8QwYQAqNNrw2FBBNhBuLHe9Pa9
2Fhmdi6ZnBemQaEz+uh6NU0vy/rjNmBvcqJ519U467uM6drz15kKM2fl9tVuHmcO
ObONs5VcfQ74UOQZd5F4tisMm5xH3r25VOQ16hOivevXUEwmFP36spihnaKLp1T2
1OCUMf1QKKa9MauWRaoyMSoxjOEKnHRm8G0qWAGQ0gxn1Z9xPg1X9Eqemqhaa/pI
xk1UrZs2Gy9iS8hM/mO2DoYPoKfNhOqSXu1OtlEIsZ3IB+yu2XyybZ/1m4SOdiXx
gy70Ge14WbT9BeyN9iJJ6rediKC/bxVZre7cf57k4b16g97kuK81ozlhxHZZZgC9
ykOt6ARUxHz/XougqL8G6FLO7NDPZD/KVTdDtgE5uWzTBgEzNqNmQ6IpQyVOlAiW
P5JcZ+eIDFdfWd8rP0cDhgKpHC5YXtUUWidQOXDcja55FQxkOV/ZsnEaAXCBgdEk
Q9SVmu9iQiVL9PX+/edj62AvOJhZpDit/Gp73f3iHZh27hEl9/94myBsuQgcnVzO
i3cHN3bQc1LfR1vDJzSLqQJB9WsMCs4EYR++nezTkOSWSJkzxYmPq30/dGrdGG+n
PDLOQLZwEESmk0RFXBblDWhnS8fBu5b0RgO3MhL08d/uhBUSlm3wNI5JO4ZZV6VY
paE6XUww/AOAQCIENOlnyBw47PFj20f9KjfONOKquSRbH66SbUMFnefmHF5GeKPm
VJ7CbtRL5eXH2YVGYbw7i9dnmLV7Gf5Dxpxr+uVbho14NrbF/nuCv5xurkgjBPI6
9r2eXcdx9T0nCTPDJGPMtpkfeBjC30BgdRj04UC1paA5VvHbKq9dz/uVbEAsKVCp
vRC7xKlnvWkBGekCW8UbCRD9M3zqvQtBLXzjg4QS0mYuep199RoHg2Ojf2CUPQBF
CzUvQExz64+OVatFl0h9LjHT6dJoPrCKqWi/mZA10+uhQnJivcpOB01/4Xsc6Hj5
zz4CnG1mXgg+q/S3BB9oOssEyiWDk5Nx4Ks4JLCDCn2w75rIX41gHCsLtRNcib5S
PqB4LQh1mlvbg3WRISlZLuhm/oABdVBc9EIKe5Q6PEuwS//5Pk8VGRQedWZ6rxGu
k39Ad5/00CQJincmfE5/+NbtuQqCsngpUWsoAW6LLKL9u57+8W1q61E8hOCRV3h5
YmzS3mpmRab5/N/Hdd+xd4swNUtLZc71j1nFYipoQ5yfOUNhQFTrlBOSYPdxpvOP
9aHbpQPCgMFbB89bHGCKrFMpJk1RQUnYNufp0NYlpqC9UfVCo03SWTM2QlOMSAtS
h4AWOZHV7ynnCO1kPa5HUqJJn2pl+wsRrLDgz7WXI+NpcI1XwkOMCMrRvCWhNKjO
0kAHSSy0tYNW6/E/piOtfOe7IX6oNOcEWsZ/pX4kz6wPkaI8hCVceNlr62tB2POr
H3SHGT4+whYM433BPmjYLfS0wTEc4PHXWHHHziOOuuw342bNJfmKipstTXJMq2n7
VIYrBhT5HjNlStk0MklOtIm2mQxPyw8w2mI3A5YGRLsV0A6U3vDsaJs9yEMW9EUR
p4YXkFSt6heRLWCrx23c2paNds5hvOtx0pwiJonU0JpVDAEZoXp6ssMfLBiBKIS2
e3Pd67M4Dc0vGHNazbXf1g/ujv0SGzplOAJTsP86Vqk9s/6/gLRIu0A9XTmIf96S
nwlQ8UHyeA7heO3NdU5izWwRCWl7Y2m3zkCb0cQ9md6z4dEU0KLLQLjEy9Tnj7PY
hZarmQKoQt0CryB/i3q9PTESZPNHSwLJGZBS2BbW5bP7qryddcpzgfENwqFUr+gg
qmohSkoMmVRoySEnhC0Ae7aweg0KO2K6rSkeUrtplQLgYp+LG5CthGh5eRbH/lKs
DTSB4wPv7FwLiXTrYij1GtLd+vqxnnBIoZtHCBZrwiFRHnKJD4mk+3xAYlQ2wuGw
Qnx4OM7OWtmYVJWzdHTXGrX5uUuqXjXxB5CNzUvYZFUL/eb2AeW01YkjrjHGEi8v
fE4W+EcHY1cKsQFOZb42rDV9beZe2nFmjhddMjJcmloxraJAMOAeLFP6G93FMBhz
6nb2MbreR+KOMaTe719Jr7lYF4fOXAjU4WF/nkN3J3b7nxQqvjciCORx0UMvLqkw
E1d4wE1wcX5aVzf7BnYpQIPLGqI5iYgHJfGiGYt5k1mlhXjbNviQ1LDVojoCQxUW
sGH3+yJ+cAI6z1IsDZdG/kVf/XvnlbJPRtmYHjOTRI8p/BeieIiRrA9+H1Hazzaq
9bxijXQhoYuB3oR9U9E/exEAEZQs/PAG4+Lvgf8cP3WVxiKq4AS/Lyrp00Heb4Zw
J1VOER69cGbZHst6vwaIO9qogyoiPWqoV23Nn/lnZdXxk1FJWRpxg9DGeRiUcksP
DcVlN/Teje6RTpZ3PDScLhpoBERfuIVAfr+PKel0CmfwlgVmr9cxXRKunOc0Sz+s
1bN5ekXrrJwjUMLJcrPipxfsUFQt38JSqVhBNiVTm4g5KUYFRrSWt6uw4ZlvK6KI
LTe4+X9ZYjAb+rqCTdDLC4DkK2N2V2CDWQ+a4aKGK1xCQABaPt+ppC0T4HskHGhV
CQ5uTtpuoU28YkHGzRz5Rej1EuT/MXl+7y2iu/HsTJmK4ibGQphLyAt0s6KFc3K2
F0EsCe2fARt1IVaG9qhBreo1fevSImn2pPU/QrBVp+XsQtn58TlQEuUgigIA8zoT
7ZYYnmgiYl8RETbk5YqpGoGZ2dqQmMLj981U8I5Ls1cj7x5x3qLxc0d2ONEnbU8f
zS7ULh2WaRMTDFDvQ8vbrtUCjwutxmNkIUZJWNpGNJQj4W0GazqvuB/NAV5FBvuq
wd4YSmI7e2QNuOBXZ3DeGLdWzw74zj7LzygjSVm2+gCajZc2VkqwdP3vzwnHPYXO
cZmLJcOZCvoGP8rskO3c/G3HNtvqh2zk8v5Wknyr+hBNwASDeeMcBm6QD0M22OJk
l77uC/tzsER8/3DNhKlOFgtSaPJKRmm4B/WujeFM2VE6I53pXOVbOLB5KaWNCdJn
1epkCoY/onruHvWlitGUMlwgobWTgZ/acPDGdOXq9S0UqKI6acl1sUUGoka625Rj
hmuJeyT4ItFs8xnQjD8xGHlqB9MaolIsT9OXS6nUoay/8Z1tGX2eEC5/ZKalTqRg
Ax7dmRQ9ijJnVqeldg+ecXPemVOOUp08Y2p9tKYIBwWbDCKCZu7ppthnIjIiBuc9
Q2r75s2IAgCdPrG9T6i6ITR3rjntrNWbVsd7jIxERbEB5b/Fubroa3Y2rWrPQYgs
Jm/awJG1GsODR5/cPwrm+f0ao2+UG0snPKByb1nMqj9Bgnufl7Rg6G4EluuaxJlv
RcbE9RFZoomjveU/5BRp0VPRPgJVZhij+UP3goEMNhdu84j4HOqesNdndXyLHqpw
LXIZl31HYjXUsdP/woXd8pH5cFOBDTGyOlRWnvYTh0WMtNeUvBnvXJYgNVGSaGW4
M+9ZDFBsaa51uqx9vBApAIjunIKI2Y8VcVOzObo9kbFSgt47E5LuczJ3pPPhQ0RE
r7f+lvvT/IJXR1HPbqZy2KBDHiXJcGdzobHVPNIW3LrkCf589dghsNV2PpyMr7TN
GHruCoihgSCl0i39fn40N5l/1ss73YYjWB9J4CZDrJh33uRynYjcU4REQ1RzNeF4
GYg6eSt6fxcPymHKEZJy77JYfv506WZc5zV3S/V0naEvH5Wwyl7H0UM7Vo99Tgf4
8XovkTe0H7lxLZlFhFVeF5bEvPxFGx+fbpSEVDNgMbrqyg+9O1NUUn/l8U+JR+0a
Cbr57KBNZLvxlPfY8JyNVoVryRRboODcaearbDGJdP4N6j0ZtRRdrAUdVLVFBytX
453Tpp53ICGhY/PJhlyLF23UGX6Cw593Imhttg24dMMr2DS9Bl31psrl1I47tClw
5/DSNw8ahVwo/sxJerbl2ZlMtILjVH3Dt+PfZsJMvxIhK4reZcabmqxt41yIU6Pb
CLjAJKm/1hVHZFlpjvpKBLr+W9H5vVZc/tUPRAP7DS+wsiHHM4/L+TBKp6f0e75y
U4vl5LD+bGdJhPX2kO+YNMC/LV7Bw3KEt/3DRY+Zhp/vRRKgnQ91vRciUjoiXwVi
JdA/l7vzoeirSU3lu9HmNggFIsDAatz391/qkqYhhapYmOybq9tVykoelt6BryB1
SsLi5Ojov2V+y+JMFVcbz2rYMZP3D/5lz0V72OniGx/OtGVa+mrs3D4IBr41fPFV
v9+SCsQ0xLuBl8XXD6OZoHyQLjXrL8PpynrQAZToxzPr/Hvt7YaZ6A3jS4nMxb+J
x2xqjXrLFIF1ubYpG3Gew5nMRy9taku0kbV6PDs0PrjhEWhGtMGp9eAU1e5jS03W
5vrKNjBt7NVPyi9MWjSNNCfcFrKT/t7WiEoGuXN43efT3aweeLdwTosQYVoMV2sy
3+FVVYNLVkN4RRXMX1oJU2O1RfA2Jpa6Pl28CXhq246DrrUdQbDVfmysL3bQsLmR
TXaz+1DZ21b4yei3VnSYFf550c9Tec337bSLQ36KQH0rtB3SZrEz3pfYKUYsq5vp
EnmaSO9ozrzJFq/NzxL6E5er2CYZTUpHG0b/A+L3D0TZbjqpaERqpXEFprbJnwmw
mlA8Y0oSRVMwg2twsiz3NVALIdy0U+HAqL2Bz4gZrvmbBuGUpy7QWO46EgDVuI2F
o4hFzTUXZ2dN5wXxMP4OVWY9Zsl7wcBEq5cr4hgP9OgJwiqhdrp3r5Cs1mQs/oXD
8ZlhmXFfcTT9wUbsjvkdKWVlshDFrqxrKCjCxEdXKzaNQ/m6HEwQuAWr/ZjIYe3n
m48Mcv12RlJhXwzGQgqKkUe/qvuYviIaG+Y8GEWkI23CyCyjAZFW4+cRAOYvTyFK
RvjYthO4rabBNkkvz893/WTTY5B9c/ubeoRNldICZwx+k63qOx7YQgHjwTffYf5U
YzTi5MPiSUtJDohulxgnagjO4HxgZ2Je8RGL9ggoMi/le8emfj+wsiRYcj5nDnGC
+HaQHqB6bhTalZq552l3DMk6aTl/HLyw2+tlCzGVFk8yyU6XIFfpM0cJr548WHR3
wxVjI/MXJI5wNBanYhrx10YzktnlKx3AcPEaK5nWxlbD4kgoeAzKCITtS8QbfLUp
IdhvP6mpd7RODoXbkDTkWwslBBreoSCsYv2HIm48QaE4BgJO9EUBgBT9/ga1SCZU
YKWXtZzh95hLbDYLyuvkvzU0zQhnkHfnZPwDPbhzdWvuP7b/9IUPsEXqlSv3Ndex
ebbJp4CvbWiRi55S0ohVErab9+bvlomhj8vKoJNi4VIJJBOxtPsEyf3cXj+n9XV0
mjj+DWCj9L+/3ZKQGP3b5krnIl8+m0ZG65VCfNhmx+z7AmWDcjO06fx8pQDrWNsX
c2gKySr/Qro9ZFPD8pYXlgRE7bufB5eSs3B8oUHcJhf3Cpbyvq4wFgH0lw7UlGEc
Tmy9rWTUKV+g5IBfo0KKlTTcSmxC6mfv+W4w9PckguwU9XBwtZUTwHOqsXR+H6aW
zXXUMWtCudLJ42ycxAYFhzGH31X8ygk4mSyaJaGQ6BZLBSQ3PMOpCQAhk0BmQQXq
rN7Alw/lysMCp5EfcpUTTclXV0g7Inm3pOm7Zc2sNmrmH+JF/XxUejLC6/eVH6bc
5cKsLVgKNwVI/Xfrjl18ROmNSUJ3GJJKSi5oB2OUZBZ3tFItGOgAFL2dCnKoxd3r
rLSN0ROuJUZB85RF0pbyncm8AMkYldQIW1Sc5FrlJe6j9KHNLJpnLV+vjGsopjwe
d1KwEl4fHlBvbZlrK/jNdkmDwHcL5aRvS+QjPAgu2NyUBi1/8jkwnnIwyX3ninDY
2FRGT0l1X+3YtMdEnr49oEY/1PnklnWPj1pOsTtQ3X4gvnDXIXXNYbzPo7hx/Fj6
iP4Z7f4SPjWtG4qxIt+7wTHVew4Nld12DcMzJ5nc3xmNm51kLIUBRu/4akAxCwhJ
tY/1KaXXqZlUVSWodWtQrIQXMA1ZqMDUnbFebHJV9YHIehbySRJsa4GKi8w2EaY0
fG6rGHIk/k23AwvlcQznyxqnUvDG4nyhqdzVmS0trgCaeEmE/2opa6q+Mq1xgYHg
Z06Ycv+oGOfcDr2Y78BCje7SF8BUPBJyGxQSkGrV7TKUXFEaryIaeJgw+Mtu5flb
hVJoag1loiNccSZ+aiZ2H4Ra3I6MHlitKC+1SPvOQUpel3xrGho5tDDu5V3G67Oq
OJGWN1a6nxghyazO6Eq6N1wjTHg9CDusunxEoJUN9Fni7e9nJXbENF7Uj3X9KYTm
rhdNJjfaEhyCglvOtjDA0SBbroOgQRzPoktPWalW3izMzXMQhvPfZKjfepqJUJNx
H1HF4iHs6HH30QPd+YfBe8DyYxpFqbqrmjej++eQt6YOMr0kFXf2alHTyZWMt1oT
LGg5QhIYeFzdWRdPVfYOmOUFO9qGQLWlFyskr04nluApQaFZ0Z5jgna0G9n6WvCZ
wsuu0mlmSFxEUppXHqBDmBwuTHr0VCFNQQZEzl8CG9/kN7D4MDheu80FKoNsXBAZ
zwqYDstFs85vXezM/TcdORAkPCBxgwJKJcuH+Ju/WV1C6HiYnMWi1aeMrL0dookX
SnkThRJLj7R1bpPhYA6hyJqHCzqrGjCBnXcM3phn6aYh1GtpTdygE4AiYMzmUZlK
a99rPAueog7TSQ8W6kwdeWXD2u7YyzsG1SIdM9x4j/ll1dj50vRSyGeOGl3r9095
K8Nd5bx1tX+VK6yl+oyksXHpH5iffwFMHONMNF4D2xz2tVKrritqPh/DODbZKoI3
+avRTxI2vgl0moBI2+SUEIUiPoJqxnjSvZ1gr6KlJW0htexWp8PVSNl556fk3uXV
OPtczuaDdXZvuktZhkhseZqUJc5J1SR1nloK8ve0lajPhRZVxN0CLCdwqUSsSbW4
OP2DqzFO2yTWuxmPVXvgcYxJ34GdIstubKKff15FKdOZKhYURuLZI27RHmLvziJf
ikkdDwiuZXzys/SeHBHJb7zpkIWc04Fy721LLLOGg/HKy4aZlap6ieLY7hTHhtt1
DhzgeoGwLZw8Idgq1rLyjTQQl4TNmdIL4BI79f3Gf6vBq4S7UWxTBYTbgGFwozJK
VzHc+SPOBMLVHGU4P8QLb+AQ2oav1tR6mJukMUaG5VYCsbF8jCbfTVwGzmMJ7t1g
O58w/VNWxy5bhvbVBke86jGNoSGFprocsBP9Kdu02b++x8DCespyJP1uB0o5esFw
F3s0qCwBozN47KtcJtQttJE0B0FRMff4jnhF+iORJNDiCxqgWsJWeEyn9/gE7brk
DlkmYFWk8GrMU+Xfm4DLvtsYRTBJhVsLjN8XMU7/FTGw58Lp83RdpebaTpiewwiq
VIbX0IfKsqp6Md8qp7vUOfOVPgJd/dAL7BBJc1s1qWvdQR/UjzZXyp657e0Y9jAj
86OL/jqJ74eJpE4FfbGzVI+rV9nbT0y/eHptPBCj62iGYGeGjBpmk5mLcwAbnbZ3
aW8f6mgArYTW9ph1oYDX5Lc7HN6+JX1PdxX5kiC7w7WSxdlhna5uGgl6BH3N63J0
P4MjqOiObgxJJ9uv7eraIFo/4K74B54cGkPqwjzWfv3fxAV3+K1a5jTqOXQ1Z58E
G5aWjrDTFiSdm1xibeoWneUqU25OrqETyneMhTylYqAIws0wknW6mM5OaWAvc37E
BCbevmcFm8F7fQYw6uRUCVA7e1AcmhdzLy3XkuxhGgP6cQMtla9x1JHCcdJxs1OF
bLqXeci4GuRp0QXUF33uv660ud4J/8xOA0A7aCdI18yF0wgf4smFFf81Wmvzv/lh
3knnolzwP5XV3uFYGfuGwqcKKacU9mj6razuQTr7nK1dnqJihlh5ZmFs+VCvIL/Z
nTvv47WPcylh1zsHdg3rvSegRhZ78uOT40T42+mqO46PcJsZ2wxsV896TgE6YhKp
alsXaiabajxmMnmR8x08IM3Ns1EB5sTSRI/9oEHml0OaJPZDjemV1GRe+304/f6m
hQgmRw/+DeEo1Tism1SU7pkoRQCcoYv+GRKMOjzN92A3BrdPzFCXcMyLA97Mo26r
N6iO38FVKmDeqjuxv6cjYo8FDJG/oKutfl9kkJq9xRISQ1cVfONbGzItIP2inYRY
4aveFREeiKWTyvLkBtQ7s+DUsKRruLho3iubVhffREjoBchmsP7lAUPZDrEcry6/
DDX8jYSjkKwq7plfi3zHr+qLEjXKsQWJhjVIM7UG7vH+p5wQ6KMk04OgRDZk+WoM
JbbOHzHyaiZGA8dS1Whp9PDlNuxFJSqIoyXMVl4x2Y04uc3lmiFUJUtF4ouaXDN0
5dM3idxM1cpSZeZW0pc38uKCnUEYtv20l0NDN5elbgGO33zE6d2F67lOa6ZXqA7K
1ckjifPxD9+SC+9YSb2s3VXY1+Dr4VSwLInLVKOuWyY5bJwX9yzatbkPVSd3lKLW
MijrWHixNp0UE9J43HWUe4Zk7iMCSyGQCyUrc2apJ1yUt7qYnzCUbm27aetWv1dl
DT1lYGJlwDfJUZiV0rjGTGyKpBwNGXUf+NWrjX0uB3fKCxXxXedst+zD1qMjNCIg
tWgA3rxXR2pOzpBqkHMULYZr2MTAEkiOJ3n1+jFx4KbIrDd/GEWDQjIlYfNbqqHX
CcSrNoOXHm6xXDkK8eDKUDYHqRr6CS305G0r4+VTZH3S0OTKOcYg+7J7Z8f03Vz/
UrYSg7ViYRu6kjiJ564zlcLxTJ9zpAxCvXu41AiY8Covxk5zyta9WBu8T/y/Nwxl
qwznJAI81+5m6Q6j1vTAcJ9WnVtHsiJwpw1/AmXMfobhAsBSg72SaSxsPVHPwKHd
Jqx1c9b3/QCo9Jit/Awg7wY2NVSHokR6yW59DuwLxfNjZxAQ1PMvZ/1aS73taw8E
+EBg1u8/5ElTYpyzFMW0vfcP///5fIP9Jmr2K/haJqJHsrog3kMogkIhK+aRV2j7
ffM0p8pZxi4tzueP0Shy/n2Nt/WKMKTTnNJEi9/q4EHjsa41v1xX6PiH+eXpRL3j
rDNwlSBdUqiZwywsTtZ1R91IYHOoxBzeGVXOP2fBuiCTC5D4wTyCR3AKghryeGhJ
b+wnm5DKPJgoog33YIdScj1E+yY1hrD0gryYIzriSl8QmZcR+M1A6sDxeG40w1yQ
mNwVDWP0Q1GHG8RXqDAvt8598Lde7IKTCpOapsN8U77vdbmrNQDCVR9q66f4fA/w
QfqZU5gpO0q3EVYtSOqy+sYenM0MMnML/9dmZAwhsks/lcDTgFpOGOURLgqrZCbg
niD/ZKsl7YLErmYL98d6TF9V+iJuQEX33+rpJjwuytyBJ9OWdEKta9VRgCzKjDPO
rNJ0y/ukwsFMQ9Dp2e/7JJHNjtiPG5qPlUdzndSPpQu54XoJq42mmNxJplQ4XKO8
jGTUL/grwVMpxI/gRxZXgyRDIBQdW2qjSWkVZ0WVpCBulYGLMNHqFzlwhVJUKsd5
3wPhwbIre/sPTgRsMHiKPvrz66OTP9fVlV67UIHDxxdSqmxTbTWqY9uEe4cz2wbD
gCYHkiPOtEbX6Ls9mQnsZYvr8mtgl3wsHUSm9WJfKvJDr2/joFX6xYMDFwH25Ezz
BkiaocgTmuLtl2k/YsAbJLKTNMyAjzBKP1M5AoKwfAhmvhWQy7VixgbWFdA05yHz
AVKKP0GwOIo1VP6b+tVRXlMuN74PU2ZKJu1XSdoiCLMnnoS285paeNr219XtIGcY
oarhUo35iMySiAWk6jXxQU768P7lTTO9wNX3J0tT+HDAHPpGB/R06bYaM6j672/F
mkttN4MwdoTiMYNYZRbF1IVo9R1hNbb7EZyAdyEZ6HWPGpfAvkMmzrMVpL8NKYtx
ElXBhmi6iXUf5+6mFeReyQf/PX7tv3WSdIPq1pA4hRBTVccoEpiUXMKLHBoRR4r3
rtS0vCQ7m0j668Gc0HoMaaF8z76+UFK4z179EB9FvRYboyka+aA+rGnrVcy+nEH0
bbPLhiSSLm5X+DlQNv14XMVCrREku/cQfyIaX5+c2RKq7PtfIH6zjWmxALbcsokc
HFJCPScWcc3iIBtTKmTopCST208QdyUQZRTgcO+LqGU+Wnig7pNmzUWG542xmDJk
U0OHhIO6l1lj6YqLsuVdSS7LUPunbg7VhjmhGNjQQQ50DR7sbs5AdODg+Sdoe2dR
fDoaf1XOUHXpnq2kaDNqAwWRezK2xnvB7moKS4zmVIl6Um3YnqmFeiODw0Q0WSml
JF2hphpB5bzPrlTqTWZGR31Fk+8dLekOf/LgCrCo1iMSXvr6siO81bPMIvwjB7Yt
GGG2DQvsOuHa6uACzTMgbaRLOoTTF85SOfIrLlnilscWKdy8/HUMwD+oeF9obwhd
69acTnXKJ/lwfAbplljxxaL6IoK05uY2YLHeDd3Qcxwqf2ukHdRuD1axEMpEfZ1c
HRmecIRoIdOjSQg5dCg3NgdEfZppEa5Wkr30EKnwJOr9kt5DswImEq6ELdZDVwR/
fPmk6R9vxCCr28N1EOK5IyhbzR6pvY9c4ZO/NN+9/fKYjekP9JuBJpMbN9o9VxUl
vLvzXCckdxG4SFE5u6Aju2kdWwDR6OBg5vbFtJnI5LgeeAskQPyf3eEfkMI5VIRm
FS3QiVa9guXvsmI5Vcx0GLuHCxqvc6d1pS/SoKneARJBFPMcui/4eKJjJ2Vh9+Ip
+DNAQiebJJHd8boyCJaolgqQBtKgxbaCtsMGtGEpTNKWPoMk9rRydtU/DRPVTYTc
Swr8O/Ns4QYLWp4qL+6uFJUiKZx8klbV1UMu75Q9FuwHGlPq6x8zsUFToI4dJgaO
SCFPwo368Kpk2gmu04eqiyXi44Vc+yjD3NaeGJJie5BJP0aCdni2OOW12aeu5tdJ
NMAC/pQsSlEN0OGYRQ0wLEYXiJh8MqD9K8W5Y3wDanx8L3g1L20asrINEtIAdlQo
DWr3iflMRUIK9v+bif19op79vFZI7iL3JSvOlgXd9cG6nTxE+K2WZCm18Iazxm89
oqZIOjfTiP5klwsf/KcV3XCvM7V846jSDEll6GeJm4hg+8jnhfId9zLyNy53xC0L
2e3Lbg1aT8XfYtCxs8R4fdQf7qr7Det3k1Re2MPp/sxD5SlyJ0hC8ySmLkB5TJlE
x/MKQkJBYFb3HA/DIdku3YdOBST0yIuxltF/fXLYLPlV0jptGd9cu/fIEU1mEpdk
iwfl5fMbIiUs/tCFVXk5IfAMwmD8PU8FIXOT8FBXd02gX21TnMeuRba60V/z8u2L
4imX+U5b9PNbrlM4H4sfkAhw5QmMjFHbLyd5qy7c6yu2SY4+t6/BdtE4SF83QkyA
9pBCq/lq1z4yD95HPgo7xfy9+lp4at0m0iIZCT39aHwNM49HkDHPgjSrYWg/T+Sq
f20+8sVxjbztlxnVXjaW+/aaM1MH/zHOtKYI1w5smyDft644ZDuYrief0tHZCiQh
eIhOEGqHhpxp2px/V+JsN7GsvAAtCpiNt54fjoFPSduDImLTuGU+5hdY+nYBoVzj
WIQBdnUYxOBWL7c8QAH8hUamvXtEqZ2eedpL8zbtwCZELMdTIfqiZJJZxCvudBEk
y6nI/Bt7PpVEMvpPuO6sCmECyd2v/aOwiqIuZ/Ykx5cXOk3hwe7xtuAKJFpoPzno
xdXjhZB0S+/Fi82tbWXeRFuns5FDgboQynDEyUJvG7yHCeHIa1S3qXqVYeumBSEb
DaJuDYUJsA2OLamalZxVvRcBTziLZrTxIN6ej8LK8OwBaEg44/cZFv+DlJpdpbbS
egbqju0FSOSHjIzzlCbIW8Fgacw4PcpxyOxBjLcIEZkKo4KsJFEmNlKmsHtLFhF/
fn3mXzngTG/7J2Z8u7z/S9ImlKt46ml5UPI/vgemIbHrFycIHKoyKvDmy7Wp0K7K
YsBFrFJWJXioNN+czk3f4iayfAXTwfSUPe56I8MFAbIWgNcDfswp5KMBhPCmHs6A
sDsavDAOpZJZM4Dfhy2aCKNIp/0YHHyJ+MX88kPRn9LUq/WYDaLDt2E+pR4+Tzbc
PTg6gaPqC5DrGHjjaCsMKW4qvZUtE9G4a2NLAGBhnmOjD4b4KLfaj6PPFwugbME7
lzLvIS/JXNIu+A8QYI8dacg1KP89w5rDG3KqFGvlVTxx4PhBOJVzySHRzgtesEd9
c+pjK8ZhnxGqiqF/q2bZjYSU3MMdkfxx4+sTjEmeUIfEufQD2sbx7+4pJLJrHud7
AjCgcOFMaT4ddijTCbKnBc4TLMZ1cYAOFFMydhWZLBhygnskuLmCli4pyK0d2uL4
nhRkU5f5iIa31EIaBEhJ3pR2Z6EUagvBJ4RQG++AYB3mWV0ajjyp/u6XoTVNMasR
Ovk39D358P4ugjCz4i4nyjmpp8yxyP4Tnfwvys2WXvAAKWor/K9BKz7jU9JHDXjG
gAMuVgRFp/0cGZsLNHxGHIgx3fHlw6JD1SHQ9QfybHju869+MYpCL9QAJekHqgOU
659/m3/PtiSznb6fX9EAXQZdAJVy6lUeHofjS3j0mMHVUUv/eCpPTa1/4C4l6qbG
oY+MBmQ8diZT9ZjSphluWEmh5gexlKHc0EUOvbcwUQpumTyptZc5mtq3ll7AOe1Y
tQqbq2+ejSeAx1QN5HhWbPFsgVrLJaC3EbgjJGfJZyv1p0t+8NhoJMM/CNHgV87i
95o1M3YQBzoS7uYEvZau7KlMHbzSnQsQNq4LweujqOvP1nUqHyIdBTSUrIWVFKhT
NvataQi6+ROm95Y/X4Bke7AQTSw3hJRD0lYJeoKhflsEMJCLUH0zaYUIz1jRngRB
n4uAQ2545OQneBXEI5/Prid9L9gxOP28CzcNnjS6XsJospHOLfh1bIb0MJOafUY/
gjhWKAp1mx0HvMoVr9us5CGh7XSe+L4XbqYY4feNCNx/vvcHkjE49p5VH4ac+gi/
ovk5dgXgWS8FkKhastEKzK8F1Su/MjUCaQjP5HXSZlO5IakjcQ86m3rF5THzUNYv
J/meZgqU54/mHCevOC1fcO/5m8xZZ4Cz+nviYYFkixGtyO8ox3NrtUfkMYXkg2ht
sVF55ZLNneEE3DBSu9IuEpp3UpTXdq0vmVPEqtqEp/7JlgTHvuh6IJzkPvjd/wxB
tpsLj/MSPyy3/wLF3cKBj2irJ3GoJaPGUJ3wU9bvwSyyqo/6h1zhbJQ1TQBATgja
bZUt8MAhCsKrS1hF1V9de9rAqrXO7WhzMQNLdWfVCZQFeqNdj58lx+YGUkYhX99z
bfXGVxFLd729x1y4QdNGF7CljDQ+vOMgcqlIp2PAa/i1CAeRCX4hQeOqoxoDNH/M
w6Bu19iesOJ7ECf/I5Etj2n1sMnbCGjxKu97B2pbtetzsCdmUoenFIFecRe8ENBC
YVzhwHRickIUP8F+QD1B4gLH3ayiyMOLtjVsHFK6PfOqH6LnXTeu7aCiSJmCW8fC
oPoNSESBxawzxKVmxL7OKObFXdzo8BcRohvKN4cfeRNJplQZCp5iGL1JmeCypFHg
vg9kElZ2yQtJzXuksPEGH+oImtrJFYRBGzEcMl3Tvz5oQBbB2brgM4bPKVzjdvoU
LwkopjdDAqu98MS8SCyXt7Ze7C2Ju6Q1UP0DNWuq0nPasv/0+jRL8sIObEWvxqrJ
UoU5B82P4dFiD9T7gSoUUp8IPaOeAI75uH05TJyx3ekEzMuWXEr9Z1iAwZ4A/KMT
v3eie/nhQBty9a8RaLoRjryqWE7scmDKs7rTD7TUMa7lIDeiKHNUcpBcF1H4R8Mt
eWaZA266ZW78dfddNZ1scuZBghcvuuKb6ZJIgqLe8gf5MG9oEnV1kc3Au9lUv7dc
Wfy5SeDb85+j9urX3nnroF0H/GtFx7ZzOsJIuwUKTcJHnlrjVfJcrN/YtK5l0vqg
ey5UqCewDaZ4TQ2kYB4l5ePYJyljx9Wcekb4d4bNUfht8tmvX957lS/cKaGX7e9/
X2kbtaQPQR5eY2ZvTCPWgPwWqqwjy4g6O89oYtj+FucTthTyvQtpXRReYoxSeEiY
bLHaObuqd9A6OHYU/xiwfS3v1SsAyNyLopnKzy1MUFxsKhxogD+urv3iKS3ylzI0
MpxGNeG9aPElN3/rDCTgwgznqBjAhMXmm8HEYC6smpte+GnO1v07AgLFwyXVw3tk
s5cPOhPhEKWK/6oeLQERPxcepDnjT1OLGRe6XEUuui/JTX4LQW37tdHtOMmxs3mB
WOKeQdalHnkTccWA53lb9jtpuMG26u0r8h5K2x2dHRKPjiMj5bqVCFpcqpd7LW3+
IqXXKUwYDJ+AwYS04ZDIVEfYPCZrey1/DMIQUcW3BgGnRp62d1U49+roOqNHtkUp
oRNtD9NZ5803EAMtksu3+7IRMRhtLSpFQraoc+GCr49sXA4L9sbmUrNIzo48hrwC
E4Sf8ZNue5pB5fDkSy9QdjR2UjxA9fcklqdNWrV/l4zwJZ7ox4lK2x8zd4Xfr0ec
unI1WvJuVkF2FYAV96fmvblkOGCTO1y0+BtRLltKf/VN6/iO7KVt9QmMjGCiIxVn
2OYApMG9vLWztsRyf3gLOfJLQyZM8oKPK9h/307uARI7hgxXiD+FJEO+TL0kJAsV
r3oHNmWUL9ZfnvPpVqYEcxWdHzGIpZEBu0qbCD0o/0IzcLlW98+HK2Ik6waS+EZs
IfplzFP90wX+uqWr3BM555BLP5bahw3/5kULzwAA1NMKKz2MHZMvhSedhkekHrMp
lL/Jy/LXFFztZ3d3d0sOvpTSd1/9pVYy5OD0f6RyN/VCqtYHQwVtno2gMBCUca22
IlBrg1XvQ0Ujg0oyITI3p35ecl+gPwMEekisxSL9oUR0BDLul+ccUmBiFHBPO/m2
4lymHChDmJDM5YTVY6+Nh3yfK815cJclywcBEV+o0Q64tmnX1FVutitvmjLt6KAi
GT4G+JWAEzvnSYH/NVz3SqF8pYHPCDUgp5Ka89w58OIOYMzxmzMkNHC+purIeq3v
tocgFJZvEf22iTMTXhzwrSK++FOphkpUKLqiWMlXGvR35/L9aeBZnSrtxUOXL12C
U0cJmO4ElKSkw+ghP6CUhVwnZMyvKLan2g+pzBiuBG/qLBvC1fF+xXCb30RXUVwc
o8Am9KuuhAWZPVNLP/FLWxoKvYwNOQbteGAhSywrqKODxRuKOfdPPb9EiOTboWED
4MmCzce1rTx+psrEwNAyc5DYaREpWJGgWWhS57u0vweacDcS+q5BLQOcGqUzr7NF
57QNHj2ijZ9XztZ4cTCuGS9wjAqVnDtIdZKEzdlPZvrp4Efe02xEL1ov2FfhNG5L
8IlTVKi+n5cDDK3sqwToC5Bhs3KcvRvj7IEolahx2nmn7qpcU1vj8zJvXRKzL9I0
2EzbctVdyiNdcCo+p+5joKU5FceEWpj6m9YeTiq5i0kMzMplg7x48b+QQxuaSZgk
0qudC0pt+G/7IOhUfXhkVyG73nNcfFPfp95yX5vWWNMlylnxulq3kzFriY2LMvBM
+OFHOeiCqP1tNveEJu7kKYPPZAPDXSLxgyw/zJQ1VYMydc8o5bVzbF0nEi0eE2EW
ETzxHZmlvJhPGivg3GLyIkXkJ2AylNFCg3wtKDuNL6WymX7R+eoGMOl6/WaxbiUM
6tURde7KWjTtWAPnOGDW4Imkzy/DwfKUWmhb1v3I2QVPIFXt+JdAtnMxTcDfNLt8
EmRHX33y7g8TXFUwqe4aOHe5oQOnAULiIWDfP7QN3PIHQZ9zSxDm0Pl+g92mJNAb
Pw1dVzo9r8k59A6vPknU33PdgQmhTb9eZkPpA+32CEBR5TxAbE+tnRGQ3W5XeUN5
8eQ4iyrUopD9jikhY5A+iBpFcPahbDSDl9n05NsitDzrvgeaSEmwnosY0H7UORKk
C4UF6oX+YLew2O5afhJvPt7h5dyujPKHYdtiVtvgdukbQRBU88SqF6Rwvv+5V7vM
tvjRku2dlZ78aznvcgkWGnJRqp+LjJ70ec9orGF3m+BgIlx/E/1L72wfzLFOwB0p
bhoNux2UptOy+x6V6a30QfuvzDxrOWcIp40SxqfdMKYKg9weXX3mMKdRIyyvUzNq
+/+NnfobWLchHKyGUmz4WrlqVgqSwNh0FIvmEts8vVlw0kTSbsneCtncnqIkC7uf
1kfnDbJbMYEBw67zdE9W4+Y19nPHLNz5ZuT6fc/ro/2yWaEReJZs2tdxviMGDxcQ
0ZfXam2HDacfXdL7M9UYTQylc7i8Bt2OUYGWjtp2U2dAB5lg6sm6ek656jf3RIcV
f69n9/kNP4of67sA0LFdL/gtNSwHW+ZR7NaePalmOYxdn6Zw+hljt2bYb8ZCkTHN
sYtZJkP8bvC8qNQkmO5tar9ox1wAeyHr9EvdfCVotW6mnfcy0Pnzr0u4i0RWM7xJ
Q34dxXNTcsjpaT1kjIiOlWDXBFLuUa5PWi8rkfAUByCYJNJ4FdXClC68j3WbtfGB
SwuQ0iIO8lYFLktUnvC2yMxn++IBJCfsQy2Z3n/5+VhOhorX27D/DIkS+vo20iO+
7nTd0hmnqlY3gDZ/U6vW6eoKbNpBcLQvut2XX18zAzLKPLMzd8CYfG/KFwv5lCJW
DPOvsQQLi/rtkzLav6MNsDfqWSZ1rK5hJFopWnrvl0MUtJNu1I6lxVlgxSeBlfX+
FhmC5AKza3rMnjrrBa7Ibq9qLzck/n4JcqyrwAlSSkzxciyiv8CBzSHGm+ovX2pN
kTQHyBbILPLSrnNIGTMCLqVbZhP95RQE3Qd3IYgFRcYAxI0aKLn0mHGS82rfe78H
J8Z12M7nIVUF7BvHvlLtmfsvogyQBeD3uUb3GPPaoZihfPuSXHIywPgA0jmfZYqR
HLABAI/Yj40YI9MRj1fi4iQ/NEcTiBKXw8rKY8HhNiKajW8KswJi1LtUHfeHRJvW
6B7m0I49l4jINjENA69DWXR2zGm4Goik2NOGDnofdLg7fXzXBzKV4Xta84XGwWnE
DwlTpLnWkiRlQDgOiy1cKewpvqJTwmjZzX8z85gkNzUIe2KUY0Vu+rStdJizqwAi
3GoYDitJsikobmdjXfYNc59PZsOM5oP9vUrFbqYusZWW/Em1MYx/uLd37CO2ATUK
Y9HhkUQwRzAilBqVk3FeSAFWAxWQbQJQHmkPoF+kYt+816aMaHO78pI4S2D1I5FW
56M0npDsEWLxWMhouZkjc8rwYPHVQzntU0y5E3gfoYNooTG2gs+qtW9qdSYSxmWK
Q2fhVCarGkXlWdnEh121+KPD0tbQ4tGIjI2PizpnsYbe24BJLs/cHyEkBuWk7lOb
Ef7qywb4VekTgzrz4ANmDa8plZ2YJQmSMX62E7yTe7R7MLAaAOSDhNCkqbQAAe9x
4mE9PSTIdqjMjWFYO+yEeqvHUEKdq/OPQoiblqwxy9CvQQbJci1xwj/0EdBnbEjG
6A/i+SQS/Pujvo8b0f7xIa5zOcGcAT5blIAQmsHrNwcbVHoycua9A11h3UT/QAAq
WZO1IJRiT6lO7SNEDWhfwZsSu5FYqOVy0QD5lY1nZT5FaH7KIfIO99htWhURKTLc
IVUYRHaf5LYQ6L3ogorlLggHfOX1qxMl7eZzevuCMhfGFjQ4V/OgeahguNLyO9GI
2xudOMrEkwCjTzgZtLvXkkgHwRHgOax1pazqxLLXn5bnwlD8HEJSSD/w0ETQhLiT
jj4Ga3j6dNR3GDF05Rv0cYHsFFcoNdNT9ZWTJzWHs0tjsv7gJmoa26/F5CnZsNwr
NIS4n3Q3NXVgrRVM+8qjqdnYV5KhctWgJtG/lCLz2/3HoBlolE2wuFSnIxF8FjdQ
N6piXS4fm7LS77+rQ1ZKh9CdSemxw+pzsi0rqPmUM9QGBSCU+hdLZBi3pBcKoemp
mEidTB2Nsp/s7FTfIrVN97ukar/k2lwzJXmW0KatRlDQngrqyIc7OybGxiI+JwRu
MQSnjDleuB41ao3M00gf4vzkAfqLqry6L5Q+RC53AdJlJ5SNOOjdKCUekjyHfk/t
wdbq0K17DNOutKonigV0SJBehfULbKtRG7BZxWqjZThihEgMIMtP/7YxCdrv/KE7
6lNhUSUR5odVjVg+TlD3qokxVmR0SM5IeuLkEezt4169y42mKFnfL7ntgYqBdSZI
3pykpezbagG9m6ET9ZkzkpwFMdUeZwllXKB/8/Z6Sv6qLkQJdzLlDY3KYfeNvzAX
gIpebPN1WDm7xODkWvax+FLROEGmhz9wAj6vUNxyfLB3w9UHHVgTHUvQ/YZLcGZB
Xlypdu32N6eVyaH6EKvCjAzjq57V+1VjKDGNr+pTI4gR4QdOPr6cxls5RdDlyAV9
op0HpQ/Gb6hk2XawvEknpEg4aW56WbRX3Mw1/M4oSfzUd2DyQDoRRt/TceSsFQwg
79EytZcSjIquBUPq4gwjuCTzSyispfs7K6E7XnNyXO0Q8Cuc6yIIgPBXTjt+KoeZ
QWsvWvEpT8OPBLc3qx/8vrPuQVxL0enp5C3J/fQEpIqpcHa8/m9stZ/BOmrhZC2J
QYN2N8vMGVkWRUU3ipcKTRyzhsut2h9b3GcZaSg0567XPGZuOAQNtZKJ1tGvGjqk
FKwy7kmkXEyUliweAAgUzwmI1LFhPnCO5RTP143xex6rnYwOt39Iv/lnue7BFrZl
VHVplnuPwLrroujxAh0wKWupELhJE6oKJZ8nU15vruGv42f6AqpGn7JmqUhT2Zwg
B+kScbegGDnVQPTsUccjHJHTR92Xan9LwF0PYy852VlOkcwTEZnzmhq4pbUZ4Y0j
kxPAeSdc4z0E1Shga+3EpMv6K/0l3prpufek3SVb4UtbK2hJNDF8AwoGUIROut52
thRguDr5yrHEr5PoD5BTZa6ecsVT5SurPF4fs+RGluV4qjzI4K1N0i7/laAL66rt
YS5ME7PrF/ypAY7ks3cP+ISYEbrBNQ15/s2H4FQhCjVI5TSO1GolDm+vz/YrbsdG
US9YMtTShviFS+CswuKRHptETuqvwiQWnpe9hxZftY0T3t68gREEkbVaktvoWJ8C
qrOzMiZ5KZtjfFe+G3QzruLZXFVgWTxAKzQZ8B94mCVNjvrKd2VNoyAT/yi/MYx8
q0QdExbRZbU4iogNogYDtDGdrnciXtbMu8lMrWvIFv88jK1lMJWTn/gCASdZpjkF
v9wJ+arJ98Pcgh9exhqGeFpxRM3R14JJYVKUpnqWrOBNp6gZ9mRudncUCICqBOyv
gCtKqVnVrYRCTtKAjnwm4nw3FrDtFMugnzkJy8YUtoT4IC+vNDF0E+bdfFcMfn/4
hq6ZxkNlOdpOFN+OXA8k0fpe/txfbUZvTtSbqI6e4vIprgECfwRU5RL5WZkBVyIo
Ik08aNEZU2PzcFgX0PoSucWiaWD5Q+1oU0qIzCyStS8DujpK+p8AZfzJS+bjO1dq
c5o/y6P08hyX2FIbtn7mRZyb0cSyzvuSk3iOcAGhI3BchIJHB3yRhPeHLooGFdy1
AloesaiPX6BNCO5P+/+Py7EzsEuNQiuafKeJeeXC+jdufN+tuo6/azVLpc8BFExO
H3pf6qW9zzjQJz6ta5atsHNIdxnoN/vxFNATQ3GoALMoG6kqrD377g3pf+3CZ8KU
rpd61ovqNy8Oq6rjm1NnxmaJyQMQs8fNtX8zAll9Mh4A26H1kNmWInf82G8FUWjH
9XA+ybtzzERIdSwDpNccwmE+D8DIMroEEKkvasc8uqf2XbjvDT6oUO7L9ILQcmQQ
mk14scotx2JzKC18hn1UbaAjtTv1Rfpx2FCays8TcmdPJPvZ2Z5K9mLZ82aDADqJ
US9UxYajvqXKQVktPNYO2pzwQHH3p9bANSWZUDVusjNMZgL+TUKzWX/gcIAgqYCN
xPeKLduNJdwLKbpHJ0c+rn9s46gXmA/X2KatedcVXYdbEYdnaUcFmTas2KjqBjun
wSIMD4PRg+8/aR1I27zqvjd+gKgXudr91HXgXJySDEX3QMU9IJyPjLa+vboL1a1M
7SnsnBvtw1Rl146HAC/pnAI1x43J0gj5cSpMIhqvd6esWuQxslBQaMASdmmoHXLg
jZIisEazecl81pcO51QKyD09W2PDvodQSL1QFEL0u/0rIYPkpOJJmOFc+5OrFJ+6
vMrjdAbTb9k1zOhu1RHN2q3Pch9fNVRCuXGJ85Xh+Q6DsDUmUG8J7+J99SKVRb/I
xTmjy8iaXmW1oeW6ATH8UT4QZd6KzP+EhWLCpx+wI5rreH+Fc6OzBXmLbqI08qHU
HI1ndgC7r6C5QmdPpUpzIdAZiXgYbfk9Lfss2LkYoquYMnXnO61utz63pCDQ369E
v/kFzrVmtOG/Z2vczs4R8RUVXUYdtmL0M+XI0E5wVNlcOR+uQuB0LPuZ01cEpAcv
l2cXaC1BBA4NWD6yKkWRF47tuUVbmWGIfJPihlLcTBNqLrU97ot4FGJBllAeYBBg
KHvQWoF+YYpOE8+E0mZq+CNy3nv3bWNO35LlaNKBVNbtGxXZylCpUxDMtsamXdpM
Iho0HkgvJC83dCQrToZDJs9UO48rJOhDhb26auYVrnocaWelQFUPOZFGeQL1zAmr
lTTvkSjQSih0kRqZIhMA6XI65Mt2ct6lBXcHdjbziiK3rT5yL7/fhHtUYTU4NTfs
L2p8H6wIs6oyS5SXahIY0PGbk3gkLJ0MbNL9J8I0lz6HuxRCVFzPryVr5/hgxQ7U
RR6983CYSeA6zNWkoBerB4gty9tR8uICMRH1WJvbi5GjvaRBgF0oq6xXmId3oVVf
XGlItuCjlwQDsChcJn/nYELZ2oTrLBX6ecq0WQni8ue7nFhSkd6HD4jRpVOWUk4c
BHfaqJhMTbc73ln/gtdvJ2Nt5Z9WKJ7YdFzJKX14sPD/Z/xaM/zhCzto2xbBoX8k
JZxOy7hY/XQc0Fk27DJrmpqp5c6alr/K3pJXQs+ErTgRmALrnLjq1Y+7eEjsEu01
UnV7pumXE/V3TNUPEFyOfPyrIfEiHSHO9mTTU3lJokMQzeP4uzqep4xRil7O++3n
vNj9WPez7QViU4zUHXHiYNQ5awyHSZttfXw5P9YtLF1QPvNkLsqx+YM7Xg9K5tn0
vpvd64KANGfPMKU6Q/Ip32DKgsdV+8eaOr8h31JVSiq2sBCu6eGO/6sWtU+UpJca
qoa1dnaF8EZzqbq6KzePl6rYtVlSNxrRyByvchJR9ZAU+mcQ3MS4lhdZoqrryu4f
ILf2/R2BOEvSPGmadNJcSYZzu3AMxeJKM5R0ewjK4ljKfQGz09Mn1HmBDBZJBuqZ
dEP2Dhm/mywH77dhARsq6iqNsNdwxqibR4zyrcM85OHpuMIJdeKtN5cPi6YUQf2x
NQGIIbK65DqMM/XG1J2v7Wftvb3SwVWZxT4ZShCoCpQ3JJ/iBCm1guKicTYw5gyP
Sjeptjopep2q/Uzn7sHRQ9yJJfrYiW6lk6dC6U1RYme6b1CqnhhB6utpFy+gZs2P
fWtex+Tbapr7mdlueVz/Lt7Nlh/CDVszs/fEvL7VP5u/iG9vyj8RRGo9Gu7HSEqg
0VOox7wwhhfxk4heKoQmPaCzqo4/5QCcYuWHx6Y8RG0Ic1Z/vyhzr5CZMYeVHexE
SYzp9OpwmLsAwJ3sF70TEhswlrcJqJnxcRcbVG5edb0FXZAJtBTILy2esEmoFkAo
+mWSdsmD/zrl1oi/Xq0URo7m1YYvviO32YUa0d/j0PY2Ik3wXJKtywL5JGDhEtsq
2yIktncdW6bVx+BjUHzm8cLobBMiesa66GiPR2sXS8RveQ09xYNTFnkvRAfRcg+u
Wkn++I1aynyhxL1oaGk/U7UkBCM/uyy3pieYODImFoGMvbjeY5tMTtMTeDRXIBwx
HyyVPqUBKYjGZIKbyevDvLZMu1eI2rwXnLWQb1+nGr9NhzN+Yvc/4Gb8eMZAvq3B
RokTwWrJS8AV8csUIjEkQ3TrnWQNnNK/tOqK6IkpdXC/xUDkz3qa7wp/o31qfA2c
s/rItUqX02l3D+Uu6No86skRct5iGrU3/TsaWX6DhqzITiFJPRBhKoxLvKpg1kSd
xCS1TxANW+b9qFQx3O1n+ALbYF28ntsz8UVDuV9RnsXYxSzPQZ2H+GDkJS55ZADZ
cr5kBwAoOtCY+bzkTJqqgU7KHED5wwAH0JbaXg78dBvc7jyMObI+yzpUKMh+grfJ
EeZ0kEswS9h91Y0LUoBeoy2KByMrtNEQVTMPDDUgZG8ktBvN5gurLvncxNSkl+X9
d82mHHCBDNNW0jtYJKLV8LWVAVPcr0N140nYxaSNXuXap4znYzwtnQnSETB97ooJ
66FJlXIG6NGUGxTjzNWsqCehZKB5mlbkkJU4uXc2+fU5nD/Ocbh5DriqGe2zc6nm
8tYnhfD7mlI4NIrbmZ5kcHv2WueC5c1q0CvxTMFUK+JRHO0Tfxrw8XiiS8wfIL0N
Y8ooq8IriIcmTrtySOZ5X/vy+ZCfc86mvARasukHwHYgodcoGaBskT1PRkGzdAEE
jCyigScnquveE5LrRytoKdjykAaaDMDYwv3LxSYZUXkBj80MBST+xY4z8dxtdAdf
YMUWVrTbhtHiuRun8ft/Dv1aH9xwTINWv1CgfEmJCXF4pZ9TtMaJOUGzk2vdNSwq
R1+xbs69UP795iLUDpiDKO/D80EsBrOSZBBH/Eaev7EO+YL1N0vgXOyHG/pI7aWn
mqThbck7h9gr+oHgN32MtTpx6nNC744gAXgtV02it/t00mM4ii85tqoGilnLANlw
bHV8IuiGZK5qwzVXgXAmcUNDEBomiDvDDf8q4OJUvsZEt4nUN9fDQ53IJEx7IBSA
eKjl2sSCRz25qj9Sdz8M5vz3pfs+cdHmTxFqrO4Rqg9zydggoX5Cr2yFmZ+uFRQS
B/yhshQCISGiyZvotsJyPfM4gTRYG/JNnpmlk4IAA/bPLOdW7O4NafNUUU+UsJ0W
gmQV6/dOyVVNKQQcJnZov3m0L3XH2qlvELe/E5FGSWvPC9QYEvgo2urkfXMIDljI
R1anFZwRhlmROOufMPp8he23XC+Q+OqApZsg8OudKKmGKNQoxh3pBCvEnrWOMLlm
XtrBhJ5EF6du3ad1yvHwKTWw1av1zTXkcze0k6TCpA+rcw+NhuRQFHfZVjjkbbzK
PwqAt/TIF6i+cIskUrra5j6h/gBYnehJg9ZPtRF3Mxqk5U+yFDmmi+Ud/7M7D/HK
nuJmdU/2mQSgKkuWymZHnqVBhtcJDkNGUpIX3u83qQ/q6H/Xn6tsZQSMqAekQBIh
KO22ZOV0cJYXrPEO2NlceNQXl+c2OL1ov9zXS+Eh+ykKUWM3mdLqsWX2IF4JjFAu
svd7Cbgs60Jec2S2TdeD6SCGImZx8sp8hWCNSuJrkrYkSgjVom8/ri/hMo47x9Nh
Gj/wAITBiuuTkAQ6FRdkrYeC97oLW6iitR7EugZ8lIcvwImRxnZ7+Sg5FBBU3xGm
/osJok/Qc8ZrrFOiDAnGSZanmmI3ULKOWgMf1BwDtRQNlN3cz2myBx1F1c6hn2TQ
/atdM5HEqbImA6sonCTsGXXcuhCmxHD5jvK4LFMQAuqlgS/AS9Vf/sFziG82UE2f
zKJ+8t+pKjtccxketiKDOG7yZND7cy68kT2AxuG4diS+OXMC29VfFf9v+25OELLa
Yl76rLe4J0bqDlQBVTJs5SuoZitO1LCQIsLDBaTK7c77igCWuLK8LWFFnjtFjJUI
Pqh6R2gDGgYqMhKLFgXvBV7exQfGa1e64tcVHe6JfjYLcwYqiZz/e7VHx9gLCAF6
hGhDGVzKoxUM4vkR/wmOZPXO9uwIKT0jXv1WxY+wagZaXjrEUpVl+R7578vaU2if
yByrjQl6s7JIeXhBq7zsKklKB6hciPs66zm0nLvya5G5WHO/gtjB+rrONIUJU0j7
/x2SI9LkmzlSeZgGFuLNnxeMtwfW1nVqv5o9kUZ82FLqPsUQGInq/eAQ1EyDfNT/
0R4Mk3n+GXAaKPh1mO6bhDiA4bsjL1fdkD5kY3eDLpnjDbYMiGlxpDc3BE9MnLAX
tovska7mv4snU/FcE4nVCNjjq5NLaa2Fvsy3x5rDPi1nzx2OxQTiPOn4XddJh1hh
B+oef3epdU5yGQcMeyxKBP5qlA4vSSrbjZh3SdpDzS5GfCqBK3aQbpynT5q2+uxl
DtBYUabKAoyrsr5DM/Vx5xHtWOsyrTwuQwxlthd/7wcXZKy8t6OqLBJ0i4wG7R32
mvtESJclX7kDh0gCXJMYR+vhEfmgjNARFEYo2c+y4A8ndbi68t1LPPVn8iPsEVXy
TLUOjsEEfb6raC6uVMfi0NQ4wDUCFM2E/3JMZtaR3zODIa04QmDARU1ju7vplv8f
5eU2QztLhh1dJHV24WZt8W1jme/0enCRCv4FaHhsXbGTg+N8SKdjrH+vV72peWyj
Je+ptvM+Hd5w/fuGnU5Jz6A621iv5KsTah15zlPoWnZzGUguqot/tkQdBiUldIbL
R/H0deeINgnGrS/Yvg2OK6hOFlACznoyR8GUwqw0zhyt5t16uFonzy4lPn9MQJQW
11/7oNbxsSvuLrbxAgElH5Ye55cI0/OfgzQqUOqJ/GlG/f8ZLO3T6tlNS++7Ezzj
fhdHuM5l0JO57k5SHAw4HXYXFZmOosFeTIXnQLa+R5/vNLHhqAk7F/uw201314Dr
LN6srpcRU5aUW49PzaJ8rC5j4rTSJdjW7K+NlM6fj2QrheHIaj7sWb6wTrMKQnR9
jUtheqKjAgywOxuV+xQzxbG+RYIHe+xFS766HWtijR7Slj7Fc4Wdl4/rRe0hVrcz
m958mJ2Xg/TMjiQLx+PW00Q2zJ1MafEriFbR8g17o7C0PKY0IuAONfQtYVTG7Wfh
JzdaZiIPnABK9yFLnkxypFcU2K2KW3qinIE3HDkXrevvMFBjjb6VoncxnEsjNioE
dsKmIBui7Vu0acof55yIzYa+oFaGc957/yslEgrs0MYlqvrswfui5C4pVTTnbfY9
s17nP7QB75lyyTR+rsSyfxs6uJfZLlR8MVJEYgRxeOaOLNJSQke6sBJrio5ymoc2
yLZv9NXthUU6uNE2Vo3Ddi+hzA6X+YorrRVogzyGRoC2hJPg0yza4D0X6yIvugUC
AHm/u/Cq71qMczZLWCVuAzDddx/tK2EPtLCnpgaC0qOwCCNRRD0ewONRQtDHuIGG
DQowRCAPkWnxNAhm1yt1Jqm8qDlasNfaPUDi2F0x/y5tZDEakN1l/qdNzMexrp6g
u08W+K/n29TXMar3Xx3sj5Prx/jvf3QfCMroSaVdcbSdJwhfMOV+tc7kauQaIFHI
GCxvtLEqp6VRwUg1ETx5ng==
`pragma protect end_protected
