// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UUpUM63xtZu+xsuAR4R42eyI45exKdazorXlrB3J7jLgOuQMXHDZiPHTu9vYidlS
B8fIs69i+Vd/YAHvXrMilFGSKO2Z496nb7pSQdutD4iztZq9gCY+ssOnZz2om5q2
1xbg2/51F0cvfN02rTfueQKK1WAIyooZdwB36CqmT/8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34464)
xcBN8LI1uc3nR7GAvF/3ZnDoKMrc0tguq/mtWHiV5OOMt1lhYsmWHsbscN+ak6h2
q2JdU+jAkFLI36irS4o7ysbtmMDbHDTavcwdBJWrx7XJpWub+XPvd3PHJDDl1ZEG
79D/0axzjCvpYcNGdd81DnQ2kaHbkxI+7iQjMn+ktzjm91e/+luHlnH1Ngwp7RjM
nA6KgdKTR8v+XksP1PYF3heibYfRw/yfmgJovxHrPWbECbOJqozZF+SX0JEjNBXq
TBX2MJGOuKxHuT3otg3DrgXvl1/7DH25d98paewT+T83BphfGpOVzO1eXArBxxwn
E1kVcYSMUpBHhXvCJaCCIinb7u3pY4hZ00BTs3EQjNBCKuo2pOjwr1QvBgJmZ/Rb
OZNAbOMm+GISxgLeZKbxNBiQt2R3WW4OV+Fkxxj0BGZDwotmhf7zvbx4WwsFYsN3
FDPLjmiAPQrvHl9WuNYWJmyOCfrtdU6erFG5R5v+TfUwWi6KokPfbKGC0DAe7IW5
0Nl0eOXHhZZr01+chZTbQaDZabhyxVlgge7r3hcz7wE8r13Yg+ovIjeHA57taOxF
G7NFZkfcyQauTA+v8HHYiaINOSe3qKQp5QmoBgToyCMzmnuBb9wSQAHTGHVbpSJe
hmnfP+Tq0VDQZLya8tzK2R3J0FIpcJ5R1DlOAE1BCADVZuskEEUmZ5dpTGR9uQ6t
rAT8DhZvUyBAWmYYo4pPtezHTFn/Y28Pm014cZVSu2Mj8QAK4TD/YbDCWxLrB1tE
GXe/biY6v42s/4Gu6YmNf0fczpXiorsIFxm++npkBHsTttgzvQiQ+oVrEgc7jjh+
///P5iFuXX0pxecMKp/jmegoU0UsBNHboZdVzI3FBhZMCD+lnp93ZwohUQsmIf2p
Ge8cFwN3g968a/3NWWebuS+D6O7q3F4Pcbiuh5Xp5laChIfEWyUs9RJ5LQnBUYv1
O5MwPem1xobJ7pdM7p0YE21yLz8ZbtSzWNASLwzDs/bNYWWTG9PgoDVzLGq0iRCD
12PWRzU4MNFiVOhO8I7qCa8mVnNv/msNAKXonDf/o7/TZN7XmvRpvJ1738SIbGDi
qWl7om95mGeE9Np4D+mWYcOK0NWsBGviRqP9nmd3Aro5bNCT03CUKIZxGRzHQ3r0
/AwjJZCFeP67oQLXV5/2t7MhaOFzcSf9ULSZ99y0+nrjmsHCBY5jApEIR6XHVT8J
h/Bd9qXlgmw5te2MqfhR7XD8UDL8rF2FGxrItGMMKWoU+3YdbKmDaNmGLBANHmAo
q43coP157MMOwyZXui28u/b01BYXmAQRN1Sckhxno3CtJV4K7oxRHBEwZIVUN3dP
cHfSQ8rhImPGXW9zi3Nnp01aOOQzF5p4fZRZAgr+H123D6p68Pqub+3TRb633EgU
+a2HOnPvhdOIuZ0jR+nwhDTkgglwWbDeVm3EV9o5iy+/b8oeILx9Q8PTV2Akuf07
Y5/9gPq0anWKveFGdnJ7dt90x8jPp3xrHV3s996uS8dyTBwOuQ2Uf6M+3wUwbXhU
S4Aygl4UkwukkKGR01Makw25hVNu/wJc5nBYfzMDrxynHDsPWKcxqadiuaqvRJfW
8NErH5nKVwv1OxHFWliH4dSqdQ++0WJQIcIyCie9vDNGQz1JUx5OGSsrz2HDC47V
3P3a/BOnY0tvd0HBEH3nvEw8Zr4WEaQPGcOyWNJkyjFkNpGFFC89ftInCgBVDU4j
AXMdX9ILrj5dVp6zjROSrxcBjg+zPmyzDz8A2aD+BJBE9/K5LQS6iIIjs6a3HdLE
eSj8nIW0ZsQbVBn8xP9fQ+dBBaaElZwn+aA+fjINZKgNRgdDbs04SYIwDTEPwHe3
k5dbuZ3Am0Q8AYvTcI2oXwdvxCvfFHEatCgVtTjD3LFWUxuJ+8h4tVPdYgLbvXro
8TSFuuYyK3S4flaqoxI9pOPD6RCTz+0mTcfgEPrpM8TNcC2JUKkHe9TFmMFMMKxM
tk+jPND+CsiY+WfoRgP4semNPfcM7XWIzVzJt4Of4TJRwKYb2luwXd3v8uRKNnVj
LVWRoMCVjFYR4ViFjJJWCIawP4rbt3ezXNrd7aT221gVDPVhpocUETqstDwEOvb7
V/fLijhL/VkzislaJRYZNpmeDeO95YWML9p/SIOFOr8L0GJssWRtu+cTTnoQBcsG
vvroi26MaL3u6xvXiqYwilj/EbDPDCqFYVqYyd+eHlIE8/cR7rRv/xLNyfOd15zQ
mcmHKcaxNakz46VkZs1SvB7IZuLnUc9kCHoL/1kO1SfyTPRFm+cE+XRqNxa3feM3
WMZGn07gRrrQNFy74gU0kzr8uShOrJh61Hu4x6STpJ342zFadXpi/t7LIQpZ3fCq
o0VXWQDLLFAZT4LwCPrjlGzxrxCGYCJAV+71/Mn+RS8hqHpbFCxnu58JEQdnBrqF
K4E9fhwFgNJbZKliFwRPCMfPNPtpbFyJt4QjEDgPBRzAIYxd+HesDvKA9zr0BnTz
gnWNt2vj+Q5U23qFINhYoun5HpCnLgXlOSDZwKIL86AhP5pKxEfovYebNQD4pvlR
0PXjLjL6xHyawdkR9/Aa+3Q3ziESUhOBCyYSquypEMYj94No3Y2BH6L0CZmfwxAo
axLwNvLtt3lCzuDEsavSQA95DfKvGAzEOuK7PeMR0rTv3yXgFPT9qyFjXU3u+mhc
z+GRw73iGMTZc4hT3+1LVNyqmK5rznOgRB3qz8Atj1UyiMlKyiqToe6nXVpoOYzr
v1wgsf1MMtDL6JF1uxJWJwzZ8E6C2wvRQukzOHXukSt+lb7br8G5nCmdDCbY227+
Fi7HNxOXgIGQCshCyzKHxj2EqQAr7+NvWNnozwLyZVvDdSHzgr2zer21dHENSKOf
5IMgGSmKOqXBSvvMaPsGXdmOqW+bm+Bwn4YwAx9p19563+3IvMuYyJhtHAoOSJ5R
UGeiFPSCy8U49d3wbULI0bSjlkwRv2pUXyC0ua0a7NY0iGSjjPb3GDIfLgrjZLb3
8AVpcfpeEfhTENC4VptS2FlftJkfpjJfJbAz3mUW1ELiCSwb9ew79/inUBqf7y2r
wJCOiwfAq11dLsezqAWKU2CRhZYWRQ7mXpXfs4xaxfsmlsdNIYE/Xh34XB7apS0P
Mh0oSfxs90RrQOnvLMClYWs3Fxl/ZwribC+WGsDPE/zAgWqZRbpRsXqWZc3ALOz4
etU8tR5BA62rJUG39PLXQBLQc0aDmGPFxsJbkdkbYC6IG+lpSwJgmyNlUw00X0pX
k+SMFibav0yqtfrsln2cUlwwZwgUxt3QDNPy21QYkWXDNEgszUSB0fRlqvQOuO1K
RbgfXWoKGjioP6vf8Cj+nQW5cKoOIxYaCiXopUTaf3E7s0m/pAPr6b5xSDH3jWY3
iDjSi5SLslRBDi1PNtk5EDrAxwtLN5COgBQ35qEfvBAlpbV5WDeqDyLjD3XN5TcM
PNbAtwgDwm2DwYzOZNkL2XpsLFK+azrbxKcvY8crPb61av7B5ES8s5dc0KGd4JGL
JsdFB7WLxqFkF3ovjfyZ0LO7BYz7zz3LuiXIOeKf+IM7aB7nxBbtGGmQBqv1fmCN
kv/0hdxqWjRCFLZ0N2YKE8ImOOkYzn4465PDDeYeKAwcruJsLGnEfwJUJJxCNAL0
DjiN19tKl8etWFynTxREvz3Y513GAGlRqKrbV+XPXzd+1jeqkf4FiaTu0EJJi+JC
+v+9MEYDOd8tNGMbgDPrYjvlrdjkziMVSdjXhOlX0UjS9Z8Y8ZnQ4Sh4TzUwr5X5
YqfnSkOcyxhddjj1U0itDupmo6G8XYRg4HWhdp/o4QGRA46XqPQzzHcnJiEdKiiy
lXK82NsIxmYtjJSew/AuKqN+/RGXV+FNjwqd9HFmka7QETxYptYEjpDZyyQn7+7m
pa9/QWntC4DL2Ygy3nI9sJcZLudahQWz43KFMwPuS7q83Pda1KHyV16UnFVuldFt
lYb+xw/UDDLi6+LpTN3i2GEWr8VMofmUPzehMZPo2/LQedaj+X3bGftKOCA6hT+j
2Gcke8CflDcRbM1H8Gk5uDvc3qpJ8u5f3oisFWdCTH2u9YpBbXHzeRiVov22stVM
pzKJ9kDydsSG7LdTNT4VYiNLSHH+vSaqIa/LHkb0P9op5R4RpvpylvPfQ6x/fVFJ
I6KKmWf5xkkBmB4h/3c1ZkR4tBsUgfOdin7R8fKIkgOAt5DUIczMPmul+YG8dI4Q
z+06dOHl9GVoow5JT4rSjvU5QHedyCOyOaF/ymbQbxukCHDBToWTKf7Wh1SMw9Ea
PYoa9GB0rQudJVsZORCUxc6ac9Bm348JczCNL+5aZwomFaQVhzYdr++Mx8rFxnlN
us/EoZ1JnA79DvbkA5uqhlPVgAALXDQcLkn1AKhl5yupfNw6DeYPQsVNbiv0AAm4
iRs4IwBnG8k3i4QdZPbqNlUGAVou25Mk0f/dAzHmCQswBZ0m6lY8/z1SJWAY98jZ
58rmTo6jRBHTbS6vQqS1orfkDJFhWPNioIUXiFR47mf01arvQzJNQUj8seZT7u5c
8dzP2zAoNwfPdSs7DmtULTTiJshaGeN85lUO5/EjUvIfgieemweLKAlYHS1cvbEi
es8gecjL/LtOnXcuunbH6lFK5aCdEr2S5hz4ONuBKr39OAl9vZow0JjCY3LYTFSd
M11AnYzjOoedbvgSWF+dIEtnjajw0fiac+SLN7zxJaXEsGWrbdZTBnyOjhjiiKG2
XjoNjx0ow0fCkQLL6IqR6ik9Yn5oHy/Sy19blAisS2f3W5njYj4YNgtpxFPWnENu
2GWLA7uNfZDy2FGQd5LdkfWyEes403LEnH5UJlnbWWXMNrx6BFig/1KQSjg+ARBG
mECLwTTPWEZOIphuxsBJulQsCRrZnisok4IWATuwPDOgDT8wDu2JJsWMvN452A0l
Lcv8m4Ds8ZPDsqkI7krVSjYVtEgwO4rygqjEFreXCcHgdKjs412atdq4+po/8wJo
GcDL47pHrGxUBFrUeLAI6ELit6sF1WXazpuIgK8sA8ZZE6Nq7uoqsMvCuT/Xk6Jj
QRKoHKsqXqKQxhiS+3L8lNXdwOUZT5pQidNM/B9SlRJC/HIXUQoJFy8XxV0/n9K2
xFObz0Q0RbCGTMqkEeX71ma94u9OBjzFiSv2+4GnIa9IwDpm/k8lXa/MMQAU8zTW
qW/L0gz0dWh9dqBdKeh06jODaC87jjWiWJ24wXJiWXRPIjbTm2TCDReukji1yPJX
Z+7E91VwkvTQLsOAQbf5rO3l2tURfiybkWwMDHX+ra139msmnGRi+Ek4Uf5el2kC
+u4v3x0B7hiF3COLXXiA5Wb/UmFVQCGPuaITfQoqtZpen9mQoH3INyuhjCdD662r
JGpAhSJxJKfu+0NiCYhPhDWzpo+U9rvAVXx5R99sEi2nnisrGNNSi6WX57jz9W/v
9ZIpqBiA8mMymWwPkrpEfbsVoVAEdhhYNoqYUd9xAH4mKGWxYzYWqgmvpKSuTgk+
UexayTcFfS5S6X72uePDGEOYjLnDW6e4CUGn+jHOXmYbQbwrzxx7ZKb5PVXSEVjs
PEhcC2syOx09FpJ2LfzJs1sNH57FiUOhgTSomvfW44b/lccwTpMp6ZSEVOmLz44Q
HMF+gXHTGJMpab1Ql4ihxs55bFwCTWjOajYGu856BmTJl6iHWcAezQXZMbawJrml
ZkRHPOaQtL5TPrXP/itRtE2O9Ry5c8w5ycgDXQEYDxtCMed+jFecOZ+PNCIKpFIo
sdiXtzUbdxDqqi/46SRLw2QFB+dHfES/cXpTPT1gimy8qOiqQxhWWWKzhNe/YCh0
V5hlTxeyya2nJHAsKVtdO16hrook/1yIM1Ua02OY6SqN8ufvzsy+PPkcjEuv/OSr
RbWIMfDWDgZfzbe9hBRt+3moLhbU05pW4gcQ1A8j1pAjdZvgjyWjv0XeP0G4mUAG
9QJETKZu2e8k4DGiSakbCxJpXQZ8VwVhuchVqDn6vvSeXtoi9ZNCLBaCep09UogR
o+4L3f629zg+xc/KepHoPV4xPyRMmUmCMmudtE/u+7FDJKleDdX+JcLaIL4jwQaC
oOgJcQOTnEo5HorRXK1JgHc4CWH7EbrQkAATcDtx+UwGndsup/pg8ndQg7UNCZxc
E3fIe/PJUVRLcLoYeQhB8beAUvz+CYFGqmyyLMtLPMd67lnY30GV/WwHxJiuFQB1
56xFcLM9TmE5Bmq5h7B2TJobYloF7H/X756h1foqxacYzpAmdglvMPkkq8HPwgvn
bWxOoL12DZ9J/KEgwB1dVKemkr4t+ulSpf+huROkeGsS9Lqc1uc3oDvQNET+UWl8
ObHOn0gaoyMM/ULchWTqk/sczKeKY58cb0cDz0sND8/xsYnDoEBH36T+lfzQungM
nlvq+2NnZftLmnoPaFI6moMoT7+Bj+OYRcWF+/ybwZDbYsv8XPhcWIpvk4/0DZRR
rajsNMZAc7u9eKklwiDmGwhfAp7RF1MEXDTwLdeQ9dhdT4WOFnHafkthqmvaFHtL
bpJmshLMdc0Yy+egU4if7RvfRFhrm5RJ6Rsc06Ln5m7985h2NjFKaW4rCO/qEy8M
r5BuwI0Tj9b6S0Wjrz7mypCOCGL0fsUoAGpbEa+gIka45IfzF40aNUEvwW4bGpuM
m3K0OkhdI9Ap5yepqA4qkr+G0eneTdCc9tjEukALW4UNPOdUcKWZJpYiqWdFOrY3
q0wJL6bFsKNCmg7MOL+ytMTXPocPDC3qOcrjMFMU8fi/7qlArfidP4W1CsyR7sP3
WQnsd3zinocD4msCfAdujBN1370q4etbLIy17TPPd58wNN9rTWlZBTpD0KNRct4e
+9rsAlh39qr2jJjUeuxnkpZS1L9jIsJwiINylUP7aTz0xQXVKcV9mK9OaGCd9imf
vd9X4uGMEebrNEind/Jr5Ix26EFW/POs8JWdCFxiBmw3ZJP97TTyOqmWEIIzXVT6
1D6HqBKK8+guHWH2BhqyVk2a88+5LrmKrtNFVOjfQouzO60o+Thinm+bwl8/ikJo
QPSCwavfUMIUG7imSipoagYPyTEw2Z/m7Cr2+tdlWMv30XGMkdVqFakN1yvwPGxq
9E9HKZ1JoqTB52ekfCwcggkeq+Lvtn3aoO7F/5IEJYCWgz9F6o8ZqA6NVckAsa4q
eeFnaa4asq9bEpTOLTflwwUaF8K6mhfM3hxH6bflJwpLiV5cJ9+dRWY4uygGn8AY
jyJZadJlkQykAc0AarVVeJXjZzNoXRS8DrPQeogiVARsI1XCEhzWwMEZP5RNBmu3
RgDGmv0X27T+yr1HuaVQFd5slm6Spya8uUF3mPKKLdpWh9ytaEHHY3YzZkheMmEa
sbgVasibxQ5egcZWHwSTmyss7wHJuOYk/AlHTG9jOLkw6rf4n1eFlbH5ohDruOdF
56zUREGq6gs5oAkoVPTZ0I8TyJmHeO0PnwFhC+TCOjnhBgAyLxSaZKb9liHSaoyQ
XDe/oq7eMtwJ2DM2q2nH8fHijQKMBYH9jvSKp0hzcoqIziNRg8AwahBkzRv6dMHH
ZKCm8tulOvh6w4Rn4Z5YUGp75pqFyog+IgfuwpI74A+7CL4US2l9pv1O3f8TWkDO
Xv/mamgq9LYBq/12e5qsl6+MyUpECLIZPKEYcjYEd2IlKPECfZ4zwz76UktUxW/H
+P+XUVuAujtZFq56RGovJ6d1YeK5OyGkZSnuhi2DOK+0QF1R3a8+J8vkwxKZ93Q0
DHcG+KT/WzOK5oMJDjq8m53rR8kQLsOVWcOpF8FqqVV5USc/WFDC55kyMC3nPtOT
P8FS6G/rn6Kp3mGBa1fFoZXG42TEdD4yRU/payTK8K+i5qbhXYrX67CBl91G6vlR
JyZX5nNrAgYeSr7FVhA/GNSseQ8r03E1wJHpIFHctI76pUbl/45u0lrTMIW51//k
GWkPCKGztm/NmcEz79LDa74OgwSpDuJwzGnMUYmHLiyTE32go1WYz3lXS0aj7pTg
zVQqvuGUBvE+6zUyOhz4oQCZTzS0TAWtBgBAiD/zNx5fP1iozBxqSLUCw7+ljRQl
c2IH84sfiWP/UVQiWdFgd2lJu/5PWdFhH0WXxqq7IbahmoPPPP2mU4myj3F0oocy
n2+02bUfXC30UH6N5fZEUl/eRIG9AThC/OuivilQErXJv5sd1qXsVohSXf79NeE6
Ll5qs4TKSGAdR1up7vi8JdtWS2qHkUOZKgpgdMeCl7hl5LoobOjS61T1yCmFU9nG
6MQfZqZU0CpmD1z9X/z/EnioYMEBIjGQLuCuBt/tBW9lPIHV8loN08acgQl+7ll7
s/iMo0lBXa/61ysj+ZRjkLO3aUwzQ5gvhqdWljLeA4ALhQ0tz1Z5d5xxtsb+taBt
A/crcnfWo/7Y7w/TdNX4tHZz+seUlysNQfvqpzJeXhJ5vENi3N5jwZcirIbvR/yC
slMJCpPtk8V1lghk3IHIkmd0MuR7ZUeHkVDTXJth5o6cDGxrLoHRVfRRMqGcE1hb
FosM5wq6EpsTJUlD7NeH1oDoix8VM8H3HgEoDujR33Da2BxmFDlJcnEZe8HoKubl
KP5CoCBHvil7ujgQZ2TJjjHN4yhIZmUzwQXDGyLvLEB5FTvB3PA3N91c8isHdS0t
axdVTKinO43+bnmpTRUV6DkEcLXw5fjI23FFoPhM0tXe6hwkpyVOtIXY1Tb9YaL+
BM3Yh3YBUrRS4zH8jxiKNbg2SJYVe2vqwCmqO88dvJirCj8dBBwd0hKXEfFYJCby
WD+fWMfZbNurrB9Yj+2jaXv48bs21HUDzJmPmtsm99stcERXIKDhEXIKDVBRmnnH
BvZvQQHSl5EX7bRvCCQo9uGKjNjuOGPMeJMXriJdt4+PT/8fJhAnQ5qt2NcRNMJ6
B9lG+pPpE4tqGzh6nV/o4ZADQnZSSlMsFHDSTma09YkIyXkN5kPQNvbEGak19BFe
IORRJAwjqbBRLgTOCZvKREjTwn5VCfRJGRhUHpn+IZgpyM45kDBpwsZuaXcPyjgL
PoXI1K9G8xDEUVCV0HtKcU5gdrRthyxchDaEDEve/opMAVeSudjbUwONBl/WVBsS
a1D1hyWpFKF2QHUNLzbvp049bdmK5Q7q2yUGCHfbRsnBUkS3Im7dxZFqxM+Y5xvV
+uEJIHkqpPays/mJXvIfevkSY7j+g81llrKPTQG9cz0cZ4Rd9yKIWqMCkhDwAH8M
0ZPhyvIzZDSkAAX+FrF24h0ZrIKYqI1U9sEB12ZtGBGtnMHTdbol89/BxuU2EAfs
7DI3LSA5zohSQLd5XGLA3zh2xfU03T3gStlKCDOj/rAuq+8V9NkzyP3T52N2u6Oi
Y1lW9L0dZ91sHYq+xAnvDK+xX3KEoDfUfUQYyNh4YlFVLbgBRjes1I919xzVY0bZ
AjJma8ai5SqR/sOjgwkVaLpPbH1OHYqfbt/F+Xk9Tuyrlu0DtMffthKMMs3LOtr0
ISC8tW1qSYPos0d+cQ8yvlMoQcfpiwrTPOhLZXQvMNrDr3SzRQ1K1smaJsEd0MJ/
e+knckYxs5ntu0B8fVcgFOXnt5dKbO7sqf+Lvce6ezTbddclMM6iCUNDZKXbpeuO
GPrJcZMRAqbpi9bpIkiN5pNAhYmC9+00GtRIFvatlrtivWoApkotcz7uzsm8UCVy
jILzYlExuCeEEVwZtB5CIcTOkalbQ0XrYCeB5B4torxC2O9gyoSSvElykv9fH8vm
MUMwVTnYUxOXrB3WYVRcQYF/bH3vlIL4PRZxMViXD9nt3upcVrWYS8Ivk7M2Q0sH
WWOVgCehRvW14JauwUbK5Tgtu6qqNoOHFxBQOsUkYVij3oz1VqLuiyHflH7lR4B8
5me31o2hYhD2YOmGsA2z4fkC20rd+PtYEN6aQo/nGrajUVRKXPneEHBljPc0prA0
1OT5VWAu6992htWu6UJ7oYrBn4A8CHE9I/2vvArgqZQj2sjlbTPCp6nTYV0IJHs0
X15y0E6RnmrHGgvOPDZId9jsR3HxKfDjXGexWBc0qV4qvqcatZefNqi5SXuHfHiu
tjD4kwcEJipR1Y5g9FdvOuJ07jmUWLZeACOrG6xWzrRk3zige4syVcDHu9h3W676
q1+2wP8o/Kx84Rz+aiUa6rUY0WDuLqLh0HNCrHYhEB1hd30alUJUezMqLT1Ivr1L
F57UluxKvWpjezNVtO3j1lacFHUm+3vVPNY/1FG1HdPTR9w5u+VyxI6XB1+6TNzJ
SuxHt5x76NZmldBWL7c37alaHijxi8Uq5fvQ46pWdwFiqp1LBBhJDrhDz+THH58j
spuXpPKmvSKiNdEjU+zhOC6ce6mmt6zQo5va24qWx2Z2J0gGzwVtIcXm1xr179ZT
M2zkPv3jlpaBrq3iPuAMqkb9PRDZSj8EesaDvXbZWq1MkqEvWjxjQWZcxhmY/C3x
Eha8PH1Mfd9nK1HQNuarf3JElizbaVvN1mC2LaP0a84DH2f4QDQa8fcieHkyIrMo
0CTnFO02c5urLuL8GrjNczKlxWjDiLYHtR8nkwJ+1Rd5xYfrh7/vbhGgalI/EIW0
9QIRToo66k5oL7caR3fO7GB/N5ViT7CHpROT0kgTAsybgv8q/8/nGXm5M5kFdKLq
bylsnShEEKVyN3+fTntCUXJmoPr7Mx2jDuxwjMhPKcTd9/lDmyHFDl0H3EhySXrf
GumFtuXdGtuwYtvmZNrV3NdwTPtCze5BKM4u6Uqu8RhQC2K5ydhJoVxDUd7a4dIu
nT2RTH+mQZ2DXUEBtd5vc3LFqQD4dIMOaHFv0jXJ/Tg8YuzSOe35WtZTJ+pEEp/b
SvMvHqqB7xWlfG4+BfEn5xjMrc0BOOLfekDcYDCYrXV0tMnD4zidL5Z5A5DxdwuT
PjPRLzm+DIUS8ayRSRomI6vD71Drb4QAXQ259CMGZdCxwjGEBoJNqXNCOyFJPf3N
A+4wz/+hoiF9c3dzOw4aTaPTlT8Z22yUku2khBnN+1iU8bF4s5EhO4WzliRSzgIe
gQmEbkTSNeNnKAEDUzUmQyL4eJNqPpcKh18kJ3QyathNeMs8xqZEc7ArpxHHiGF7
f5YRYLMetlhapUpSLuTk6jtkQ1nqSTsSztRuqXXDdn4fN/jPmrrtG0zZtFp+AXQi
mg+ihhy4RglgDwBXaVO0bOqEw5VJNVeq3eAa3lmiDD5Mm294Ac80dQ4eETpNOLxR
Y3z9w12hgvbz0IMHam/hVz9/FQTl3MEleyeAh4bfSBIFrUoRm0Ei7NFKtsWorTzC
Sz1ljRKaUblFK8bGtoJRvW7faI+rYo9Y6/fftH4AP2NtrMTxO68Srvi7bfg6uYy1
dClQHtg57RIF46sMzao+VyUYaD2RrXb1AfB0BfjtTlX0x/P47czZxzxcN4TkIFaD
Z1H+KBuwW8BdXh23tJu6uBfyAfHADXnwG0jDjImDUmKpSDzxHs3BKqpUcarS2gIp
RZmYmIoYifEr2MEcuMh38xDzRUcxXfMHTBoa1J+zkm/OOJC45z7VfDO/8wxI53SK
iINukzYDK418lfayz78PdUHlcUGOVXa5PKvlsBlo79pI3iV6lWUJ6GnwlW0jhb6u
YmAij8MoMEF9kkrZoeeYJuNyDKbfmK6NA6NoA6sb1J6pVFMS836xVjK5Wt2qnMV2
fz0AHvnE6h3sF5ACn0s90pboVbVuYGuoyqyfS+9hVpb7Me6NX09b6/Kz3FAv0idt
qsWInRTaKEQAqCGwv17QUnsOrVDn6ISRQS2tRFJmNgIrAwDroiy5LGXZL3p5R/yy
dpsThJDLYZazbqW86vqAegYO//xplRH6hYbijXglYJNz1/XHhnK0LVdRQTQMr7YP
NLt0DpAZTwzQgbet8DV0vNGzKZ/E43us3elC4Ynco/enEM08sXBe4F0RkXnxQZSW
y+iFnB9W1wB+TGqZlHb36DbfqeHvazmNWgMNxFEbNynM+Ghka3OQnG+zKg5cFpUW
Jhpv8rCBO8UaEwB9uzbNOscilZAnDs7CUc43qxwJPoHm7YXvZd2agWqciFvku83l
55z5/63uu8v5NJNs5D4nxL8iZzCBSf0y/CCUJDBnbIaqwsnmX0UpM85N72RgXycC
lCXpjH1S1Tf52VWUP0kDQSWOMfHk7bJkWpl41/rVL8G5Gar9HmQPmTl+TMhq3Thz
cvhWijGJ/Dc3D1V+p4FpFSQB5J5NVNnB2iGD10FqAu3W6I05oPXgfQBH7glhXuCx
KXOH4BI26OnhWcZhivY+oJ2MqPUEZTWzvpPFjgZUC2oz3uEel9Bi9Favhmk55C95
yQoi7JVY+OdGnZYZRR0BGGYjWAsag+fHekUr9DuuDvUsOohzaLhAPASxvjzR6CmJ
ayr5U4vJNtu8z5E4ITPQ7h0omMUpe1LKkMj6ffRlApghZyoGvPNC2oSEkAa0BJzh
c1BgWkMAZsiF3QhQ5Ts4U5tirIdI17oxbE2dhKkKz19uZ/YzW3iJx8AYKLzFO99H
hESxqZs2Kqc7i+5gZdgC+bcB5HjXL2bsY0tVi6/TZ1+vQNBM4tJVkElEjSBS0S8i
uVh0agrezWTRzJffDf1QfAT393FAjbWXHAsgBd51OYtWQMB4WVOvLXqzvkOk7NaJ
KiQ4UqjWWindO5PK8P+SW5LuW6kGJhvWXakO8ZHqXfov34IHnkjnVJX3FF7dac4q
6+9r8P2ZqqsV+o/f3O4n2D9zAEochR76ibltzLmKYwnaYxYqUns8byhDOhK88XUe
dedKIcLjKOnNFXzMqQDE/2ea8cvvXvT9BWReqkcWdDP5vkH5rXqC81WyeIzoDz9s
2Z0sBtyp2aiTqi6Ek+4d/up/tCw8t8dmyRYPqXGrpT7MsQcBlnbMaT0Q2DlY4ufw
hG6M/tw+eUJEmuU1GpgHAGhV8TLe/Q/M7rIuPUX+bbAI1LhqSVNR0PU7IMrWzhQj
G2jAXE5npQ638KVE+t8xa7e3jgYSXkGYpL4puJC2Ycasrq7eVsjO01wwzCrVT41g
jhREOUAPnGyjActJDVwmVHIRQju0maC41UFFCNhrsfK8CO5TCqaxRHZjt/lPY32O
sgDWxhyoJVeLWXM7kTiG4xGwdaOt2svVvymlrvI6C14VfAO7SWQBPDOdFLqQ4qgG
Ne6pCRZu0ugBioDO08bc1fWWqc3NBI/0cAa4IC1nwmFM6Uh8dcbD5AGFQsWOeREM
kUrxeORgJW8aKl9S5egOgJoue0+/qT1ttA0bKtv5gpL8n14AeSTxLvi5N3cesHkw
lDrKZC+asDQbJW96zgjZyxvXiZmQLG6rHNFgeiqCXc7ioxdpN48XseyftjdYUY5X
CCXIZSCNNKZxkmIYD+luBi0lq9xArz2JHadT7jWIS88qtm5vVs8j6eGeiU0NCLyp
TNEumGMJrBrhkZdvY7HLB5u2PG6QlwqirXnCDzc1mk2uDXt044HjHVTEm/5/hNF/
F5RSa2ooHt33eQfIp5LbPKte/kNimM3wHONxdldrCRTYQPMzHsOS+g8SwIcnZP70
bhRSDgwVXlKCubLMusDTpw2K2KOLBTZw1e8yrH71vuPzdd11VncwB4qQydiDkIGA
AcRHbH01GJ/ydZ21sv8MefOmH30KrX1t7lFYonVRGwbQx7GB8xEUvid15DyOpSIh
QS/Y3Fhx3FrxtwC5VLWqQ1Wg61bktqLjATrZvEaycWwMvu3PkGfDPh+CBdzP6TCZ
AFms6dl8ZyLosIZFifQWnPECXKr5Y10LbJiawMRaGyhRyay1v5Mx7swlTvfSxfS+
G/bb/edqQkck5xAJ65hOds2x5VpoQjKNN/kAPHt7h3UJNWLHWWQEZRv9jvouVf7M
LSxpZHLuCF3P3ZWRD4K8mw9rGiVrCv1HPfr49F/kdN7mlO70BZOe9WoqXxdw5iMe
JivCkQuQwFXOi8SpPJX7iNVqSak1Si8TSuQbR8Iu8w+KKGTPbft5EZocg0Z7K5ln
ceVBTr8a1Wh5axhaNtNwnQE/pN1nb0J+seiN/B0OxCQiDJ5uwfv3MX9EXRDy49j4
l49R0tqU55GURPauCkUTLzIkULqMz886DCMNhaeM0ndL0jaV5De+QLMvGBtV4Vci
kKSqK7fDnwjHLaywnSgPwwRGwQsdECRu6d9eNuRHy9rLafwpLGBX7yLcdBI4hkQj
jtZ3q3pTUc2+CYG6+r4vWmdK542tHnS/cig2KUYoolqkporkj4u9uYreb2Xf0Kci
sCWjwWj52mFjiyOSixLkmt60pwHe9QQV/zLWaI7XnnVIKoUy0WKwasAclp++81k9
AT+kcugywpisbzTUMg5YpC53aQbsGZRZA0MXDPiuJchymOKpO8SRxNFUYtGJxcME
a+i3W5HinyK0I8zydiOLpE0GjvlKZxGwxYUui4EydZr48eLmncgTBLnuNSZMSRz9
hAuWVT3iXl15Z42AziiDiOW/26OHN+qRdv92rxQuteJd9xETQBdiCPkzfi5Cf5nM
Ae+uPCyZdx0mFSHSesYljaxr1Qd3n+j527EZ1LxCaqCtRK9kend+qN4JwWR4wuZp
Bjh8EHsmuu5UqQ0YyNZNgypVLho9d+/kTVrauv73mzOcdy8t+qTtlTMdLUwgABSi
vf3azqAXIohUKkj2IBKtNQ1ZLfkYnOPyQ/9oRg+GIYUdoRTiZNXyvQ5j1+/SPED1
CMHo0iP51ILg8jeZhxYg8V0QkXICy9OSEMq06E9qD3Pe3B2/7G+Ta5zqTch8CxrS
5JAnufKYRrSHCzE8H59tVwTwYmi0nfG3VRV9AP/FfKoGRS8VNJwdIXRIZuZ2U1Pd
7XdUSBFJhnKGJC1LB6IQtDEP2BptiQhfFlinvjc9CFhQh29j7OgPmKyvfD5VRl+v
fVGn/gWZ7feYUiX7ai4evK1v7VPEZmJm/jN8tQT9+tdTUcc4n6TIfNBCuZ7y9P8M
rTPcJQYOYk1z84oPJUbFUvyqhnnXCDtdwbJ2s9tyhO/6iTSkyOf6A0J6f/ok3OGy
zdiuYLMOMqu2MzgOGPMK31Sq2x1TKrPUTwQuanIt/7XHLjFIHYb1rFz1B6DYjrqX
eHilwzZsZ93BYORivHEJEEnuXwRXXPgNs6ChppSjZt6kQ9vf1OtGvbruXmSZM0o6
X6mjrgsi6qIi4RrSTzPNfn4f5pcqnXDlGK1Hm0hBNZTdpiYmteOuHUybRKmO+PEr
T9+FNnmjDU4c6p2/XehqO8NC4nA5jUgtlr1WlbEV8mjSGVaTCePXVnqfxWDH+HXv
Vo/XcFk/Dy0U9zm/JreGYb0RSIeD1c0QZa2HMNYHyFBgXn+184yyofeQgzaXRnup
0J3isGdIjuVxglo5zyGp3nMmHKMUVK4/5OPn3Hb68bf9YVqJ4usaDiEYpoPKWmzg
KFU0tWOKBMXZokCjDlmDTOBdt731s07Gahc9yNdoLRqQuFq0tXtfmjtq71I5Kagh
xVLfeCD25pe/j1vzPIOSeaxyrpP8UpeSuAHIwdNLBhRr/Phr5lgBcnfVNcLKIjx0
2Mco4eyAKkkzmT+P9LDGYj8TX1qTWrUEKtIKJ1DAhV6O83Xw88WEvNgPcVfRh5Pw
itCTAIHZ6/fiT/1TgHKoKJh6Khq3U8z73Et+IB0xkfodqDp5roKqHmqyXBgRLUbq
j9x+RNFVokbiobKHwXxOHG0L7y9+I5FF2ZRZnFBQKU8/HMnHYx0PQBuUNiKLORuG
4dAL80fP3oe3WnxPaI2kWbGtISCenspZKUvruVOKwVmnOss1ebpBX30nQWFNWPPr
7W6DTM16FjpTzZeR0SkbfUWUTHEWsUxGX7bbb5Vmrpc+aT1MLBhS0G8KC9YYJ84n
a/zY+GHn2HILCsebLMPzpw9U3cmwdsiczz8Vq9Mc2sMpLumyiGkUeURen0TffCXB
rOICitLiaWhxGfzKUE/9sn4BOdsj2AW4DVEluJVMes9OUZEWKDDp9MJ/nn7tEseA
SiBaS2lJ/XHyluF76PjJ6OjR+r99v9CChMuyfGgtiXtIMVD183CTYdwxeqQENScf
QbN0pY2II3gHdBzEMQD5Z9ihe7020ZFwia/q2RZVHlx65lbgZEsG2RJ8ZsTLsqmQ
y0dY//uW6cKv3muX/L5nHSsc4sONkNjb1WenJglLRs+eBxFi39vE43ObzjDLMakO
m7zpWI9nFo+egajxVGxuNIeQxqMSM+BANLtczAXYPJTkyLOPKFqyXEy6teqin/ZN
CSp7OfkfvvaJgc4uZXHFYfiy22nfcikrGaOBcaALm47C2H9TRIFkfSgjhsLcCi7V
i/mCQ2QC+rU+FT831/DO8VDLZUxlXJN8CRuDAiUJE+ibOVCqFeZX7uRqqsaY04Po
7E8jtGw7+09qS5ilvwV1qqjJlwN0S28ytl6NdC11G4PfdYFx1yVq2W0Ub88n3rZX
lwYkUabVRzF7gHBNK1Y+ufoaVSHBY+ss82r8gSpo3Hl0YfkkqMdKNyY/f0rOd7qD
/ZPuUVbFiR9H3Ftpem0OZaLNdibvSMjJbyWWKKUMcfgeoOPB2gyQvHOc2poWCB+X
K0NnOh23q922/WeIrE0yr83VaERXJ9oSdXX7r28A9tfrIjJ++VIqvp9cogRmfPFr
+WAtun7DD7HiBqOBLXkaxJ/O6GdSEb143i86GdllsZEZFJdj6zA1/eYsZxRGuCXb
suQPJyuXqS5l1Z1zoOy4QXfFmP9GCqIiGAPYiMUGJ1MBgHJ8qSzwftbORsT76bls
cunz4WDB9VO6UppLMjNPBSVoH5IkMA+c5cRRvfRQkAqDb3HWJLr03NGI90GCyljF
mzxFP5sZ8ScT14hvicgFJ/big+w3gk6hFm2a+LqusSqkbLrQDPRrdclM47ampGqg
GC0tWz67Ztca2hN181CN09BhjseQdJgRtB6k/I9WDWXLCKltq9TW8uUZkza8Rv2i
88zTbBpLjVRGS5L4V4p7SJ1ird8okl1cXm02P+U+8wStUNolufVQXkru+bJ2D/He
7wqOAvtXsdT05B5FtE0ZxwCHEmtsLbrMkGYuPrKwopfxElYBn+dI8mv5XSHp7b/R
qDONqNEMnszjCn7rJItRFkf7VPMVZuHRJG/PqVbQy+4o7cRsO75prGrLuDgQGLX+
9aY6TE2NvdaXK5Ycb2RaEIdOsJLCG/1sySNlR1r/At0Qj/DMn6QNoPJkMYyEsKiK
qbv0mmLWFl3/MTagsC+9Hu26vPoghp7idGVlJA5BI7zZo0EHsh9c6ibl2YikMZQy
OPifQQ/PI4d89TJwKvEtyNbLmWtAYl9DlPZWTEoC19I6NCVXF7ZFMcMkCqip/k3R
d8oMg1fEistzb8nY9aUXWaLPIl/117U6hU7//T/iQ6hlqrv+shOXF1s7/zCj+A+Q
PKV8AMxuQGsXmDjILjCtROKiDkFn8jqAWK9XPEW/h92uZ8rdlDENMPleoVmTCHsh
VLZIioVIEDy9UO5EzN2UGm1l8YftlmN+ik8IgC+386e2bunlf5JkD9X9toOCHeQT
IElV57mje/rhSAt4U/iNDNCt+Kwff7qiIlhxxuSG0L8YSNp3fi+sRwhfmjaQcWkC
v0shFSxIR/3bgswxHUEUJzILuBuCDfofiwIpZUenSXFYMC2pm81zHH83+zRykdmJ
aaLW4Z1vO+vZdRfM9YKIftli77WVRymVIlHxlZ4nG6W/Ds6XqdVe/lAbJ5C7SY46
cRE+iTfURCBaNAUzKWMHapTiCDeJ9/xtCf+g2e40YD4TnpMrLRb/ZeUnvFMXBMDy
nTcpm5yuoq5QcUecDm1FdUFAJqQIEu2XHfDkpCRg+knX5Uwb/43Y0FMJJpJxTlSa
R2OBvwOwIyI953Wki+V+lJB/6Zk+XfwxKU4BWkDpyiQO6Z+U0CKer6cjdGsDterK
6LRMujxgj8KeXsKwWxSeTILRTSkdv7X6NTP2K/3sPHD3S9Sc1H+l0FF2mdyDevsi
IjlUeeZiMc9sI/W95jOhL8CUnFkxxgBK6zt8ZVEPB2OtvFtJGVwFbkEJ8CYdltmn
86gatXI3gJoki79F1k05RNSISvO+fWJRuExkL+s//auNk0TTGYfqeI7L+zYIUe03
28YWXwHIqrUNznBEKwS+AucI72ocf/Ft8goEwrAo61utU03BNyeIzbXqNc5Vm8E7
+GCHKQR5K8OfqR0q9zMo4Xg3EQC8qefGJbx8bFEH9wzA583YfW3prXJhYctUuZQK
TS1/2j1KZLW78t2eWOJEFh+Aon2kRmiB6wY6Ep1BmXZF+zl3StA1NHV5A0jfxsl5
XWvlq9AoYsteXMJN1QqD34A35s2OMOgXnj/CfnO8Ak+dXuaK/E3DnlGqj6siS5gL
vqUnYF0yjX9zSsdqFNXVW53+dxpPNWRpsvGth07eg1F8etWniR2anPz9Hkw0+HHh
Mm5MIQHs+H1y9EjVzxHda43HpBV/Te9mgw3eQzywvPiBnW9JwnXd5rUhveopIh6h
WrtlwiOgpm+3E7nEwF0BfnWrG0s55+DjVf/INRFaUQwoFJYAsN1NEWnH8G0AI9Rk
c+yBaCUemvGK5zLvO+BbGWDpC9OUmnAHk6r570cvBKLc1gxb4WRcF1mmduTnwLSJ
eKeaLg1iz9WOk6MdEas+boRSCvciObo8Riyizaxh3HZpmqL7Kjm9IBdYroUJK/R8
Dua3dX7oj5k9dFHXPGPal2LA8XB/vfiHCCD6Osj3xoQVVf+IkwLYiZrJeG/M7QqP
hW4q+wr8WRTww2J5hfR9zAmkYxykNEqGIhOAvuR64ls1qdwcZV1qhozcUUvrikPt
XjMw21apOEneTQ3NoiPiLO2FRU5QN9DcvLbUVQGNDaFL/eZj7ppn7cyR+Qhi4i2W
aX1icWvx1jIKtWgQkHtRjNFIqblgqIwMPuQwCyDj1Sp3vjmMrGQk/6L7+QwuhaHl
kJ3jiNGvdbt8dSZZ+eNOFlzckFc5TAzsl2zvJBPOVOWT0+rg1pA2N55O6iINTkdi
M0yjxoc0IS4NStG90dqjrMSi2GHD7A13Kz1EVsZly21mw3OKXuznWeuvWp4Z5ySF
fK2BwsLrAqK5J2Cp97ZAnpoP2y52KcOXw+NjuyGYM+BkG78cQd2JJFiK7w+QojIa
Lwt9/OB/DL/+zjqX6lzWYjlUTf1H5cnBgPeMUvd9eA7sf1PectZbyxnvlJzFdv0T
aUeiyn24H3SVWdTUCRXksMeoVzOsM//8c10hk8EE8UPku96TVWKmcovs1s1Yyoj9
ri3O/cfNPlBFrWeuY5hvbYWEXEa/B9Dj97GLpApp61Eow4V6Y/fWsGhxiLFMkajN
NXmOK/J/Fj4jAQs1FKlsENaU6/N38SXVJhiau61ubfjZXfxbIsS+yEkhHV4ue6Lj
jZU1MXlSaBZZTcwbWwah46b6AJphk+Y9CUeMEUZZljlCp2aouUa5N2u+Y1NJrDCl
4XTjuwF4IcYUsDk2zytmv+ByvQxQBPpSNMMP1d11Eo6d4y8Gs2FYVdj5/+ai3ksI
qFBdeKSBzKcd6DPTFEuW/4hQN8ePil5iKvz7D4v5PIl+FVDDEQh5Sr45QcdKzGzX
dSne5RG7RNpGuTPaYcA3fFhDfKkYX4F7+J8QQbW1nk8+F1s2q8NXhkpZ/t16d2hg
vetq1jOgHno8dRB2zY4oJJoj1asVZwfIPxNkXfZDYpczx6gkx289CAFLx8XLSX00
p9N4hAeI0Kt1lOucHq8afRMchpSvmsuPX30npZ30bVFem3MHeHX94CX7qMlnQGSI
IU2EGpO3dTmH41z85q/CIQSzfZ4NyGMBVcC//mFrs8vyvdpav3kd4T8NRQy+DUp0
qEOVj/zF3YdIidR4qniXF82DWnRrYiapcmdRZoC+xLo0cEX+pURzpnK1DEQv6lMy
9BwmduxE6z/1rNRrt8QJQaGjrMV8ap4iQuPaZm8wXDdLjxkpEKFCGgWDtuINcise
+D6yUMxMtzNoHPT9u0AOnwqLGRUebpOOoKevgzNsx2e+niWW3nSWY580hCQpt7V5
HLJE/mXst7UGp65gnj4vmTsvCQM4IkVEwlhSKRv7qxKSaBqYGUyMeykRyKf677dM
vqfoSJnr13ipsE4bS0kE8ba+wbqe9d7zaZChwPWa79FZb1eACQDtmj8t3qI7tZ5s
YQIeTfiwpnXuWCv+oCKo3+qzbYDwK5cCKTphG+SHyPp4EMGNjdqrZ9R7SKQ9ZF7m
lfpDB6tFu50a49NrRPndjVkElyw5wv4p8dsXLK57/kPUncDbwXK+HdIPpeOstCOG
0x5cc6luoCA7iVYwVn9XqYPKGBHPsfKafkOuN23WeSu/Rm5/e7WXYLzBDBKHmRI+
vNF9lDgycwNy+iL5vzWRZ/M6ooMepfvbb+Yg9diOoRIVuiXstTCcZ4HmmjHBwpf5
XpQ9DfvxLcDcuIzN+PICho+XiEresszZXPAD5J3USxqZcSmxKb3RD7f6HN4ziLjD
9Ymnk6KB5vUTrCz3wqskWvpqZnVQH4j/cW4dogXAa7vQyTiJQjoBoyNUuVgUamM5
INFDsIp6BgongQqMjX+P+Y22SnV41TDBMtehq59BUE2wbZuH6yLfqOHAL/9VLTGs
nrCPUNn0e/c6h0/ZjW4fHJIaCHvwB3kULeN2KZ2j381wlhrzg8/REUKNCKs9h7wr
Mp4cxvIoXuZg7gJqlUvamw8rAsVqx5+Me5dg3afx6NWW8f13De96vJboBS0Lg0LR
bp8LnWaD/K12ClauFrncvLv77sJMtV2lFcmyOoIw1E7XqOrbdXkDO+9XXnSQX7Oj
Soq1Z7ycucktMOVgqPu42qUT3APN44NNXivezw0KY2APgRSZ++tco376AcyDuW9G
gygkCyGldAYUUoUxJm99m8UaT2bhTONU4bcsfjGIvo1qjfgCBLCkT5jp7N4Q7vzt
artQRx3RYvLQnb+XjFzEH0cdau0K8FQyoKSSKl5Eda/aGbM3hZfAXEwEGysZFxez
rxv+lXjgkHfvZWuG9Rz0oaYHClxpvMGhPPd3KzbdPtzKoP0HWanJh9LXRLa9/Rw+
+C5lLuPqobcFI6dswjqJpeVfkiyBw98yIDjjWUJC1fxoj6HsrwaG53v3vppzbp+T
8SXbVOz//XdWNMnN9KWTNByvfvTpAshiGz2LQN0g5eQzmIJhZDTnXNcPPkJNTPKX
Fv3vB0NGj3tzjQUjqXEPZ6wq8EfWlYk/6FatZKi7raPFb+6Q+YctII7GfX5dShjR
6ikQpVHO5RHNT+S/ic2AQXq5Yj0I5hHPk9Dh5ngT/e2NXcta2v/4YqyyjcaRukD/
+Y7TzDAGec/5UiOyohZwT8Kqcdxvbr68SqK8RsTadxnAFiV7UyCwNCo0Lp6L5O3G
i7AJyIQUJ3u+OwYoJshXmbCK7kU1lGVlGxLcPLxP9VQAu1qnlGuJ/ZhVwCkMjO1V
TDph2FLoGJfKVUAdcTz/XwV9aileK1NoxxnRX+Yw7tqLVHUgcH69HtV6xr447ouy
jDAtif8tqhba+heMT4xZ+l7/QtTFK+FAnzuaPOV/Tr1qNRiCeG1NV1mUuuIPFtt2
lCGrPdhrfw15j938kDKncQm2s82FKOm5HcO0sjTBeP5NMezy5aPTlYViNfeCIqVz
RfZDiagBzoktfrgETDNncxeHPyAPGsVBZ1U4OYgo0z1Nm2L4tOOXi/bAEqOXocIw
byZW8hyotZiI0BrNoLHFvNKJZlSX0fW0fhgxy2z/O+dsy1MMS9rrw1stCIQM/Pvx
MAUCEiWdb14dNG4hxy1r2hgM5z0+UWPdmeL0SFm0dz7msQzeYk3mfgZW7wcJxGQf
feul4WMKMOelQQW/4kOSvPlRlRV+h37qAZXcS6W84LAIBOqhM6JFPIONEHlFza0p
ilDG5+QprHnRL2NJrQ2OO5JkwWNub4bWejrxGMZ9Z0c0iSmbpI+4yxzYb9TIl0Ls
lXdzf138eRVxWT2cvTgnN/eAuN33YdcTd1Nk7K7h2IUZ5iJ+5gHVWnfYa2QPmgif
Ea/ZdCSZx+14PsVj6SZ52YzIU2734iAdpHKeDQL0QjO6KSDDqJeQxg3irfT1VXDu
R2iU38X7hkNi9DYgwjRmLZdQrT4iu2J3ZXI4W7DsuvN53m3cAMnGN+XChTxw7Y71
N3XX0Kkgohl9xrt07YRbReU/uVwtWVb28YVxdJIFoMF4NgkrASmMaHRTqaJ7C6br
QmP97m3+1/Rf3+yRAqvGJNhSGiieEza5SJ0uGem69/5+W3VyhykdnV5y2HoJlnMm
iitLhDRcR9zj7kNPOs55rM3Y4+X1RiB2ndA4tnTbB1YXdWEYSLZIiN2E+uEWiunl
8l4T0Xze5OjanijnayVlEbutyZpATrNyaoIvNDSHFIgdHZeE1qSQrxGq3KV3cOn+
8NfCAXxZQGD+xxdFEm+xziSwK+fAPdhomdYFEBsmH8pcXVhWRwNAOuvKjX0I/I78
nVrwMqGkLK9nrwpYaTA5MZx+B+64/w+3aZWc+3EYlb7ljeG+A8YHlfIVCQrQqf7m
imuCXNSAVmdyBGuzIp0K9pmzw+lIfEJifUyVv8XI20cqvGNDDMBbb30C0EQWrubc
OzZLjddoxoxXhC0ITqvVky/t0Bhs3x/NrX74aHp21DlbLMTOGWerj5CCegF+emNK
jilpcwhD2t7rF1SJmgf1B3PozjOIhcmQNHUKU12jZ7rdANv0D/3tRQ8HdP3Jr0A4
9BZrohvCzgt/5dYMcvTHpaUCfOGYXZ7Fm6lzBK7mZAwGLoZZjCtqY/Jc8ruuNfqV
qav+k+hi1LloaBckGo9EqHHA75/bo5U0mxosuJleC48p9xeQDSE0lCSPz3+YSAtd
JgA3Ziv+StUTv6QHUQX6AFFSGqIvNzlAja/k/HoxNCGuUMBMXtYRw1W7rneiTeEJ
pg90uXEFRG7Yev3G1uilIbLxekZxMs2Kioe2pyw93US+EDSOPmi5WQupuOunL5Qi
wrZ7Hnjp2WxssNVspFhWeA2tcvLsJwwlR4cMRE1YflC5ZR9wm3UKAPhNaD942ZlU
5pfqxgGR3mK/x097PqfGJs/VhDV7/TPd55+VEGAM7qTIWzF3qBsBhLzeiCIIsMHK
8/ptgUgVTcoyZiQ8k/02YIMh4NiK5P1fvnlfM+ZzeIzvp5KiFQ0GHtkV+wr9L82O
KI2YWZeU3tM76Liu9SrISGMUDiLiRsXV7mPGXzUwfNZnt2khMF9kqMk4DRf3mfJq
FUPqR7CiHZ467HyG756ObzH9i2NdapmTNpvk67LFHy6pjHyLdvEsrAijW5ePCX+D
WfSAHh5HDfISCzmwEYP4/RQx+WkkS/JC5VlqXQk156pRgWGUMd0f3td7ORgh/A9R
G5ZTkcxodmfrOwR8C1oj31t3fTgRWobao9dRkoYzsF2/n3hEbs+yPCOFe/sPJPFY
9enqNNsJW98cWY2bVocOZr4k2IF8YmSYPQlSezYJvl3rTCfB/+KXZmMBwB6xrwk6
GPqikXUcL1zCIUm3spL+b5T00Rgr/jcWfOAdESXcDmEBo86kWgfFEB3B18ACssUo
yoZJ+RJfxGEsBiqQLpVcbU5dPTxq2LZGfNPqWzRPFu+2pwy3Nl73v7Z9GDaEH6XI
r/f32px4mEPfUxt4RMRI+jelvwZCfvH4ODrwWaBj/G61dJA6L6ipz6nq9CdA2PTy
U7JFTSvdj67AXl7ih2rEWWTJTEnUqz1O2WfGeUnXlsKDTVAcgbvLLsolfdr+Ojy5
0/tk3fFGjMcOCH1/+AXBT+AHA65rtl6uioNt0HTLPPIOtvvyUtbb5Whq1nx89vLC
TgHMtwDWg1VxgHAVAFsfomb2YUNMqyzB8nLPjlS3Xmd8jXmw85HpPkQFOuXZxmKE
q1Ek4DcsbTdxnd59JUCeXBP51sWO6rpGnVyCKtHno7x2jawP7uQQFyGRaR3l+dqm
bZLndzg4VUZjflVOZLiUzVHh6CP3PweSQhrm6t6QkNxVwZMBTxPKSzoP5DQKKkg2
eYm7hDowgAVnFm8ThSgS6e4tV/SLc28x7+B3VOwPXhhYMTnusJZk493SufdjT11S
I0IhtRnAVJ70hxO5j1Zar6QVCmW2n0sGS16yNVyJiUbxgQ6hKeyxgU1+ui7HTXLh
v3SnOiaKtQ883KARqcRiyN4+n9I8tMACde30MSHDkh3dwluj3aY+yoQlyBtLrqDG
2BRWGKQHpkDqxViCDefDmHFrSqFx0yOHI5Vsu57Pj7VF8AEUbgdM+JHTC42rq1X0
AL3DlYbEOeWx++tOtDtDUoD5ddBdSIo763eep3NubqMNo+hkRIHcfuG+tQMplZxC
FqYEHgPDmF2FHToa4ByBdUc6Wh9mVGTHRzdxTZku6WFElxX2WGspFo0jMD+UPibn
fQPnmxgw52biRVlxvOOAlhN447ruZn8EOQN85PSP0Au8omtGYS2Z9AhoMwgjgbWb
XSU0tFUokAjavQ++gYmKItXXvkVFEqoYhWBS09Lf3dxkQjbCkVITiGxerejnkV9H
mtVr4iGTHkgMVkv4job62s3UtiPnvUa8NpEUyMnt18pPUPMcuPiPC48sOGxlzmzJ
Lkl8ouDuf8/+jM962+UPcIIo64o/0gHSYExQBunXPbziNgux/Koh02jWMxtCiZ/m
n852dJ/cbp1luAZ6JPgav2gau9NkCEtDjZezFCM8ByqntGSwf9umyMeIWAUfG/QD
UgBLsC/VkFHlcBCDG25t6EXIhb0KbmkxXaXsWYjmcQAlqcrJHZX398P7d2wRZMsV
/pgo3XRKCiqRsNj3/cYm1/vyZS5T8Vi5T3A+cMGaAZkRb7v4Z5evwsZV6haNH+Vp
EBzWZmewI/VPM+rrzq7BjzxM6UPhFWO0JNzZPeGdDwZGA6ArbdbG0E5b3JutK1pm
RZM7qw+QarSBfmS6qfCILhXV4D/ppXWvPxN4ULZuKYbB4gqejfnWwXEnWPwYbl+u
S9JA4Dxq5J6JoJmJvDfLe416FjCL8b0+kDe080/3WHbz+CMdlFFNNi74YSCQ2Nid
iOckhgP2AP9vG4heIc+VRLzJXI0uKDpShU0zdOXY4nitGCrC3UKdqNJCN33Z6cj4
30jaxd1V8g0a1VBQoA2DEld4NRzQdwzQdkUXu6cLSxWleffiIsCGv+W6yXqcBeWV
cHwQiTS4rNJfHuEUdurIiP5oCxd1ImJufT0HeHOehjBXajg7+Xk1bKHTZWgSNOIf
cPeypOdzmVtA69oI0IkpocCOpXN23Qf8RiQViqxmAGTy/JBZx7mSKYNz+tQUWhh2
FsiSB/fxINDKg4YWer51SE9z9drVReWHNq8s37C7dPjroCu9t6XBl4RINqlg84z/
6LakR1XB5/+UV5QXOkuCsXxQTh1lm3CS2/ECge4EunBFT5ed2c7431BKua02iphy
OWVI5ebUuSXkXSCG1XSTOG7ByCkzWw9nqfhDpocFlglhN5nFxPGqakjjq3zBimzU
RGbNBm8XTm08svBaWDFMC7FjKXuelZ435qLEMBJBpOEUgJYOo5L1iRE7da3697UZ
x4flOV3Rq50aAFBEBVHzF13srL3DoazWHKJlBpqS1ke8TpoT8YQoI+n+E35eapQL
Znhp8DK71YQkLhSaO/0kaayLaUZ3nf3kCpzZO89cg8WxPHPG1QkEGeH5+XrCmc7l
QRagfsAJfE0v+sOvfT3YPb1mPxnHnOLkfQjBmtJseko65dSMtYVqBFupPIjvHnyJ
U0WQzVDX0fCO1Rv7pLNCiZMLVwBWXIBnuwKde8U+ZkCWwd8sKXHuYX8jcwu44c9y
zS8lma8UmAP6ZumQTfV1p6kgINWdR5ztsU45ZqJ+5yYavsbscFmcxFasNJ8jkeXC
brNWJFvA52VUgjHJHb+uQbagdi4MF+amhslEIFZnvSZQAbTfhJbHNqK3PimwNLiW
K9Ttv2YXL1gCNjCzDLyiVSPWhsfZkeTaI2X6O8cmTKepKzAeTZGQBiv9aN4HIQN0
68nS74J1QiVL5aqG8OABS9IObKRmzeKaa8IK6rNZF5AY/TPpPtIkWE2NavpSkIXn
MtTOsfdCCGIsgYj2U9oSaZXmRV/a/1tM6U2LY1j4PTQYtqSKZLPvwjKHUWU6xgc6
5oLHEqR1pwxJW2VdJ0f1dIIBKoGx1YPapQDJW88fiJR4i54n2T0m0MrFb5kSybdd
8ykS1yeZRVTQSZ83zhUsqGrCykyz+HS0O/BIwQHLgmouPFlyspCe/oJI99JyTfUH
4WCVe4QCbSJEIX2ECfX2ALW85UwR7hrI+Hj8ouoEs4odvGwcZtlyIOceNLeco5mV
EjVW7jmFpCjOs526lFEsM7mBFX+e094OcnQm1vHBbLf16WJWar29vqtTp3NB9hIu
amtn8p+HY++nY0lfEnT7FVOzdcExL00Gd98WtjpHHgbOZq7qDBYTPc15uJsmrwj2
QavAlF1EaGDitTLKA5gSHdRaiIpiXNBcKXvz8Mbg+RyrMHH3PhPcxQ9Cuiol5/TH
RpZmOhj0XzOXB4ZZvvPPExcjNhlRKFDx0KA/eIefq13xy+Kui5r1gWa1+QWrXSoh
Ibh794dvlPXSnpi31yHQ0wsqp+WY4t/zEwSeUoGqVegml5DTkb01eGNLwVQW+yLY
4sOX215PoDcAGwE0bdps8SbexUWcfwIH1p4XJ58ldU2Iwkc+LPqjj2Fd8HbJf61D
6FL7K6D10LLJZyyYvZ9tUHCbOMow4pg13eSUg1iJnkDQFbZvIdjsly5sMem8LPXT
EfipLiDpeMd21ZB6TeV7grG+sOOjGiIFQ2IAB1dEXAQg10orVXw1xLGjPztcvvA1
oUA5fxIZ2RMT9oU0fbIawBHDjwNqIzmmHkGlI/Utxg1oJPwslgvhtuGRTs9alErW
x9HDVD6puxDG0TPQWtRtXkQ+r+/Wh+6ucqdg5o9jQDY6waA7m+OsudoI1yy9831F
9ekMQYaw81QSFZooPaMG4sR/UySjzIYUSqOaSiWno3EKeS1EgkmydCGQ8Pa650LE
KKnvpGrQfnYuToshaNayug6vzCRMiaopGMK28VYA9+wDhoqUvRhG5yALMY/mQyE+
ULWFf9nsJ6FVOqQ6sMFG4/4qXliHoOMAHklGEqvjzMaO4MgufoAwxcdYuFp9Pq5A
ta/I2ZqcaSNJDzZelrvJzZtJILJTPN9NYDyHE5ADYq7NNu0kV0FPBlIfnG/uQB15
zQswu8I1zXxDZ5XJYQh3j3rb8unue8u3gZ946G2SGpx8FNzZn26RY3aJTUJdoT3o
31HRlATtMpzWlb6XdFqqt0R1oT/wRczTf7IC5D6ZRfqmW3kG5mUYyUMViY++q1rg
6SRr7ZPul9fit4UWrWePje+skM3a6U1Ru4zkrn3rMUS62SLuzKY+9rL3tFW5c8R+
zk6zWV/jI63FavQYc7nKLp+rFlML2VshBWVHFTiXKXma0RSLS7eC63SAO9uypBLK
GoAFp2X+EXdoyT01Ju/XP+fyCj8m+4YdZtnEiRAOrpY+I2CZdmQGcwaiiLueKHmt
6rcH+F8WOMTbE3pADHGp2ld+y6bL3C4S0nVtNNM0NzGzZaLTwB6MFcLMW5CF8PNp
pInoJvc44NXzrGs2TfwcmzsirB+325Px5B8RE1yzXtFT07YeoDfJ/BO/qUbk3wQW
CCiah/q2uuHX4uRaeaGiTR0i1Y+cJTU2jsXiNydfopyAciK1Uo4rVFv9odKHex1K
aSzl6uPYhUrpKG25g8j83LemXbRnJlGaC4zsUBO1mFpdpwSbjgifbH8LAcmAAsHq
pz4W2UGqUKIjPYj4hBuYB2bTao9EVGkeS0LbWseaWO1U7VIuXGRhR/78If20tBGE
vmwlxF4xCeONipwAocFLgNwRbVOcV7jEkklZjfliaek93EuM7RmMy3qrdiSbB5GO
pYeihBu2v7RIrfdl79Lyaghb4Ix1mz7oDdwTxoV7vWzbp4zMlRRHAKW9RGPP2Uec
Ys+Zu4Cu05H+T/RS7KdGLar6eyk5kyFtn1D5RCkcNNEOJ5Sm0nl+E3CYFZwe6MAJ
taqK2SbfFff+9rv7JLx/LZY4IXRR4rV+umk6BkyC1JrjxkX007sukQz7Cu7aAy/B
IPvkdfw1PPUkb23r8uurjB30ZwSmHQ3Kb739AoxT01LQK7TbKnzjw1Svw4ifd6yw
OiCbkQGQplW2B5AiwkLrMPn1KO3C9MHKDZeNO4U3lOMS1+5gnXRuk9LU90cOdR/W
gER4nmkPuv75pzlhC8ZXtIgtrTrBRWH3hkxsTV+R6cdx9eIVPsQ8XGfb6gAJNw7m
LBozEs6XXCd8c0ILgVMcIWRatvg7Er0GH045AOe3mnnI/dm/4K2zptEPg+KNsRV9
wzNbSTwMa9/v4fgRU0mAI4XJg++fPE3+GDGMv9PEwh7fKsoeCyt4qU0D7KtonpYE
Z7jAAfKxn2ewslhMh1TRnW4cOULNlRWYw5zWiI0X73PvzIA6wK2flWhQJnX4Vmod
EJ2wUjBBYDtwddWd58f4q3C0dZV7mCbd8umRg9f25QOo3CxggEZhJn5b015UOPe+
Md9DlaXn080M/ItWeQwp+62zUnunklDZ++eijIYmJERsH3W6wky1VNE8xv58h0Zu
JDGZXCMuVMTOShS6bNxRL8HFBmsTdi2No8QNcoiwEFYNzkyhVBbOB9DFYDdtrpM+
KvvrcUfrPoC4Te12A1+BFf3sb1BURXn2BBL8u60jQbPUg6yxTd/KWzLdyqY3lw9Z
nsZULoQc5tM+n+Kyw8ouvG4IaN/CQld7r+iuXw9fRo9AOiaAQw9D3p3Sija9++91
IAYMmHUxf+3vxlX+P80MrxD5zFQ40YTlOQFC9NIcYeyaVBBhNIqsRESXc7NQQZUX
2eudEz9rDoTcbU/XnPg1O5wfsIx/7K5jUBN10Ppi7UETEvrZsbVehroBq9vco+K6
c3LHKuZgvqSdiSm1x4bMCCTPp9K/pK0pdEkfyebIPIZX0fAwUJvA2Dmua7irPFmR
EgNS4FUqp7Xb3QdKAF3KdrSCUfEcdZ7CHPrvKYx09bZKt8GyLZaP+kw9+foDXU9D
BTdWbEE1QfESOEQ0CkVY8V9nYD4xp4fg64OH57vxn3cLxALPvm6IIiCfltZol0QR
BMNUIxvg23HJn6QdLbPXafDfr+3keQqM7DNpDdY07WWG/WpZMPcnssg8wyCt6+S3
jO+ttTDlTWWSsRlALJpxYFur+Oz9ieIAW28QRntaeaHTXBEQ7Z9ET/QRfw0YWq6E
BJSlrsRZwmDFlbVhUvP5LgTTrPBrqHcyWZS8/7n7DinWAyVUbpTFd5Sq3vW5Cc/K
4KRl1QKSM4JiIeGb/D64p6/oOrHO/aiMBjWInb4diRlwkG9Dr80drwzhy1Na2e+Z
DcI3UCL6+DLHT4b8KRWYPG8ooqrdpa6TGl9P+OPf3PadGU7aq8RAfoJm7QjxNcEq
NZGjsp0g76Eb0IAbiFccFA/znU4N8GiO6l67SNNGgaK+xKmiWOTnerqtUQRNMCNq
GcfgKt/dbbFkEZG2O/3tRbr0NlwOsW0oQa7Vs0sh7dDbBDDPVXFmaKUeKpIa9LUw
XzDDYtvtKqjR5zKOOr73JG6SU4rZdzeTbLYzj1L1wgySESgMou/u++4Rcu2pYulR
zjQ01g6gaXWOPSqRBSyiX0Ij0M+C3Ai6E0irkYax7CMvwyPb8CyLL+71n+wIwOC+
rMIZOGZNJXKPyXtRZuo84sM6L+DEh9S1EPArIFG85XiQvkx7auUmr9r5aQ7PApvi
t5GHk/nezlyqg4VU9ES2CQeyKQszrV7VOEbtlU0OqSuEdgCM0P4/mHyoKq3iL6uL
YlIwNv9ePFL2E8vtFDonc9ruPfSMFcaanjhunkQu0bjBtvmURkdBCPtxCh7hgsRf
dqyAm+Jku3uk6r+4aZOL3ve/3cux2Ri/OZkm8Ye0McrwMW3svdCj3LAZQRDoarEd
A7giLVyOkGQ/+U/8jVu1MvNvxkzFTtk1rCczYXT2V+jhMxGvSzfO3wRYX/Mgdhd2
7Gz4icux3uP2+Qc6+lymyDv3eht7OqUbFF3gPVDYVojqwXamX+U/5P2erp0MQ9p9
z9eGWxyBUNzW4WiG0msXRX09PkLVIypgXjGvKwCtVl8IhngYL8nZM1Xq3OCqf46+
l9JYFSpw1IsOpWHK9b835hitihKxRhA1JDqZiCnuwG1QiJTwX9iqMZ8jIj00Vcbh
eANfGIC7j26mTGIsqcSmJagNQHTsAU76BXfuo6eVW0xR/YkqBkUSmNFbot8Okibh
+KsWqPbDhBHyo/BbOEejPOZkX6IZzRelEmbvokLozr+iPnJk+SGRaMhwGMos0d+Z
dbXU0o0UXxPhuV14wevuuqxcocEdrPctU6+bdv5JwgS5kqVjBWFlufcHvKthP/Xc
cLAn6VnBCeIlURq3nORHoKwXQMdrAATFqWZZ401J3pLKZF5mGgm+JsbsFNrlx7iW
jULu/xAZ8VspyTpC5FE8VLTFefx40zqR/C4WtPGiTjXphNDxVEE5dSFP9IakkFMO
qT2xb/EuyaPm5nQmn0hsbtKmeG8/tT0b2a62CrON3MqtJccmIhYU0j3Ik/kgwIv9
joWgJiLfzPsNI1O3o2tw7aUk4bBgyjT5WsrS/1Zh6EiEEv5DHoKQdKhoRedZEIAq
vF/IWlEIi6SExPLYPUzuLusTeqbjBYDRCWqiwHUtwqcTGkwDokU8W3W+l+P+jqs3
jvukhExuyWqlb0aj4WKey/+4+uKd0vWBliZasmPuqOP0BV2QdjEzriEQ9lADqOYA
I9VXrE+2eI7DiO4Z8Y0il3vL6N6vMV0xveE+36pmqVojb7CMwfFUcxAjaGej3IeC
g1I1O0VjUKEBnPUkminKaDvbRZFTKxRmnsRX3vP7x2O2idPL3M0dICBJOWZxeh3e
ZZchakL/7csUv+dyECROo/46rQQxuLaVW3jEzI719lGuQ6RuX0WitiSApOd7zVb8
110wzYU81VNuDrMMXgbnupNWwj0wzPVWYKwt5mcbyMtBVq4dztv9xUbLHocZYkal
hxguu76I8PHbLhxc4vnspA5fy0QcjfBPo8xIgmC8bLCujumOVCFTLU0vo8uAicEc
vNC0L+GuYf3iEWsrQ+7BMG+fiwkD/HM8GJNuW9nuaKRlaBYK087r07FsmxgIdSiB
PuTpFP+pzJVMdO/pGlYEG7BZEgVx0S46s+GecswOGPk68KiqWhVCSqwngfkgI28H
rtgDjiSOtK0COCYbpd8HrZpcwhHZS2IVAWDbEUqdr4DHFMTTEEUtCilnEt1T+0M7
gPvZnPxCxprkq2v/6xatQBPc+xbwLftRFD1mi1p0hewUKVwT4VTupxV2BHO0zGYE
aORctyIHh7t0Zlbq3Srlqd3/Ny+hDUybeqS8ZyCKNDFATlGoukCOAnEnLWrPEExS
2yDOzQ5gwRPIAZv9knBHWI+bTpalxs0AadItyCvz6Nl3S7mDvpM/cEtCEZZJpPLf
ENVxpZVZZbrbkKjqAmwnkHDaTCYkEryXNEnnOZvw7f1cklm546OrttcRxAvEtBqg
1eyAFoX2ICsnL98hWfIwx/p7Wc4Cr48KSuncKYxjRZVLMj5GDZcMwOKSdsbQ03Wr
D58IxImpyP+aEq39bdir/RnGjjVD/a7LRud+m+IfsOU8encZPnmCizyROazrfBNW
QIAf7Iyz3PGN7Imf+8BvK9qDpL4S1nKvLVvKHqBd0wAyxtHyj8QtCrsg637/bb4x
XkIJho7p0+AjmUgeDV3ATjjGQ9xGWpUojHiroIXKLEtwByuWaCBLtyfGl4rIwfqe
BMLGbdKi4J1Z6nSjHfr10w8cjrGvmpYoVeIrQoucessGOSZhAxaf/MeStZUiIsZx
xhv9YQIx8kqKEA4XZhGQrOGlkx9NEr2OGCJfjWvcZ4l/xq5rr3GZwlnbrJGOunBF
zMn5USazMcth6bnjIcDCcN0sRA4yT2OyNbvs5RkntWihSA5kZilDfQejGCNIwi7P
sCWP/eTMMyVu0YmZzkcr/0Ohgfg+HCVBWWwXemgZoM0cLjarQYFdl18s74Vlwke5
ZFMD5mtaMdlZbXxJ3e5+d0sjNKz0k5NnMN5R6jf6IQOefkXSNlQ6A/EJ5LpzpIpt
rAhU9bsISIbHUMU7VNXuzzwj/BRGCL+EFK4NlNbyK3gM/l4PUNC1qnE+PlZTX9NJ
9BSbg5qERkIKR41ky+MbEmPQretcTy4tSBoY5Tqc/eNnpb5CUtW4a6tXicouGwOj
tWSKGXjjoRLZZIySO3d6+lAaDWcOZhsh8RQPIKKb2fgrz9GwZqmBtzFjFu5wIgUB
nPH9CWjHSoKAK4qUeD03ZxdSvYh6eTxn17aNlHQVPbBN5QpWxLdgrq5di5eGXqiN
jwpq3YIxQErEgpN14PLPAm2vIWA6LuNjQxj4PPaMEhuP4XLA4HQcGIKrx9SirUYb
YfxHH9q6emmN0nqoIyg7yYL3P9kRw04hqPJIlpBk2qbAkdELdVMe0mPYwOLawr4d
+gsLG/vovTXNwtj0RS8Hq0E6KLiL3dPEUmgM1S+NmvefHVSH5bpwOGSht/f1Twd1
/R+wILCjZIGSRGPOiUqWQP9fEVDD/3SzI43slj7jR4ntCrpZHxCTaa1h8z03TXRJ
6FlZB8znWHBv/3NJzXvmEn4lK5xsqifIz+teH+c4KJn/IWRVzMzcCXUXRMI1wYYy
lFU+BO2g+PWvfBBUme7CxwtX/0WZDfxsChOLc51aFkuFUC/akqlqjL8FPwu3JD/l
9a/anAnMTc5MJ5Vyxuc5uo7xQ95Fb7JLZpO8SGi+qB81Ct1qx62oHGd5iiH8GU9T
qoyy+tDTBwGlQkBW+cUDO+YM2ALIZYuOE4MpNxauQfl+nu5CmKNHykbZA7DI4Xls
YJDssvJ+747SJRB/LeXQJU0Z1dnqnua8JpnMc3SAU7N0Wv+VJ04kdd2AMLiUyz+D
jWRlgsyaWS4qmBqbGDomqnwq/VIDFtCQ3bZlFq13+IPKEOL0Z77c+QnQajqOTV/W
Grqk/7Ghw+0YvQl9hlMiCBU4YzPLfk3nkfgUHpKIByMLiYCbjj8w5WfXS6KvKeOm
XgrPlqKYeHZX65PxIasDsxmzeJkCxJpey8eKaZv0Hwd6DeO8fVuKDM7xZ7cKG7bc
KKbIf54NoGCvosOQA2/6X4OpTvDgM3vcq2o3/HMyov7pXBnbfRwGoxX1srPQY6Ur
t14wPAHHnANlSTHtntoe6Pkt4nJhmNUgEUxjUlpkgpP7IHvEjqaS507YpXve8SML
oV155IZyE/ioi6YVf/qmZ1ZEwGrznYeLt6XkgCVV4iXglpZ/0Jyyx/QEfMKtpwx/
0S7lHHsDFptDDxVQTUupeRhACTjiYb3gBjyYy4zIJzmQV57N+qB2b671HVpdyvro
AeARd0XuR3708tuKxziHitIGB35u/ui1316xt26Zp7LMs45/elqOgQ34nj0Dmz/p
hpTfhDsS0Kp6YdxE6WNi+/VqB9A6w8YgdDdAEs3GZHrxTuLYn2EfxIcpjzD/pg9P
Xa7CJUZCsCaba+PMETRHrCFb0JTrpgIrLgQMy/DIVMGJjVnnx3qMvfizg2fknPvj
7jNEOIM2+LdNhuKXratOx6deOQtTSKU423fgrQk4Nlxywm8CLiMaEJcX9Sfs9NXp
CtIMwHLUAGaJJ/uKg3HVbWNko7yK9O3xquVfAvdpnXTD3Qf9J/zHV4LKnzHBp4fY
i8wgsknJi0X8GZaf5Ecdt6CSyi4qVAN/cl6319Ca88eCu2E0TzxEyY1HU06QB0Ob
zRAynx5EP2+K9qQ8Szw5CRZ+4F4gEa11oNFaJ4Pt21ZZKpEj/afMlmSl4g8K5jdg
e2k4gYtIGv/WT2L7WBqe9+1utGZys5c+TwC8UclXfNI3tolHQbVslHP5nM27fcIG
wn0UGlslyu62ELUqY6lg1qhkDIx0+hD7GfrL1ShfDJSjNIiFiYQyhZqeGa0i8gTp
M8JPykHPA6frZUE8RI+yjv0fk9t9vNpBsTeLrw+wjRV316w4PXtSPM7vBiri6s1I
VabtKQUhddWJqJyjWG4Nx4lnBfiJenu7e1Myuattasx3VdnoakyPmEeDLAATR9fC
QB6+MuJQ5OACvpy6JIh1jhFQVDltdI9r3ljTlUQCr8PvxtamSxBFy2ZqeEApV/J+
ZwvFuUoxoiEYeKJBvqlF3M/3TLnQUzmrEGqLW+yE4Dce/ObxEhGDyQ4boCzS+XgI
CRCOCLlp4eToEw6cf3TiIPwZRd3NWU1QH0LwlggIfYYw0rNraELdDj8ajLo3wDYk
US9kiZSnuBJaKLjGv+0eYIpgkMdt9BqCtSHc/Gj0CvavQib9sqlIBso57FfbhDz6
+KG0gwgB6vXLmiQGuD1/XXtI5b/IcF7dwshPyNawtqdb4VCW1IhaF7mkFFiUwMZF
gEMcSespQ/JEVW6hjMx8NNwwBidhuusJMObHimisx0/rlbMdrFV4gNpO7c2GDERp
fNIgiDiy3L7D6+w74sBktehx2NLBOTHZCyPZRw2aevGFz0N9fuVwusb6N3+xnLQT
/8AQR7sd2rIbQvue3ZEW/5RB4q2bwOM4+BxvKDtQwTSRAAAyuqLwZNYU4jKlWUoM
tnRCYWKZgjZQQGph994hMZvJjZ1/laQaBSfspzRG0j/YdZX0n60GYGMH1EZJ5Sn3
urS0vl0Cd9+Aj5VSH8vi//gUftzxVXsLsPbk38MCbCZhLBPPu6IVOzOhFUAEak/b
nDgaTg95HOHTWrQgkIENPqM7VYKq3ZENmDXuFiRPhMKX+QMoak4R7oyALSg/Ymt1
sA0mCye3XmwrlvROUinGV6N8Zkl9vVMMQEssGIiDVr3wwfaEiZiNZh1V0NyhUvrT
TBwQLgQnh+0g+X9h9Y+FiaYvGQlgyZGaBakozRT/PFjxxRwoQph9QEsGxF9enxCX
XnjHmFl4nvAmU2NJBYFPlJ+ygUGWkXWl+waT1j9eymAKAsjqPjk98yUozlP5sibv
gzQE00TM/IqUYjuEg3DOeD88i0VMzitKrPawoQPvV0gdoACp2usbTmNg8MnevBIV
2eoL3Mvs5QPpokIaErNeQqngRPazkNWD+MOrkH9tnfBGlGxKMUhSKuN1aPU8Cj1c
4wFzD0zeN/HHSOea/JPAmq95O6/JyTbre1frhVP10RKrKYxOgd23Q6gGW4kuE9V+
OzPgKUghWeCk036gLi2f/bPB0TbdMxpoVVr7WVqYbHPGum7F54ZCTlBTaZaKPvH2
CRqfwyvuPDZUsa1TFXSb0hbawMdPcMq+AR+JNdLPsv45FDVkkl2c1brxBLXY+qFx
KnTpu3Ql5+fIPISRmpvV2OnVWQghyFzCdOg6h2j/bSeGdCIxO5GJcb+NGm5kmyGb
f5ONxNnf/wLpN9nJ2w48EAoaEaUlmuhG0eqiMNt8S5x9I2P/F2u1kOMMdo8bhPL/
aZbnA7zQKPkvfULuttqg/u2mQ7shGLaur2nK02fMwrHEqN439Nl+ROTaHmy/i9Yi
0MghPGiMgBP5noll69aAyp/VYpKQDk61dEleoU9ML9NNqCLo7OxuvLpiCrmDcmAg
00cvQjtHsAGiMEmYv1nin89IKemfNUrE/O3pYIYhPSJKNiGl6G/aKiMPrncARpr7
7dgqeblU70SdSpkQlUIzYNQlM97oXD8JmcyTwNte34FDy7mLXh0PPU41NHvm2goh
rUJVazrjnaxs0OtpiFq9mmkKN6hzc0rBO9l+1KCCSigl5o1ADogJxQ1/CdHtWyfa
Y68jOdZ5ijFY7BxV39hVQ/KAOi0/DzcUNBycUNw8fM5ZneVPHSKXbsKgVm7QOTc8
5wPA+OKKYZ7aWfs/aJoGd+T5vjFq7aoIlzNRQHIuYHFvgYYD2IkE54FiXkbPs+Oc
naQEDcYeYsxgjQrt5Tbp5/PpNMIvO4OKyCN7XwTsPiknUWoVrFrcLfRrdEi5HCwU
nO1jmF0gbpLloZcWgR72SPUkxXCY0jU8/kGYTWuvju80J6ITAxTIUH+h7xa3n9W8
2vD1qDbRJWVk6ZB4FvJbkIjRRNVMPohcksgzOFtiGLfmu64VAWtTJ2cIVfus0aED
7+qqfZzsghS92u85v8pDaQXg0YSXGngQNtontdyHOCMRGGCKPaVCxCvsyjQPDbCO
wOUdslQSDCsWBNvjeeYAx5Mx6zMgbLjkd8tH1kJvw3UpdASevQUnT2wqDWfN2NXz
MIHrhI0Q34FcJzzJXw+4VHKebC6t1g9fWFQIupil1El0pWKayG6hAs6cqiGQeBpf
isR6WGdYKvXIUC88oULCM2hvUEzhlp8MAVsVUMNQtXfaauudhc1OxBPN3LNhV62b
akmEu5k1WRpMMZBmLCsxWA/vkOCEmJV05skbGH8ydnXM+ykziACkPfUCgXm4+ikX
LippFUyfVdndf0GXMVmOdOZ177lZFxyx99/nUf2CskLpfYTHlFY5/5ZFXJX2mhBL
VifDhEnnX9umZPWlgZ7+7u4PWLEQbiXgEYnLK1kyAky/lbgIhuX7iOGDket+1d5r
UN6WkzEeW0Nfgv2IOkANbRqa437ziJh6b2xoxfbrjEoPp33miSicX0JMelMN1zSu
HF5SuSHFS1z2v74SQQOj9i3hT38p9QiHy2/jq6+QE78K5bhFOgSsxYjR1X+MYUJE
GdNUgi5z/L/BTHk8KT+9nfpq7ApzyO4PF5vSq9XhEe+3ob9At++zvBUbx/cb2IDu
MoQQxBJZIGJh9ME7HPZAaAYYKVyOz/myHzGvV80PY6ZnQ77xo9SHL84ES1OPxyJ8
/M6wPSS6OprjhzVK0otn3lkjCbjEC/0mH98RyEl1Eyf4f6bS9q7XTd6vD2R5FPDx
c5OXvvEw20PgeBqvumx3tkGXxXMMGPFSXbCBEu2KlZZ6j1liOI8l/jmKm5VnAT3+
soaeZ/6PSJACIZa1L5JwZ2yk8AmINv0mZu+v80k4VBm0lthY5rqL6F1kTHdA3lOB
AIU3CRxgP9q2P2KMPlX9ldg0Y2C4WjvvSGfCvawZgz/4Bp0IRcPvCwXoOSXZE8rL
ptklUXgslMjgsnMta/BtnxAbJgnsCehnl+Zjle1lT0GJLhbRMqSl7ICd3X1c1pIP
T5PXYnwr1jZb+OUYOmfiwns6EeFP7gWw1Q7faaSV1DrqBLTOkRpZ+0ZRkvZ99TW8
FpddlU8PIZ9XkT5SE/A0mk0EmyZETJjYp/leo2TmEtgBTMuxcnIel05nsrnY1ZfD
DLx4b13TJFakXwjMBREOBajJ8Dvmmsj9JC+6ESZcHvSK/746IpXR82co2+ERqJI2
Yd/j1U/j5onl+qS7LAZJqhsHbLpIRINYGCYzwnxsDXq6lkY/pcqRVog4JO1KHmTa
XzUrfZv3FWw8n91KgByYKGQUIYprjBMov6gYIljmU/izw0nOaDqktmvW6mTN6pAr
2FdHjGpNKxo05TQbfgQOm6TxE5LlyD1We/M5U55g3okMsUUqXQMvb8BS0dS/rN1b
oBRNq9+lRq16UsQPnegngXDbbXVsc+0I12Usxyluo71CQ5s6Ju4194nfmolTpSwD
NZBIWGBkkh7qpX7S4KcEHL/d7GrOGXlMqcg+IyT8qmMGZO9kkiXmfmws94XjPjEW
wjbb9c4IlBqdXWopA4OPfxCWm6TTltgBj0iIOWNql63mG5F4viI/uclmTbn5QuYj
SxYHvez2QImIovKuzZaXLO+7bDoxAW42ygInNmBHBcujzkgOn8Mv7aaC4w9N4Eo6
yH4hMAqbsuHF3wJATo8CsBjor+r1omw4kqBrPyq8uVDMALY3riqlS/8eJaEINAj/
4tv18oxsYiEBRcS44R0m7GaZrq1SbTt/FKgo1a7l2q5Lx8G6Jkc9EyJJx7QOYlS2
DktdVb8Q3A+0cINr6qhMhisGuYo/T3kEhu8026UfYgXzCeC/Cc5egkm+kFXtAoAI
wu3okKlatvtbd3nfrWclb3crWok5LmwoUOP66VNfMMLTLKQLdENWp7beCUAp779Z
ytr4e/ECyzhU9UNKCyA7McSZ1dIM2WMzuLTwFPAIRQMC1ZXvhE/3k0HV26M7yZWE
wTxmE+D1fhFvCek8bkLcY6c67iZsySY4yqzkeGxW7WH5GmDac9Ze98iBg4ddGiQD
diMfQBgHvDlKMfO9zvRRVOvN+odEHyodmMiZlt42IspOF1dOQ2/HITfuN4AdcZea
qFloWdLD0kDGbynYfZwf3f8fKvDivEfz3iqOvEZR7Y2b1Fa5QlMh1V0fZ/ctEmD2
cqJNE2ecadoCXEoGLibwIC7Q2JwVkByIOr9dwmtQNbgOY83GXjjFdMq0KDv7uWOc
tBXx3s1ssEVftGePeHu7lIjUHYbVc5PA8oo/t/z3lO5eTjaRxYsKibeaNuBRkjfG
2hwPy3lZrmd1UZWvoa9ML0rBoXzPU/c1mIpc4J2NUtPiaIC0mjBEjySGqjwMVuK/
Ywopo8E5oUrtDHheBhBv3MfaFsDaceZx2LzKH5DONJVbYVi1nvbuemapApnQOFxH
p2u7o6TFtLv3dVna7dZvojQRObmWnFj/fM4+LQ4XahgsKEgQnxHq2EBMaeyZyxrB
dqTYUFEYkwFv7hIaBn8N7fHNh2h3KE73fJgsuUnXpPSm65tj/02Oe3aQB8rFftcr
3EvhMzdNpdCkmTlO1tzTON1wOgh3t4vON7ykNCfuxlwrQJcS62BCeo3WxYB5N3bW
JFXC74/vj6fZNStThbLLKJaDYWfgY2TfU3Q0tGAtl6lvS/VYCgQZua0LzLSxZ4YX
a7OImTrO5i3/wQLYgGuYABHRabvDHPaSOrP0fpWqjo5soNrpRVjv+0vqvwBzenTT
+HCioH/KPb+Rj+t+buw1CPaX4nhJM3rjaokF5POMGRAtvALd2F+gBP0HB6vHkwHR
ZbeP8DDj/2B/7N5u7payuY2/l5kSE2nhH3C8Vykno9PMagvfFod2jv1ZFMbHLVWP
mrauRO19kgh9gLRCc647DMaXNXF5LBB/hFegx9wTY5DxEPkTIQb+41xSI19Joath
DboJ3LTDxMQeeztxhxLvwDcl6FLLeDXq8oW0G49Gm+lmzX5rpWdWIVZgVpQeIPV+
0l+IjaQ7sYMD0SyswNGLU29l78HrCklmN14n3UNDFc3JvBOjhOlxEDowy5jvNMTk
cFMNazQDGzWarSMA6TeoaJ21W9zSkJgyH1LwTqzphVotsVXHT8z+PRk6YGtHqs4I
mRIXRIeqYkd0h41NZoklN5G5ud9wHJsKnmFfQYRt+jgiySQboZtnAEm0utmvct0R
mm7qpZdBlEiKjRrJ8+jUJNIKFp6i2tERkF1GC189etGnhqb2mcRsdk3s+j58fjKI
Wnsd5uwC2XALhGVK9Rc4P6G2aus6db3eQUNuo/hNVJGNQLt/j0xHU9lXImsPusTm
M1/FpZyWErMziyC05cDSKrhRb+P4myJI7FerWCsF2LLKVE1aSum30R0UPe3R9sCi
7nu2mILC0Eow76RqtFaZ4nryaw+hk6VTh4950hhSl+RvSvghgqeK9EZpXvRPcbNX
hv0sQdUCYRfX1IFPKan3rf83AsVa2iH5y7y1YWwsGiR93JfwDzz0BvXCj9I3k5mT
ZTh3s2E15T9W19AxcRYM2FxG9DGmlgC3O+UN/S2l2WKiJ7RuBM81UUSpJ2zIET5F
2PtxIC/z6J5D5Hbu6KeRZbxA1VUPYBcdV0uMHP5xhlSYjkvbF5uZ6k3B7bnB+77f
2TsGB05J315qMs8dWcS8pqqLChDf2TvKAbBMtoJF8m5qj2l3rjX+SyIR8ZCJ/Mno
Yzz5DJPC/gde0pU+bAme2X42fcPO32fVnKB9pFYN/McZCOiM99Srd1x5irgMzjNu
JlNmm5izoFD0veC5gKJuCb2ALh28wcRV6dKm0SdGOLPb8WkEE9nw7BYQtaJJ+WgW
bSQhnd3IJLtYe5FXhxoeC5JU6qKS9vSz2rglxMtzaSY03Hv7JW6Ioj5zMyU2uMYW
pT8SC9N/lw3/10PN+3TDOUCXZahuI8F5pbrEvcHBe6v/1yLS+OnivpbIY7wyX7D/
wFxUVjjOTA0m9r6BgSe5jYxtkCYDQFe98sBk5xbL3FgbfbT3xg+as464Da4n4g42
zEwYxwnSlXHzwoOOu1htdAaH9GbDB37oOCWd8QbiDgOYtCiYz7e5TMTZyo1uLZv3
TXS+B7Yjl1O+hbEjwPqhRbUTX9h+7JXgOqlIYjggsvQ73dbNyZ924IEeST+GNODs
wwQfild9jePS5EW+nrIpLXWDGn70hC9uRu0LamQ6s87LsfHw9CbdU+WBLfZQHEvG
+9J46JMMtoZElg+QbX1Qh7S3I4iY9L1CO6nbr6GHjzARfw4eo+LKN1K06PMUWw/Z
KJ2YBOxVbezLKIIg329dEi6Ldq0JtmgLpnuYHaR3aj5hA+a78ktRnmBplMK9e6et
+l3SYeWVkfMEyKkwIcAkRg8nI7SE/m3mqb6x4i4iRdQOAbMqsREjig41Rr1vN9UL
dQYmE1aMSbio4OQ4v12EqUFxVRvR3TpKMIAkRyq+g2qGVKJuC72hJNeBR8NzlbjQ
Ufkgq5RzN5qiRRWC00VpxEWSffcCb8pnrhLOeVhSl+a7rlNPzAHGprdMnhtln5LI
WkIrgZbEOWjxLElo/xOZAhYCkQDUkbC4abiKwN5qg3Qlnqg7IsnxuG45KKt/LKXu
mTUj5YbS91eeDkxBta6+Io3PqifG/ban3JMwR1REO4DUaARicgTVuj1alpcRt39t
S6TWcpb6tbCGeaWFgd2qEYSN4voaysh57nwWHnD3O0MVF5K6RyHSz5WKAAGvjYr+
QOdyyOScg3qP7xoUPPIIjrvETQCaV7D1mPG5sKdSXjtN4rX6RdM4m7hDSAnS9Zsx
/9+Ts8I3NzfA56AiC8z2N61KSpVJCjUjI1fzfBkXKl5oY7TieuytJzPIjQ3FSwBn
Q1UWjFfz77/2+GcbU4MOmqKug5+qR2JKvSIeMhzPIoNiu3JjE8spWu2A/VNmCksf
sLxr34YvGO7ZSHkNWrSDcGfSuYUaPjaUxeDV5ff7xFn7KYuZxDi/zU1uHQKIrTXA
gF97T2z5YSArS5vrasgO425vHcuHn9uVZDYiqX6Smqgm3tBu2M0s8Ff18VZ0Bm7H
O4aBiZWr+9b3hXP3IxOw5d+Z9l0zyMxGeMwyLili6CCLGspHHQ4TgykCragdOIz7
6BEEE7+xe8eMePa+5JPFvpShfpN0S5xfHZCgYQMCqnxsvls8nSxuuLf7noEGY9NB
RmH2SgiMOM5FsHV0/eblARdV/oQ9Kl9ahTb5VWovVihW5Rq7Bo9BuapCsE0DtoNR
Ad/Xy5N6oUdwO9wNM6fbnFcua6FeTjgOD5ylZ90aHfJsqqHb0KcGcFQJoAz7e1uK
wOx0v4R2oTZtAZ4co5v5VryegS0yAHad8SR2p+Xd1Iey+VL9JO30ywwc+JnHmMES
IlKjpk6Bc1J2tSdaXRIyZf5DrRM8Nu/hK2iwjBqPX+LfzNnMjNWVTQsRUTl0Xycj
h6kIChN80wY4j8B/DdJmm3AVmMJtfxTm8k78VMtF26xVeOURNQnpbQDOObIqZzQb
nhWiGYbLN3/fBIDP7QEDAFfUsf2RfofQtfinj6hKeRSnQOh21HGX/Jh9iaRNHQKS
Ir82q9/jF6UdgCNcS9/kjMRcEJOi2Zp2sumOiyRg7SWZbG4h+uNGpd5GM7+ggjFa
faxIFiRglpE+VE5tEu9axQsYI+2pX0ihZz2iSYteyWjykwAY9jDxZfmO+3TTarB/
VSfLohcwqzkqMa3/4nJ/U5RLXGAybq2cr3bsyWm3NdjDgqwGbx0wfbJLGyZB1dK+
GfqrPa3mZg9CPGJon/mttS34IGKnIwrHzw5SHinMLYX60Ldp90GawMm2qaby/Cuc
bCi7w2bUXGx7OTSLH47bjFJ6M+pnc6JN6oHUX9SGebRDZIf+NwoVG7kZTrqcQZfj
vixRGTMvda/ehYvBSskjRyvXfMz8HLQqY9u0fLZxSAaxj00h2vrdmdoNPyAcNTBS
OQ/ortnDLXrV/lB5Wufwbe/ECJUynePTSJ6bQPytRADIpEv0M41753A9Gz2HBxKx
PAmPxUK79L1msi39oUCyC5AwVzmJM1lwzSuNmX8R7n+5/lSoXV1zeEhXEkpEbztq
BI9bsencXwvbRnq0Zb8Sc90bcC6UZkw5lD91vu5Y1cRZqqHg6d5YI8bSeU5B3m83
yFga6G1xe7+Rg/JgSazn3uAPDPQScQq+/M51REpZ2x8LTvJ/kbwH8BJoNmPjy5J2
EdUcitIdBuoycqm4fhO2S2ZZKEtqyM2ErJhgiU8/4og9vp2SgjApQJIxreP+dvi4
slUMvV7m17b0jxoKfTrESIOXVjTmWRIG8K6nKggVt7j9mM5vURk/mPTPWBiPfonJ
NQDwqJIm0aT3lMfz/WBETrQZxkVhi/osz2G7GkU2ZMFC5TBNrH/E5HundfHKkUOy
ym5NikIFf/uY5OmImR4bzrxgpMpvdzwUnhaHGfQ+q3v4dgcwwkiToFOf6N1SN66a
TcEFj6w1YBweSABSLAP6s7e3eqCr7CLaK00aJE/6UnXhiEy2zmkf9Aq/N2upsXbq
fLF/TXuvjdQVfoyHzk7HYt4yDujFNrnu0G12T0kq6WCRrGJw6FWRIdp8nDT32z3H
gIC/yTphaPAOLQGrTnl+iMI27sRvTHepxgTD3SSsWNMVXqthSzsCYuH0QM4B/sR2
f6I9MMoLidInXvreGlrrIVprNnzedlFyZdQb70NH6LrOz+abNauK5oOob4/Js9/m
ZrJ9EBgQIVfeQ/QqNfoaJw73Bw5zlWlAo6asBfCL61o9Ch3QnqaeebEoXhPl9MB1
5Z7ULINP7EatSKhObZWG8XRGPpM+Le2Dn84U58/+oXT74xY3OVQ45Esrs95f7qMX
eWpktOQC4On2a4yW3McQEDHM0aQfOcYGymjke/9HLJEtfYEePAj0H6u8+B0oWFuL
roUJb8U9mHMrjCIeVR3zFE3NYYQa7HOhLXl9FTiufM0H+yjJQCbNfstVsU7PMmdi
oPkwCyBUOKlWLb/8ztPCdTa83cBPwSzhiwPxXcmzRQKV4WPcIfec3qdO1MlbxfoP
wWu1c1UVCXPAg3cPE4Z6oxQsUr4yRl7iHxLMy9RKjSeg+cPo7RbOGl34kSLGF91r
jaH/CXSD3PRYVR+isMwbJSywxjcSpzYYwpCZ6Qzu45zOUVT36uErFCZfwhiXNzpR
vx/d8ONNdeQFqdqrpv6fQcY8QZEQ6x+cUkFuuq8410uEWTWcAwlcvnWmImc5G5Qx
VN4+N0Rd6z4wco02tT1HmWsiYi6yJNecN1XOXq/IKokrxd5Ufyz+GNJhydqMF4t6
oYpKzTAENPZtbnFP0aSEoI6z9ro9LTyWHZYFN1lPX3RUeEqnXZDpAyqasBPjQJh3
OWOXkA6RIYCrbH8nyFMEmJFxHh7aYqWupbABhsqXmePKZX5zC7kSDqIXnUoOX02C
N1OXqlWvHDO40LNMR2QRMiUafb1BzVP2sx7oCAAZ3KW1yheCVb6u9Xl9ndLaPeoU
11VeEhyTj5+VeoT9w1zqasLibtoTviNFZVJZkqEah6VTnnSV7pL0ywC2Gi86VJi9
/Y8JIrtdfrfVlEfdoB2VrU1qRHeMHATBng9SL2F195A0axeL+Hf64s8xAv7sCdXZ
yDb7b5XVqzALeiJQ8xrfrNbJmcMAteRGGOBhahJhy+JufZdp8bcvghUsSdqB2Lvu
i0vgKnaFUawhL6Vfm9UljBbNloI1wfd1vN7YeWtykrUUtYGInbk2EidU751C7LhS
WT8omQNQLyeZZr3PDxLf1MDAAiCK/3rzZq7mpErVKIuxFXlNsfbOQDusk0k8+V6b
wz8JMRsPO2xhJHwz1C3zInJD7imPeL3szuxxplZCQXxq0YeTL9Vaqm+slIRgQ99B
DPE2nK1hJ9oACt/0wC4+4kZFzH/UKcGuZB5PTTbGoV4O+dp1pKFuo7TkGeV8vikM
WTf0/tyeyvlAvab7bc6c2RSbRYNADzEJVgxhdzrgJPtkrjej284pCsUOWuKqxaUI
eMbTWfDv3b67HmTpyD1tFIiGCrdKajNrzcfgGJSECOhQ2Ycbakw6JB2PXYiFoXGz
SwPn3WlyoHoESjc2JZ+hkcPuwx8F/We51OHhSV7rXJwut/1yQabp0NV09OdBqzke
slqtfFaC8HKXSqGORI5Mi0W2Zrm66s4T+YcDplX58ox3enrE02V/3fO6XeU9PBLK
0CbKOcHqe3jpC2znhgAMZhlPLCGg2oS328BrvmAYcdsI2QabUx7UkXFdyurYCqxB
cmKjOBCtf5UESppmj7tSYNYQwBY8r9ObSyFjnQq3PHKv5bfSWjGAo8ZaoSD0zB97
1Uubiur5wxmiQz+9Dl+1PWXayDBK3E5TEGZW+YfIv//Bc9FFdeKpP/asOcD2DYGQ
AUv1+sERs0OaQJcO98bSzAfHYwo2BC/oU2Rud6zN74cMDBv+0OHt3ufvPZn/I5ir
uysn3IMicX221YQ2/QBnqY+nYq4TWDKFsJZvJc4ixHURAQrHBNrC1QKM+Ahl7mXj
CLSL95EkXdswmBhTGjPWkZ3lHFbjBZ32sqDLlkmTjy62Xlzb2TL2XL7LmHukDY2e
gj4+yg0IYj3O+siDj7QitS3f9wkj0+zHcQJh/SK7+5lvKhCCeVdHEv6bgeyMMUtX
bXtvQCvMASE5o2mi40VIhDyHoTahGWxVxctT7NY5T+iIj59K9BMi8PwcLgfqH/Vn
mpkqse68mB5/5QyuhTN74enE5OUi+m6tVg1kH0JGxCYc7jy7enf1zIPvyfXAA6Ky
q8XgKCUkURErwCtsuIe2g5DL9VRq0AHi8Jr/eSwaWbrwdqxkboNdKGzKVxJv6XcA
o9z1U3c+ovL5LedSbRNJd2UCFr/gwqxxfyWCUMyj5xHuWviAn7rSd58vYUG40gIP
mQWxs09MLO+kkiYqcaYe28ZAQ2B2uRPUk8vWl5c1i5fwES+dHPLCe78p7uDKGyY8
7FebzhVUSQQTbCGNlSX7Jc9UthOBUXK0hLI10Tdu06USy22FKCv/gtd2+RoWBAih
OmaEfv6LzExrVKqCGEOHzYRboh7KePr4aNWVQn5hOwZXX7MHlJUoxQR1ovoJ+8jy
oO4jMLNWMFdD/ZUihIYdDvqdwMFfRjQVfueIHZ611fSDRxUpmXuXHN6zOroUp2er
PyqVvUPojFUJ4LjJemP8yAoxKqW9YO1bRZ72+jLjiEWS/X1pSm5ystp/c/viOTQK
txy8QbnCPprwgyOvnxtQZO0qgxd3M3cfI397jzJBvG5Vd6SkhhbgLTgSNhsqeWDA
QLPpvwOzluCbeZEngodjhxYIVRL6DLrYNGbKNE7cJooWxZz51oyiut7GrUZPE0Qx
ZY8casvF5uuH+Zsu8IBVOHY1mZJ8PA3AD4S+Vn84JLy6mPWCLduFnfuj/s7cNxuO
KsH2xXLzqnoTGSCTHjtprH31RGWbASSUGudoXyccAC7Slj1W7eUIB3CrzU19juc3
lAJ2MkxX8uJ13j3BOs4pKFccHdpr3YICI4IaF+hClxMbcWtzo/qtXo00Tz2AGidP
cFXzpWfgVxbDjjbHYbyWeyDvWuurJtJ9uBmSZHJnxPZ5+Pj2LBwovZNxU0OiS9t1
vezi1PBF5gPQiICVAQft3H9oT6gFM5Bm5mAb6UsUpgHYJvEPwd4BlTWRoGP5gKa3
4v/KThEdulmqNtD/uayg3rBfsnrXyuTdIp7WMVyu+6hDZhPckmnXVdY5mjh+cyRQ
dYo1KHJfac3kqUeM+oAh4pfTHvB5gBiXbnBU1evDus4nINmUpSRRjm0e/tAeWJpc
+loXiugyhA7fe6CSjy/n9HI7TZX9/1HrZrQ7zTAvfC/7Nb2hwufVEpBg4LrmrcUB
alcyLkF9Rp5El0xbwRpXJbsDFv7LLsYB+tNsavZqwVx0rlwhbulvxitnQRhjhWkl
`pragma protect end_protected
