// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aqA4JNTASh33YLUv5OIkiHRrkf5NgX9C9YBD1ScRIIrdIbmJyQGd/0jW4UhcuM+W
rItlLW7lZOjwaMEUvNMkXarvxsc5gqs46tSyazYLPViJVEy28Xg+8sP5DXCkUYvW
OvDX4ycss6FYx86oqVQvQdN4YSKscz4MBUQaIrXKXGg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18016)
d65RtIx0YryFeNLO1HposduuueYWtQoE3Vd8o7DwYUssVA0Pbp7lMOOd1gbyTQ0m
9nYi8FGA3A6S6VXlNTLJhdINiDx4kEo2SrKjB8SYk0y9MYCCxJwdjjQLr1udFhou
7CNb/SPcwrAK8Ye9xAKMsGvXFeyspKKoe9p8Q6kJcL9PJ4e/r1z7k7x2Dlnuw1xP
hMy50pPpOS2s1Iksv34J5Wyi+U6AKLIEuBM9QmheW4tdkScsBu6hitPXWAZN18FU
1U5LvPN21kkqfbtqPt8xvK3iMh7+LbcMetB9VRZB90Q4+5brNGI7aQHPoLq2Qy01
/C+m6XCSiLrgYjH84y+whUNvL/yDf+lZd/LmPfQRUkaVPUOkImiGsMi3c3Svf26o
y7+yzBC5ziugW72pBx6hfOM/xl07xd6AggbE+y5upXS+Pnm/v2L9Om1cd0dH+N3y
tH5GnYwwdvplb9gAUCQCsrKm5LsSgnPuU1Dz+hD2liE9oiL/BBL7m9t4pakwQbLj
GWs66jv1R555QDIbi4E4JHFrRrvI87eYUFxrGoZOOnASDRSGvmZTbmha1mrTIfWz
ifLWG5p8EncMT+DO2v6JU3Cdqjz8Oml1jAAZYZpOQEo4s9MzqNxt9o9FpwS01KEG
0/6BowODeWq5oO0AncfSpz8fmDCgL7aCSTbVrNPwyBVW47A7G2t6HUiyrvxy+OWN
495vLVnSf9Rbm1tTUiagT2W4rO8DTKAB+WHo7OXjalO3zazT/XnmaAVhpnV3bkJU
MWWNc7eWOvCfy0g6RPHBN0R5HfaWLjj2Db63bL8LnaI0BOEMbxGADgxNrderNTao
pByyTGGFBk83WBLDjiEvaSr+uFtaIdEqoLwTSR2qm7zSvpahnrS6R/sdFw8uNN+W
YCK09LGpadXW6GBcz48d+xG5SsL2PgPGqzgjWtgSKC+Es0U+idDolojiTx3gr4nM
u9NypTsaYkMflfLHPpMxYlfCv1FOHW+713sqtRXvUA7Xdww/c7OYogecEM63kb1Q
pfkp7gkhM5LCl72hrn71qT04acu857yOpz+cfCV7L86fSqEML5QwrVVuWIAvAWyJ
07scwkomgBMEX5pOi0H8s6p0aSo4fC8iczmQ5wYev4XlRv/8gFSK8IWAvM6rZdwy
BOcTuNv3czvbnrPIHNzzteUvY8p3QQ2xRtlizlGg+DxoTYTkgrpIsm3zR3l1Jsdx
rc6KTc72YqFtksGFTavpwFUmu/OFK8cF7pRSPNOz9MmwgoTj9vNf9eHHgDLz6cZb
rYK2ybj+rPUfy3yrBBf+dpqPG/vDCe6B7/8SZT+KWQbu+lMU1AiirlCWQNgqohy5
Oxuefb0d8u4mbdQ8fVOE0o+3UfKd10qT63d6f3gw66td7A0/tayuTmmAAWXYBk+Q
/GpUWzo2fzkkUbJy2Qqu/1rxXHs6FKHCi7vcotfmJMdh2RwOQo+RKbPz+79xccix
Nea6hdAIfnkI8ngksdhGALrq7XrnYxYQGNUmf5sI/kN8nZgUYDoxWqH/kyEJ1VTM
xFPb6/66VkjDGKMspy7yHul/RYIlWathAjZ4/j4+mLBAk/qdtUVvycWmY7duz+UC
iU6vqETwQhanOGPKpOtoLuNDFOxJTXH/HKRBVWFc3drjDplmPewf22ukoMSbURUk
2nukFSlhcrU5QTJr9cWMrBt9KkbgUwLmhAJ6Bgypt/i0V/QR286zamLwCjy6jUqe
5A6gNBcDkfwRy0Z16m1uKmTQW1ZKrGowjhlgescAGL7GJ5kXiXIrjtMAdPb2DtRR
J404nJb3PoG8ln5NvTt5YA9G/f4wGjnpyi9O1mXUhRoWmg17BHH2qw2U2Izo3Rrq
61wZ9/K7kh6fwRlhktzykOTEQh8x/b48j1NoMJYAoJczaQHhRVfIramSC4GrVODW
KbC1yFBHQWZ8t6kQCZ6vzmbG7ob7PW1H70jLhNonTkzuGdt8m1Z9DKrZd47fDFe+
vZt1TnqdY53/IZxCUK+rXWsj6U2IDjPvUGHnKOX8Gf6IgFJRHXaKS+z425LRCy+8
FiSnwSy1fO0jqA7zcFlMj+ByjVxzODWJNe9RjJYk8efZG3WR2LbIZe8TMnLrYWp+
A54FmUW8BXlmKab9S1BvrdD8Krryh7ryB1scgMqx2CCd3PqJiLLveUw1dU8k5tST
g+StACxZZwm5Llz11Gjjzxt1/AorfLnay9FGWkF34PsXziHpvDxEX5rszlB6/gvd
EXKreUVfVj131Vtlrhim/1w6wN4wvExWYbqalnzMcUxLvybE0nKoHJFuWsysHPWn
jJAyA9mZLm0mNF7skOQKzT3V7acXR26ut+GrJ6P+9/s/2Nq5OGrf5M2MPafQyp5X
4xaaif3nvXSJO0G0AAbHcKOohYej1M17GvHJCDcPUAex++eXdtlRVCJ6BU5FHPCQ
rAuKpEvG2o+euDC2eO3OrrqMeqxcfWWch3Si6uPnm6TIzWpP2AyN7iw2Bm4Gcxyy
iaEc0zIrkxYputisp9+HU/qXCTDnEC8uNOPJpJCdccV7Ewh7K6Yt16AjG3YmDE7H
oKNbrgAa4ljVS2gF1P3kB00TI7UmMCIgJf5cJIsdGVc94GUIx5tjckBMe236G2Qq
FRzWw9pln3LZiPxOcuF6WQl+8j9YDZqBZ/m+cQfeqNGc+ZWmX8WBfYSm4X937Kut
9bh5U/IRifgQ/WWhmKyaOr8Dj41lrzMb1r6vDhTQuXerTX55RGDao9VoKoKdN0cm
YSINX5FoFswpIj5iygMSggTwi1jC69zskfqQ3fNOE06afhGzMvUwh5LH8XcaMOA5
pg4GqqX0z4BLJpJ9iIH4cJSuPoCICz3V/PZ7+wg+A4y6F0UHwizzB5uAN+bLmU1I
O3zlcyEfHyJ8jssBUh16LoDcKnCUVVm6ErOs2QI2A7j9tvJOxUg0AENj8MzZqQHy
HgZzvyxySArWKKO9ziwCdcqf4WOAPwLiLSF8wC8u+CBxfx73F0WmOdNYYcVhsE13
CjMc5gycZn0T3tBlOHZiWfHmnbgP206ewX3tNIHnP/sztVaw8LkNNTyl46ssmfaq
lDKw/8ssYmRg2/oW6xWGrJUjb60PM32K451PX2HN0a3dNcNMZDZUjSaWYL2ObU3U
IEmfxsEfSSc5NYPE2pXAX4rYVLbjhwRUHZDmZRWzZBmcNwuEsQSFz6nz+PW1ciz1
dtp10+qyQ+EIcm/x+eLvOXKDQbS0KilBUNGONcMJMbp2hzy0FJsAtlPIX/YyJiMK
gP02j8W43Pl7Uu9zWNP9K5xoIJ8m8fKA0JrYRNpyS078ReqJEd1WOEfyAtftHFxZ
gS+zG9XiP50mC9cJVd/ocXfALYDGuqatfoNed1b07h3SYxCi1M+O1tGxN86J/eh5
UUOJy63bAOHaSSModiy75e/luDYpk1CApaKNqLtu+xTH6x+lni9Gnr4lhj1w5MwP
OnOwy0BcYNJdpEeLVavlP0zvjQAhpn4+fu1vlf3zQW4KUWOhU8SoAECvbrW6Y4RX
rHt+UvNC7gsxrxui5Bz2jMz02wn5SYthC5aYsCYhNQWiqp1LtLrk5rpz4yAaBEBB
cUcnWVWiodtMNJCgy+gYOdN/Bx9DrdYKdwIYuZgpwEP67Ooor9nhqioBAhq077NX
zUTYsvx/md/eCYzratZA9SdbB26g4qq3RnE0ENzCjMqxYydMZYdsyFt4CH1Iglfm
HcP9Dth6iUaZLHi47ygjeVNs9FY+iaYTY5T38j3yD0WNcc4nMXU2t3bRMYGQdCqw
P7KawqbRUtpSzMP/MnXTfdCicFKiinABp286WrTVHeD0vvf8mE+Jxy/FqPQhvixy
sdp26SQ1g5nJMYBcxROxtgof1QEIHCt3IKMOdGrpRh/llDh28BhSyGKtCDg6InZa
lpv2SXN8xM2arKCs/OOVRIXiDDjqwXbIQ9LPgGU1o99PQBeq8Nh3mpa+ICAPvWcu
qQL2GQ0MYQ5McV4AKSy/NjiM0wwzvF4Q8f740aC/FEhxpXJDRABsf9LuMMGEve8y
Qmi5ZEPusfgvraKIy8A19Jr7AziYnjzCV9YQyMPfJFQm3b8k/rSRyO49FCH9wkfL
/6fKDqujwmoBLbeHwtwg+YyzkJTIwhJjb/MnXzGqce6BzEEljCsc5Mehk7qUsgBN
x7NsJ2bh3kESCvt/3HEZLGNggMoV2Dc/JHjnitgiTIAykBgrKx4BBYsJmrMAABma
+5R3wD49uTjyYyWDtBBR0qqo9xDWowwmhwB5Mcxsjb/IlpY4LdawgGNrXC8IqPFy
3IiTzSMWMm656D/QO98T92CbYyzhSt44M4Fh6u/iEs+OTJnvFyl+DObPdk4xPEuu
tZoffg0C3BG0n4qv0qibIFUaXa7h1T0c6JzKpBtq1KMS624m4qarGPKdVPS9q8HE
8meDgHx1pSZmHY9vZOXcMdqgN7uYGSiJygifylaYGP6kC2y9EMZHOd6LxUbcCPGJ
J1a0SbvgJhZ9chj0PdBlpyTgff2tyQkqUIqTPa5ZSiVTiYK25SHNEvJ7o9CXurtz
Lgl/lQxPBt2jt4zii1bsQfEpv0mGEf07nqdrTySXx1vBQdyq7kreYmsjmGvBEgne
NVrX/BJe9KnJ0xRiQilrE2Qs2lJGijvwcQNfUuG3lM2Mg0ZDPFgTijJfU7TOqQ8Z
1+e3u6aM+WRL8uhkkU1UPhe4noXTOGGbK3ZMFHfpzDzyrBXGQk1RU2rYVWgEksOf
WeoO1IblMnYAOlZ/Iz5vStMge1ywVZ6oJQqh2USrVPx9masiNDs6fTffmP08zCnV
hW4IWzP06n45oVJBVgRPpUGH9XmNajBLeuZmj/YbXWwysTuun1oTayab0xXkIOs3
1IHbia8rPFwmbGLAHhvFRtK9buWHUidXR6kVw3KegZE0D+M++NSJuzFq39SklfKF
SknJ6a553LCsV5vPuGlXhhTVtFVQKplWgFXn4tVm3GECLteKvgmXP5ON/+XseP6W
U3L86NQoL/5iC8RVJJoh2Qgc4ca5smfDiVOHZNeNqinbgM+lfgSRy9N/dDliWb8U
zaI13I7oP2l7YpugAQaFFTLbnd88hPILYoh5MhFoFNoNQF7qBiDK2926wlZQzGPd
1nH9Wg6jONAw8+t8Kv2WrdGBfiFCVgBobm+DxA0I6nVkFLrrfRq8vWrVk4E/U49K
KiRqaMSxFSyCowYJrVUe6W0uuUtr9Wn6Qn2vFb1eI+wAK409Pv5ng2iNi4A2+Orw
8fQt1k+d44Yta7Frln9UOdjUuLKTbpzYSOha9aE3FwKmlu/mW7px00yPTlIX6McQ
0gW+qb4YHg02/La7CsYeNCg4XaxBir203kOVKy/nwUtrNNiKXoe3JvCVFzSfLoR8
Ch1rdYoPXP9/d30kDepg4MXK7fKcigBXSVzeFxJlmlpbRMgcLwCOpdlIQuzbbFfk
ckCw14eHz4kyypsDC1BD6XFAu/6eIxhCTUy1mVmqthZE3GmqX3OypqEBw449TLxI
LTYqYqb99LugVAqSP2kB7Jnd2dyAgSMVd8cOQPw30TI6rkzQdjOLOtDx1TIufZ56
1Ldatid82wO7O+ZbhvYaZjt8G5Lepd93kmYSI94rTd/cCTNHDhTJxYHehXYnI5i5
VrC8svmnLfrw1oNBz2JjgaxZYLXU1N7E6e7xdeuHxUIaXQPoRPhAnA9ddAdSnadq
xnfNUZxuvaF/HgkzSRmDMaTyKTL11BnGAsWUTzSbbcSlVFwj/IgNHLklOofVigAm
XPzVJs0J1dsA3iR0AJ4I4gVZfNVY9BeDR8RJGE7VXCGRXgmk3/ud24p3HPZEVrrm
oOtX3TCBwcBTsDYKYyTCX3dVn8onDwDhwFCKowx6inLZ4qeMt/PDuzy5fanN7wyQ
ikWEjs+bA/1dJPC7i++RFmZLik2t2WghyliAlBqrvF92so9fWiIfHWf0y4Jw6Hv5
+9Q0dgeRcIwDLtJRL+wJ8Ums3doyNJwtYDNsIYHcsTa65fn/dmtsTQ+qtWK4pfMH
zjlWWAcFdqJuyO+u5UJ+YI1usE/FD3PX5RZXRP1ifZJDWeX8zJ7irUB2agrJMTwc
hU+6vCl6DuYHR6oaUkQVUfHP4lBLp7lV2507z4TFSCtzni0el95El702EcWR+8ao
bd+KP7yIIifrtldyoFHgYf+VJ8/w29PPKyZf5DRuOnUn1763W8EgTt4zUTIYppey
c0gLCF/0fFNonC61a+Qvgqvh2Kbv77ofToo8W1J+pkeeJDcGr1Z9t02XF5w9IXNQ
D9HOR/lBHaYqlqFTYSVqpV+hWRYO4wPNKw9ph1N+GrIS9308IRSNDmukU0ZmqLH6
dYfsdUEpOvR4G6czO5ps8J2ousbBeeujJ3qUwtsHsUdTeT/pWalwt2fq0TxhrWSV
TZUL3OUvYIrX4BoAdxuOVIHnfMvVfr9egF2vv/KdQI1qGegBAqbTdRiEXHgLex9N
klYLsoZS4qy/exJaPoTLYUORGQowBOSNGGoDy2K1RnCsoWBt3PcGlMrhFMhAAVTm
tgtRzXlg0mqkW49PknFKAapmm1tY5tJxKLVuWw7usEw+ASb0Xw2MSNOwXe7C2+F/
12gg0tWO7QDktmoVWScKAk93rSl1hwh5Vp3rkXK8wOpSwl7H8O2u2bIO6xbdrw3z
K2Ext+PuprnmwZvsWx0mLl3uL+aiIToJgpgmu5syNUES368arNT/FdrMQ57193sY
jc6uQjZcmZkrizRLmpYL8egYg4OUGGgforYhCSC3ScYb/mYajJIKrHMIDKKQa0CM
5Cmj/ZMMrtdSOu7Ym9PkCnbyPSQGxwv4ClEhZ4tNJRMAGzMuumLDprCkGkDc+urc
RzcptutcVD2cECARlRSJkZ1rdzudDiVClGNF3K9it+oNGRdZWGsfoIxAX67mSKHi
Ji+mQZL5geKSTfKgloGi1N7Civ3yVhANwUeqvtWtYVeofg6Jn8fZQ5xrV8Bu5DjQ
H2wdD1B8OanxWf3YflAT7pjKkI1TFpfpZ13yAfald3A3QPbOrkI/6cy5gPOgqgLD
pQdZh2gP7XpUzhNvng8qaKGfSXhVuTjm9opg4Sn+Z1qWBerWwQDLCRO+tyfslSp7
NFeCP2n9l5OJyslUv4WySs/V9W4Y3kx0PgJIqqZuOFM3ririjch9BxUs/dz9IUyi
h/ZQxCLGl1rSddZSdgRFb6hTS7MaJ69yGKMa4Dqu/zcd8KpewLtNZP0ACSBne925
aFgR5IeHyB652VGvZpQ82Vy25Xqm2KuvMKS2rvSpt3E3911y88nw3NkUB3fhtELr
cMJLPYBXTDCyR8u0tR21tdxVxIO5B0bOOmEN3xmGCoa05i1c9YLHU/6h2FZATweT
fKsKDA6XrlrK8PEVjMr4yE+/fKloUsqFSlEaHGdFlJYErg4lUMCOT01TbxAFx9a7
tGljUIxpdT0ylP++I/guaV7o2Nh7SLEgF3TjqpeDKiQ6cACH4crxktHUKxHRmDR+
1Xau9qTRdcwJQj1Y3JRIb69/vGpF80YFsvPrRSDpmvdkxWnI/2c6imTEKWh4YpFV
lc0w5eH3KB/yNWKdXoM9lIeH53PnQGFJfUACPBOGrzzx7PMA2egFaDnpUnVnGY1v
sXqB+dJrkMeq4uVuEcBqdudq9Jo/FPt70B+Nj0jQOdBc/6LHZFadwZTXOOxlUvJA
UzzX4gkrH6uWCJr7paeA+nDXF00silx5edG+6LRD9iz+l4MYAdlzFVtUHVG2ELWU
XPo5ZeDddM43xEGLrx25uDX4Jg2kouSWLJulSmIs9/7m2vdjAx8JrBHLlhDGmI2p
He8ELA7wd/ClNJ/qIJlvLjTfNOBqQtcYk+UMdzKcsLx1UknWDBt7gBcXwvSYYMrN
wTDngBburumzroAaStUzfI7ltqgy+QZQ/z1F7f5prY1/Ii59gQskMv8ACHa9Ws3o
VsJj/lgBC7dQYLSJQuT2FWG33jsPAPmGKfx3Qx7jeae2+nu7l3F5zQb9obLJWjKR
PEc9zq6mWwHeGu9XMsEa6p4LFyyqot1sC884FU7ur+FnYZqQ8HJYn4RvflayCTrd
VyOmr2hKSsRUAS4qMroI72fKQ8zTKpbMMCX8AeTNQ2rLnXKIBD/Qmi49OeUj8uuY
GV3kKovMmLYoAu/Hak4jSfAveeWAVG427fbbsZvlibhu/NFzqpDPxi4LhCe1Mc7I
wjUeQ5PximGVQ+NOxHvoqZ1Fzmw1/lI5GSE3lP4wrmIK0xio1ztsFnOBta/qlafl
XV4rjF1Vpo/yB5QjQl12CvLqCwcdNGhY8ioaiLf9G8fXe8DF5QubbgSv3JLs1yVp
NODIDIVHpLShG65GmqJOiUAhUpXM6XRrsH00isTwdOPj5erOVQT5u6k3DXzdSbVe
o5z+vBrpmCIfOyiIhoFWeN0vMM9RhvurJDtV/rk/wGkbmfjUr93MSXOY1xeEMl2N
qNX2xs98dE8nmDpU/q80sLsD4bEvANfDmV5o4/U4F30RoP/RlAzZXaaMTSisP9gI
gKJwxRZDKK4DYqBCYlTlZJYDyxpuywFeYLEp163KnbaaLae7WhnfrL2cokGDkL40
R7h3uwKa88LNTM//CL0/odH37JuM0Bpu0mxgPiKSGTiUp5bnPUAsdCHLaydN35EL
XVEgQl5koUfICUvV3k2y27bQgVmq/NhCq8eS4Rj7OK4P0YIpk0ib2lIBWF6C2rY7
4gQEkd5Sb/hVCGInph1L27uu8nKEFsZRpjPFJPvzpMu0VX89+csdt1+Rg+XPr+HQ
BRjRE6pOybTgrqcLmWQRMvud0kn5NKejoZ4iOFM61RZiML8Mi1uPl32QaxVruUAn
+WQCqqL8X+JQZTYATMXJwDNe4iGFTKmpS+5X6RQnJD44aqQfYXnFVzpFbZA8JEGj
Ufxta2PWX+SyESvdasfaPuQPcDCPkO6dvuJ0ICAFoQuWAnBI7Z8YFjitQ8vxBAxz
CUt00txBwmyiwtvF3XYjfqe3Q01wUN5E2MpEbe6dsu0wl/a3rVoE/hAhoVHsuGqZ
edf/ND32PZ9r1guoMinwbKo3VxP64rJTwvi5hIruoRI+M57XC00CQzDkeY1f273T
YTO5O+zu9EpCioHotoTeiPpQerLWspJGQQPT8zB3rNYzHLfi+adF5mqnm8KOAxiO
bmQB8h8QuhidyGZMz4XNq7qT7xFLUUBJ0lz8BwA553WrUy/LDx72QkGaxBuPNDG0
LKM89i7QMhSZycCybKW2qYLcomCktLQ+ubBvkvTyNkH5rNUn7bpbCFb+pap/c1jj
T1VmDjhEWWgoTVs3HYsrsBKVC9n1VUnjbBwBSfBzrAxJz3pg8/eoEAsvz2U9LT+n
X5I5ujq2/BlU43+qDLMYRA76L1asWhHgiABYUi0p694KWTLvW1M6r8wKKI2hpMGR
VPvMkUnZPlwNjPVBParvx1JXA31WGqT7kqB61+rr99U2/GWCsobLjuBNWE2Mm6+Q
+Ta3PVZiAYLZnHDxau2toAQer262G74aoR6kXpiWnzuNJt/GLVr1I1nbMTWqkl5q
3BeDV3wlFlB1Q1NH1wsanuO/Gl4cUmKqXsXzH84FEzO3REiVmAr/yGGxW1jE14FN
cddHsGkYvTieNV8sq+Dh2V1J7ZiPStVILuMMnVfyh1BltUbrDWm/ZGb519f+R39Q
dzhJFyaEb1KeBCqNg0fi/xi3TN9DWB3Xe1MZUmtJGCgKJWQroB8BSrT9VZEBRyCU
GEMevyNexi0xH8Pt5VEMzUQAI3nLPXmb1eBYENKtMGN3Irytw5jEItTUxzp2otQB
r6Lg28w/cvyGGVUhs/VCTsdz3O7AcbJvI/3HdehvgV7miahrkooxWxT3cpOeWry9
7orMz8b5eNoQiRDUQ1lSPqrKcSLdvwdnOnh+/iKw+tIVCGAweyQrrtOWvvc1Ubq4
9JKPM34q9JqKgxL7Eg5FuTbLiWYFut2zr4b1oWziMp6WT30nv8+g1AYGUWNVV/vk
xmX/L5AEIkm9yD86C0pxjGzDY0qQJ+Jbo0s9gTV+7fnjVh5k0uVEBOl16ewBnB/W
kbfvqJs0WQB0z8vMYBt4zkG2D79AX50xxF7JPwp9cbA05AjZrUHRCIl8c5Z/AtJr
zB+YgAtz7sGdlOev3LupJyaKjPdhAtIU5ZlbnfxNK0qD2httKGPEU1sTYvR3IzUC
ep6eV/1GG6dRoG+OU61987wgqV4Dpcde+hZVadyxd+7GJx29HQtPU/WJ+11G4ZMS
gGXE5e57d+KuBmu3BKZW5BNcmWVsA0KuiowqhuGGE5NpwRUGZCcjyKhqdSdPHFuK
h8uD/78Z4n3J4IzFypB59nu5AWu5qkc8qbzq7SyBB66GPy2eJbHM1iBoLqfp9v8W
zr7MmGbRf6DiY4TbCcWOKjQ+xt3zxmmBkYiIEpXRwRKfsKSFFf7DiMigmVUqRsWE
ukVZpZ9rfFks6lZtGMB4gGFp3TkSgYer7skhF1/T8u3kx2KV5l+ieRjy8r9YNwCV
bapomamO9u8yZbi5yLlXG56KTC6Q37qZYsEgrm7RB6xiDQnmysGnYdfbTNYl5Ure
2xgDNoI7nqnUtWe1blhLj/y94FKiOzFrZV8g8qF7amH9dc8n/vlnEBTmaVtB6Odq
uZMCM+b+NQRv2k7sYEm/wJ1qly+kcl9X9ekE8qgJ8QbvLdpGbPmKllHDYaDFriJy
b2qgIbz0+SC+QKf8/w/v6ajO5FbHLTvM8rY8EqiteUHC2AVg2loI7083Lx6FmP4v
FZFWSXCcagxZp8J3KS2m1dMHtoEWMEehyhLkTBJF+ERA3vxrpgBv66kwTNbL+mkk
sBwAAyLw7HLzYCiueMa2kRWTmPk3zGeMqhv8kAROKH4EQdjjfLS7E9Q19a8VyEDg
jscQrP6Oc3luOB6L7UvNQLEaiqBvUrZz8uiGk6XhNF+yEvtYtGGDSJaJ7RUrW/PC
5SU2pFYvW/LCatRq7Yy/xes46Lj4Q72bJ8dkj3moI3avqqKclhn3gK39mh4kZK4u
iVgBvSmPKwEVQ3bV2J0NOcgrVQdrcaSExNGrr0r2lip22VF8wycrHesMW2fvMxjD
94M2XxS5xfgDDQYtvu767Fw9gIxf2P1FMhWnq+Xt1wZCo2qddyMDcAEG+JDG8zXg
ttRzXShacEbHTB+PCBAcvWL+io40LJQx6h5lPlDLGSnmrJ0XYOO9jC8dy1Ufp3mo
Qz9gR+TpJreujfsi5I5nEqLg0IyCNYHxDUbafnz/j0nZO9zbmfj+Wk27pkh1ucoZ
K1mFSeqy/3TE/prxLL7Eg3iVJdbZrtrrzshr2+JXCcOSb2ZkoAFxuJ9jVninQ7yc
BCzRs+0H0PJ2zKUra1yA5LmAuBcuDbX3qbn6YSWvG72sTja/ZXQzcOULYVYnEjPV
sjxjiaKBUn17kwijpavzAtJlkaqjsHlGRn71A0mc6D/3bEZwfJmCWWIjts676VhN
aDg0Qs4YmhfD1InizSBSQDtUaFQP2TQPz49nynSULcV2/M5AM85Bx3qGW9dOINuw
cWPZ5YNXU4Cgzk1Ol0gh8W9mrfZYPcdFN/4irCuN841iLODuIv42pxxsMS29QZCO
PmgaDNB7llwZH1LeZZIavOn2m3MdSgukwrVTB8gnPfd5+KKwcYA4Ri+3qyyJVAL8
f94PErJlme5ArRxjRZiT+MgjI8EnbdpKZ9LfiAUW5yqp8OoqqHx/44XWe6QRuGk7
AwxhrlkfDycVMiYs2Eg16JFRtLoohPM0Rr7JZ1piS0TkwG99myRFIg8HSdXGGssr
dgeQZ6O2lIuF2BA5Ao6oXWqJ38o4PAIHosjuZPBPihAoA1H6cZQaDt5bPtLgPM2R
k7x/xg4yuX7huzWCSoQmL9xk8RYZd8mCOtKePxXFRbF+l6VFP7pfX0ZvoUaxf4BT
IYw6s41ACeyTih7O7R5pusmDIKZR9uJCuqhHlrJNvnrTThwW/BVtrDKRQ3BYRijh
1PTWR0HRKG8bTVF4WM1KwF6hU3zW5wXNN9/JXmCEm6HEP/Bw2GfBHHs5LRRT1hMQ
jxNPaJsD1Jy9Z1HAbi72vDz4e1kEGs2haM5HdDKPNnXQrs8MkdCZe1b5EC0njTCZ
OZt0KM4QXpztL/0lKQNBgxyoWwSmB3lhNmjUFPirlVf1dGd+y1kBOJqJycBHkJEz
zQR5XkDTe+HqMsPupmPC3ZHS7tMa9G8WOVzHXoILvZzriXpMtdNdJnKGYBeQAQxC
1NImF30w/2LB7rQ5Ky19AmWgYPzMtUho2iUbj4YjHEwFWxEz03bGJ/JGjhDxsn8P
2b8gJnfWgD836HKaUCWT9Iqj15bvrGKKstDd3pCrR4s9On0h7Ne52ZAV2eRkqDdD
yqKAQ5SuSQUSZfrboNH3nYSxQH7g8mO5jMLLbg38gQ7tViNhhxXuXb9C5wj4razw
swixu5DzvVYCwnkxKc+AvUOi5rq3PMZx5Tc+2ZSWUM5FO1mjwMjYLTT81nZMPKwQ
F5/7ySL1OqgzuV9jLdNtIkFu4wAvS2MEvjJ1kKBb8iJYRVuCNIv48NmWxKcfmwjQ
FgvXGqoCcmqOmtkiToZT6pFPeejoZh8VM0cJ0LJz4HLmI4CDpoMuggNGQoA6C2wG
naMu6xjmJrVhBw7JoNPEbMtNgUa/6Xi+1UGFQGVWqCoIgUQ7bYBepyQlEt5F2odN
sQgu5KGM6I3v52+dIv1y+fZS8GjrcE7060XjOmDKESnW7syzAo9ZpmEjnb5/xZfX
5Ple8a4FUM8BklOFhD4dQ1fq5ywH6Lyq/2ROS2zmK3oVTaDaXWgcI3tQBjhhA6LJ
Fua7PJk5IlwVDquNA21BxqIPGfN04ur8lZ+UAZok4zBWo9e+tHoWRErkXk3/DXnH
+9EqtYa4Yq/sIzbfXPxz5TOn+G0iwVXmSDe1FatrqXzXw6rsxab9nUoD4XUq9YqL
H0LQO3B3IU0q/6jiULL68nnd720IWsCGN0hXTAErG5iFQzLl+c2C76o3nNUXEN7T
OFIkH33ld/OxbN6vI6z4CYr0+WtA5YqxfRkL2j+AuO4ckoTM15Po+X5Zmi1mAzp5
6CeTZYKSQrrFurMwPj9DJzdgBQdYFOBGkygaAaZDTWN+Qd6ykyo/bKEMAJkIDWgP
MW9zeUVcgA3DBg6b/TxtNqeQ7jKrkq2cjqlm7lKALVJhJTcqUmuVRUzxaXQ2t2Uj
Scd8tFcbHerEawCHXjyR/0jvnJhr394JO2HDFDVTUveIoFg2uIf14Pz74bpqCjoC
LFARKglePL0fwTxugoaf9f+FRdfTrP/DqzgKQhxQf8TfD6Di9sAKGZTx6IoL4kQC
c52Pi3Ii/7OVWOmcgc/yXhm+mQKBfsDufpT4puZM14TNFqeDyc4Cxos+ajPzmSJZ
CcnB9BdGoiQMVle6I6i7AkE5Map0ZZrk0Q8mu/3U7yhr/X5gE5S7mIVmmmEdIyEn
ZWGsgQDnKynlISACAcInCKpOwxOWi2KM4ADnIliNESAMK9nA3oiZdyyg19Xcj4n3
wCeNmXyQj0AjUbyQbtArh1aGqav0P1hgZGQ513gC06ty22TfhfmH3SgeGVGtuQKW
o2dAAUOUc/fb6735PJfUlvcH5HxugmxUXBdXhyUMMdqdEkNL8DAr1iZkibxCkjH0
lz0McOlOkFJ1aJ/yphpOG6RUIrnwwaNC354tuxrfE3WndfIhSUtwUBEKHApWOLQl
NN+oDPgNuwZGIltqTfK7MLVLKjvFwww0S/4JffxSk0oC3wXbAa/mjfNAU8GCKn46
SPk4TlN6nwsNyfojbH7AIdePuZF7QxXbCdbrs/KIR3f+Dv+JpTYJYXlnDHaB3Bv0
EpN3yhKuC9iLwUoHhSbW5535aDg8KHJBY+fGRedHUX/ZvkjCVsafjYIF0OsVVaRo
EmTE6XF3ZodhAPIWsthQDv5xeQaKhJ12iqfErAOOQyB8uXEyOrssO8DRhruAWPBs
yOGlgquqR1bNFcViuQMViDX3HHqoPLVX7NsegTI6RQphDjI1LM1lC6IM8qk6tGf1
mRIMA+3mqcfYKCRAOsgyKb9X0GjRk4HYpvdCNiCOPXQiyjY2mXEEIQxUopeBNH1O
x4+i8JDmg89FKw309Y8RCSWC782LWFevBFM5QEdIeLLPXc2vdoajKh8+58q+GQEA
UU1V+8wbUYCAHYjO3psqpMzZG4sQNX+InGMHsAgsxgjYgVgWGhtlL+5vLRxfqaAS
c63BAhkbAtW6wj4O80CdH8yLz3drIOTe+gbEnlEddR8DIejyWb196oFT866SxPuv
KDv+Q0pGPFGO8qOmLJFaswgRU9HCwZGtOgL5qOkmWc0tDP65ljYGmTmSb/mojtPN
GDaj8BNJgDzbOIg0iTkfx5ovhW4U18nVl/HSQWwqjKLwVLeAS7YgVTAKAtwVGLHU
te1h4DkqImSiA14dPv3T5JWUDMOxjevZNsH71Jpe97oWsdMEqIIlck82FQtZ09km
WFVy+RPzz5UoGruVxe/VQrCO80ZPQVCOmoDs6HX5t4U9tFKU4MpHtqvK9pTCi7Nt
pNBt7UVNHxYU4XBTJ0sBHN5C4vgLYnOX+vdztCq4idYHR4xLliSnTJXJV24uc3oo
xbrqP6DmgKKsf8gHev7c98c3azoDXTNzYm7QuV8FP/uUy973S4KEc+oTIDU1EIbP
nYaSzHsCgqnJWompH7VaJxZlc/Ol/b+BIxz4OPdItSwCwnLkV8UohcDnQFrNYPGL
xcy3gDelUNifqGiJLUJM+ZPanxVZMe6gl/HEoxLD95StN4Tk69OtJzB7SY1d5wnG
MuuxldA2IMhlVFr3A3fsi0j/TlHfv+LTm2t3YUTfAbtUOKfjBh+FpXIavfgbzKnk
dLPHA+YzrJ9BWfmMylv+7cln1LKAGXViCwY8f2CdvOCXBDW2GMpGrD2b2DPyyZi4
TBtXZmqSCo6vKc01LWqutdbIqldY5YUIw3z7Frq3CA6ypdfOKSlauxUjQ4BK8wZG
cVOMW+vug6pYDo9wit9uzC4gcmjQ9Ulo2TyX0rBJ/FES/6SITZ4EXvQ8sE8/qBm2
5OkaUQGD2j1RrjfaftQZQ1FbVkuPLfqCbX9n7JJlyoVp3UmfgSP79qytr6z71D1Q
FSOuJR+OdfakxllsbXAPSNaFaHtfCLptxG7MYOishZh3zuquPikdHN6alV+gQVXo
FF/X5WyTOgm80BU681eZ2dkSjoVT+acUvazCOQyKvOejNo3HyLEuj+GLz6uQjegi
FlTuAS8jF+GvFycGP7sfRh+svXo3vkiB06lRbS8aHCfYJMjxyng+pb1maacoH2cd
QIQ4IQQzmsAYWC2icrm0hj+dyIE3wSi3s/yXtBNlxt1cNhrI155LSlMU4wGZiQaJ
3ZfXUoAZKtSx3/avAC6x3ZGXDyjDAqNVdxUQbXBGoIN0bcfaM9pSo7lSMzH+/WsC
CKtPL6effzCLwv1/OVcx4XB1EgQQQmfnEAYzylF9gQl5osRQhgxtileTaYJlWmGz
ql3LrpucYr1Hk44/MFQr8MtteHxC6d47+0Rov1bGnEGtXdlKc1DbWpBIOyiyNmfc
jnWPUf7bxRY1CJkKfjdz0HawbPoAzhU8ryXJ0ztsYixtMs10asPuPJk5Trlr3Q+6
lcpZsdydfstGovdVJ393TcZdfTx8DI39vf9mE7aLjqqudCItFjZ8WxRFZz5sEqxm
KMTMxFo69sjE4E0Cw0D0iBwxMQfFzJjY3zXnmJdb52PmYekY4nBX3fDcSFb6Uank
gnMjGExCAn35aLhuvljo9iwWjpQDlqTvjjdQrBFcnMc2WiH4PM8u2/mFSsSrnPPC
IoMiMc2hYUh8QhfmaIfH9dcM1VhOE4pNGXtvzkmX8YzusLa+ykBQ0x6VTIKIcuCs
aJa/WlJYsLEyOxYuz8Glwba0cSO4XtS290DVhMTzLN7G/8suGo3wMivxkZO2www/
i5825pM0tPkq+FJCaNj8fmQSDS95BTfN3Mv4QAPV3IX546BVjfk8kFxqvSf6fjgb
LV2G02ZadJ644NrEm8x+eBd22ycBu8265QPFPSc56C47hGZOZMcuODNmBKeBxQSp
58qsQWR02dvbMTMR6leGSK6s2/Jo7XL0W+aieMlFKiqdB5iTdPGwhRzpXHNGtlru
5E/3O/Oy2AdJyw1ovAc6rO3pGyInAIFJI4eo52uF9xzlxx6MX64FuN7zNtMng9Gu
P9TFSZCnsVZUi5jGgQxqNRJCyXc7NxTCIveRBQXWBtPyLVvg8LWFEUgPE7drhMRc
dqbHgJ+SvYP+JG+/2LHGsfnTOfKYxRJkgwwgZs1U+J5Xzj6RNkl0A9w+r+93fmzt
ZfNA5ppJXd2ONgpihKbUm4m4nugDwYkK074oQSOvgIkAGPuQSPuIRbi1nQSWWkoq
1Do/jBlju6F2YfaW9pJ7gYR52IHiwfw0/+vtB5UgQvwdzJ9xaj9QD1Hwh3MzDQ/D
a17khJ1J7MGm7LAO/oxUZpF7qf0VviUiUR/BOjULcpRuWApaXY6v7YNJGZ9x7Uct
AhiKIIG9pGyUe9voGDS+JAdS104Pz/JBfk1moRrv4WMNW0NiktqAFq8Qg65CrTAP
Nut2qEINi9DdKCqWi96+iLQPy8bXztK0pzSe29AKM8Kv0Of1nqncUCdjtZ2XY6e2
lTrQaoh2ZvgIRPhbrVNoNzl5oRxZoBCTPsFZZrQqF9BGU5clXrt8RYFfvbS2Dod+
EwFfZNg7xYWvfk0TWv+Nm7jTGIwYB7hkH4K4YPCCW84HohkwKNSSnFmXtnnPE288
ved5AiSogVxsefTajnDaEZs3lVEyRECuAUlkthoHdMXk/fbn+4omCdg9utQARu4P
AYNScckIsC1JEDLJfGrLPO4eKsTqTicqQcLymRmUqb+xJ/yIAY+H1dxJzM8DHVop
gTOQbu5Wn167rtQTe+rOaaUIOcoX/IYudeQIPheUhfZ3nAETn5s8URzPtMCjJYvK
BCMJ+JiFqQFfvMVZhBUfmqRXuKsh48OLzVoyrP4PpDjj0oRZkBQOwXT4MrgCVhW/
Oq+ZITXjQkGjT0OX8kS5PYkV+WwoYbhh/r66MTTwPM5HyHDV+66+n7ae/rSYrmeO
xvILpkhRj5RshhPeSVReu0Z6j2kUiDO6N/AQS52n8O20NT30i8vYLQ5WNHxzIvfg
BtvAsxZ8kmcBHHemAg7LHTN8NCTojCc1HGqFnUDZKw4DOA/vAzCTtiMKQPxz8BoJ
qVb2CWzk7/xlgmOF5lrh2fSiNsCwe+uw+RDYChOAyyExxjTPM5pt5z991xdhbg32
5R2YwCgcW4M6fK5Ei1g/U+Z3RCHbT0r/lCBGU1oSze5B1VOpOG7wOICwFVws3MTY
Dj+w1qhzEQxfkZYjwsHTH9mJxJZDXYtBN5iirkzeW/tY698PMHi64pMUsKxJXmAL
I/5D3A+fuvtYkNPzwAH1f1uaGsqwzYJMuVfuuOiWnXJGnrefihyokxQEalCXbX2e
DWCmItULxZydsGpVLaAAAduzs6G4cHGDzcijtfFljaLL1JWR7zySIP/JPzaQ7g92
dqWizzMlbAJTgAWJShiUVUXYU9/GYw9EZp5DlcDSuai3bEnWvLQhFi3nnURC72JF
2DGOTRKmRsnoLnL81bgUUSwNIl/HRiP21LFbRMblvfx2MUlh6M0cd1EsgtPZhGxQ
9ptFiHjKxfx+Gap14yXBj51BcHooO5hOiQw01KgV5oEtdlhq7CNBE56devfjsXUg
CK+kPrYW05ORPh12DQhX97/8p2wARyG/aNQCRr644QCwHxVrsbL321w1gjqgtnuO
q4IroVcY56gaT4667LyMqblHcJpalXf0PCqh4eIyW0jRWxvWdwuVjQ/DpTOpOGLh
cxRH4gG86gjlgVVnnNtFHFVw9V5qQBeZi4AqgU7RLkngLw8ArHFIBe2NlpLVGu0q
WMUe7znsLRw+FRc6aYlkBE7mpVGNz1lQXc+0ZvgsdrLnn9AJR7fIznj+vSiHO379
KLDaXquDgyQWdBvUsKpgRTFwjN74pid4FUVq3cBmmxrfc5xVhXDQlSQns8L5yFsB
+uoa9Ee24HqsU+8Nb6s1m3b+M7sLtOeMTXdR0VK6VPM45Rh+2Uzx+aVDeCrBRLe0
2yUMfuwIQ6YK/EHrv3jD+IQt6HwSmV93hcmxq57iiiW6+7udguKBAgld1kab/gOd
ElKGkRpk6idGRI/nspFpNmUsZaDKg78l/DgSOV12GQmDYjSJ4zjxvHf73BLPFPhs
zP9D5ODROjzxYOCJRGiv84rU5spZsl+LXHlcT3jy/sKykqwRapzKaBHZn4vL5qV0
n5NGI3zZLKR6RtP+K3CstkZG2JKPFKognZocThlYhNpj5ZIU54aXRBpmvgWkoG6F
d9FX/Z1RADi1fRf37h02SASKHEZlys6YSwOYjswPTpdSDJBVkqa0uJ0oF9cCS++R
wrKC0tDukZYF42d0AdVHAcAm7ajcm2K16bi5VNLi1bDhTmGErNdwbe5HUvSmifUb
zXe7oax9yOGKExs0UaxQRSHPA6laSZkKv6EsKQHk1aRnHvDYsWFgQnkKTbErYDZA
GNzQmoPrybSVTg/NirFCmBngDefKfqTJm+WXP8pu32rBm2m7xM301ilJw+L5hPNi
IysaUAK5M3kKJ3930uplPbV/Rx3gWbegyQ4uaRWc0FEko+VWJ0qSwt0NvQUjzces
5WYQekq3WQceYDtCm9OWDy36g2kml/hNsmBRj3iBCVgGOXms102g7+rzt6a12OZ6
bbckF5qWO0m1E9rTt0SfgDYwFtCl992wngtxfzzVk90KCGetfwtkbhhk9nRwzvqo
mz8AI6tRJ77cZf5QY+aw1Is9fxOLHUsegK6MfybQWSAO1WM+6+5mQnh80HX8lpmk
nT0nXrUzPV0vbUjqDgQp9mGIymPNMiNfkb/uRoi+oXojtyC84YqTBJIT/abg/n7H
rvaxt5echFmSVC6FAzezMOIDvOJKVfaGSYlXjjP8qsSynwvAmpLrnYiOpoqHgsk8
t2C9owh5lMGkYwavMwd19lahHUJ73ejPgyL586PxzCXFzU2Gq3Tk04Ne/kpNuj00
m0JbcbUSCp92kN77NK8xiu7x5sCAIYrVzOeQLE+GrEmWTuROuB/HMx50vsNYB2kt
Wm2kpsNnF3JpCv+1UIucw6yAkDwvY0VLfCMzG4oNF8L0Y8R70c2wY1yMkcMFnZU7
yYk5ptMGZY+k/vlCP0DLSsZaLsdYBZ1hzBYqRYC6DLHdzh4BJ8bgtsQGVWNM3Hjd
TEbG7TTBw+B/6WFcuaACt0nwhuv/gMK2budDfULxNZgCd44Pz4nIyOk3La8lqhmc
5/gFCCDHHBTFhQUub+xBzBdtiYkJsEDZYhKIjvv+IT44ZlXzuFoetpnzazPe+RVR
hsg067vE73OnZ8BX7e16DzFAIllzKv4LGCBv6T7ZHHPpPm9Pa9HtHq0QutS3V5Te
17hmotZMniOKgJOuWlItkVCL+ccqsAXKJEwhnDJOaPaK8Bt+yQWMZZTxtuCxkIx4
SdlsNU+gridHIF/PgxITK4xetxoqY9kBNUgo/4dZhNsuYqb4vBNq4IqTLhQCvnJ0
Ubqt9/5dQfAqT2zJ64kPbLTQZSUSXN0EyBRPcjYudFMlIKrp1I4YULmLtjNskm83
ApDSaoXUCkK2EsL17GJICMldaKgfvtCr3BtA3tJgLz+AMU/WHoSTg3vPwf8T9nIf
p57cWLY9imy9jPCuL5/ifTfYgo9tmZGZvGS4rwWI4eH6eEqZkBsMck3qi/llN4VR
s2vWZAARfo/SGBrkJ0f0Yr5zRNOPEPYt1SR6O8XxpQ3xfv6hZIwaoSYUx2kSBeyJ
XB7V5oF243je+Hl9bGOePemM65JBDJZg1tVP5se4+ps5OMxbj08QGKAmFqBBaD/f
9KFr8PZWzvUC7Ugv1FJWN04GUI5MF3dpNdt+v9mjkz/xW3Z1DmzQw2nR7Pw4YeeK
Ph4fj9X4/PV21YHhytjXAdfUzgB5UjE97a3HDTrS7EOhCAbhlqAcA6lLUi7Si8M3
cp4Ung69mvdWG88wZ4JBHDihldT3QIE17cjbxzeOV/D8mGc2ZhqRF+eWbXd/K1As
ipRr7RbCGKCKnCm5ok0mATPF6staRVhn6lI1C6fVNWXaRmAMuHFMYVYY/t/HsBLq
z6LDROAifZBC1cM4MZorLgfCwXT+Y7b7+E3JxW7gh7er01fFpWDysqDMXislv97a
ym9iGwo9/SuiQYFP05dRJ41jarB+fFeiy8BHKvZA3C6A/LI+XMVYD1YzH1TOmfPB
0/9T2p1qoPkheS2slHqU0g4l5/IMolzD5loSSoTO0aD9UKENpg0z+IL3STmo/DED
LZUEtmpW0zyqHJnFEQWXz38JNVZG7Ve65+xv7r51BFc0jzoRda8k5XZPWjrg2xnB
JP+fG3AbB/xUbyVmfEIEnZb4G5YU9zGMNsd1PEfS1OoIyC74LQp+VEzlw9XzaaWx
ZzkXSyVgVhRFqPu+i55aBXAQQ6HJXcp14vNwS7lRJhwgmdpknGJOjbaJbEhk+hHz
Lt3Tip35KRjBBMxqFpOtZciFuHQre87nOJK72S6+daURyRHJH2NL1VUwwlzN//Vl
gq32EvocsnCbG4Ixxjm48PJe4rWOGznzhXDL8OhSwm7HQ0Gycca8eOsYAPVR2yjp
NvxpetXXIJlFmbf00zXT8j0GutUkslXS3WBJg2AibMtUtKIThfO7b05PHsapDhJz
n9r3Awi/En6w8hboHWRRWNURkxD8eyGU7AQTTEs5hvF5EaCE3IG2swwfS1r7EWB9
rXXo9WRz4v+xWsUE0Lr/ISFTzCGMHbuzj3sZihd8PXdN+XRg6Yjt/8/eDYr5cnIb
DbUgnDK2dkm96lKcfL0yvcw/JvCKZogbXj7Da/4/XkTEkYQWMGhgiQHLvt72lE9J
XaV+VqKqQgAhbgta5TCVJCFJrt/wf1/Hs+T1XtnyC2uIG6R6RKe+YjLlcc25O9bw
y19y22C2hTo3x2GcnzasJ5gaPv1bFJwPSEdkzp/iLUfXuSzaRjX/IArGnIEz6rNr
AWE6USMv6Q2tQuLPO9+NZU+2ZxB/woQtHz6V5E9lOtD0v99Ps2GBOYWJcPiz/Rb+
oj1Ve0F9kqNrKaf40N+VSnCzslxl/MD8cqBnpllUhHu6RwxDIcXYKMMo0U5YeNHn
jm43QLkYyhhQwD3X0xk0AcXJO5lwmhJFjRzRWWFlzwl5XZ8JAnRDXDUNRaAW4K/8
kCYBstEA75IeKF9MTIJPLcFdN5ubBnPvnStkhhm+TyY7fxH1OZrEEEX9a6HX3LCc
OtmuIOxCh32MG0G9RwMpD3ltwj+9coF11Vt720RDBDhW8/G9M6qzv2FbQRAe6x7j
4N3Fd8GrnAgKzGoUWFDPmYe3JmkaZlblHuuLYgEzdL33kTCEd0pkDRQf0YhOc5Tb
BhOeDvOzScBOBY+InWNB+rLm7KrHKfeDLlaXAWc9PkvdTLgVhBHZwntAs1Hvucqr
PqinPY6+dqw7OTEgSIbt3Xeg26dvC0o9P51vIy0o7pyXGMRWhagRL6kNeFqKnz5h
UogHrM84J/bwYmoQAMrk4ioA8WaXY38Cs8qI3c6Qpypa52XJDU7ZGggVi08SjjuV
b9fo6yw9j1hooOS9K0HlWCMvs3PSxtIoxZbUrdVQL4eqYjze1QdfnyfDHgkxitc5
rtqBK0r+dzormjIXuoqd9eU3t65aBnEu8AU7rB1jCpX3+V2YV1Tt/JxlIiBWS1fb
dUXPTpeBxH9YrYi4nzoHPqSUKqwePlhuS1ghoLDEh+4AJSsPcnT5R65c+/HIcQn2
bhw8xMtZyr7/WtLDGcs/+URWSiMVt0JHWvKFnGxqtMM1fPw5zzIZA/YcFk0lxqOy
okNCui9Doe07WbRijXatvDZwybWXHuhhIRXyS3cWRXNZAulb+Y1Y1rgeGbH635h+
jd9b21U9QQidQEojFrgS6SZqjvGnlSR/z05gMnZkbclYOQ5UFIfl9yYLMd7dwj1j
B9cgdVkWsyv9Lw/rVujczdZFRPnoof5fK/sW4BnvIDGQbAgSjq3km5iQCdH9Z6ut
ut4X3xCCdvHCaD890nUdbu7v79Ea6pOPBz6muiJ8QObtun27mOq0iCtONkHtnZcT
heJ+vnJSU+oViuEy1STi8x3hDktHHVgs65Kc241N5XB9Rvzb8DUsUz3oGNmBXktS
OfScUomNoz0kjGM8D1Txn4QXl3JZuO9DPBHpY4DbYD/5Qxaq/ynTlhzdN1b4LLSp
1czHULOaTkNOvoWyTSAnji89QBnEelN7BdhWD9ymzWfnurlCgNsZFJLLVR9beNqa
BdiuiI9wTW/82OnklY6UTQ0fNEq9+B6j7OBpFy8Z0LUmOVD0KYPCXwh4jfVVDJz1
Pm43idSrO6dPARbr4oSZ49MBiqDnQAv7j6DucTpPAaHI+74zrz8s6QAAvbjC45gp
W1Ir68Xd4WAsURsicikY2jxa+CkDZyCUzMRjNXjlQSOE3hyjX8TaK2fbtIpy+ZKk
2avG1Ggb3IsxmHtSiAzMnM5EiL6RgVDcjdzXVUYSNPWhSUz1pM0d76t1oJGYZlTB
JmA+L4KeuZoxTfDQ14D5ZCiHILEP86RWAlLC5l9o2oe6AxjmOLJZMxRAEAnDftig
AcFppv+FHofnC5RpGVulcs7hP4/S+TY/vSpM2WzyVM5/QVePzBhcNTEIILU6lkQE
Hzqsf33F9UYLaVMr24L8S21fseslMztj1rAHT1yaR8OXO2ygbqDEd2GNNRR+vZyj
2HXRTdanlr1jWu69F0QAtiRK7bfrR9ByNlhXJQjDom6CNfxK/L71YA25V3cLzkG+
s4xeKICIpux6MOWwc7KwQlcekJdnZuiZS+CBdI82jZVGNXu3lcw1oC5qqv0Bfjun
xiXdu0RAA66NeoKD43LDP41f1V2XF+eCLJE0bcddPOfx9gtkJIWmrXER3XwjX+aJ
zKsbele7jFA9LHgHqnlstL801i4xhMTmVobZ2SH30L6XI6rJwRKnTnYspUPCbBqZ
vhSqGkUxkUSXoCu8J/Yq+O238bfE37pbZqeMmOw3WSWVm595dC3uThglDcWXXyGa
1x1Znfk75df+U51AjXSjza0HSLQPoPBOaoNuQyJTj5Pvz+X4r2EcEk54PezZHwun
52PvQBepb15AsJXw8S7ChJkHPcceiR0KAgcuKPIS+o6Ajws37PHaLKzUJDSD9iY2
nHd1APxKD7j1kyIas8asBOIKpKoQy36yeX5vWnKBDaqOYXmzYN8dtDEOt9UoZ9oZ
CVoWEeyworuHvRjf79qwJjxTEtXqgLOcbmbKHr4f7xO6D+8uU0MNkPV9z0XVlszM
cRPzx76gCp9IMeUCusADEjMZ9acq1/77UD1OWuN2pvSpc8b5BKnMzRq2NBImApG8
2PY3rtO1uOBoxkmhgviYWZ/guY/0Q0M/WACI2zLP+qvmIkkFF8LisoH4FSHOBeZa
YvVvP+j3FHxreDgZ/50C3rGQJcq3pEfZ35KhNd3T/1I/wD10SuVQEyHabT48/dID
LSJ+puyqrWHsTrvxa1tqIGFnrm8KQaB+NoD2txp3t2Tz4pqtmAc2JusaSocgDpIf
Cm6jd6xykToK3zWRy9jGxwOWu89DTMQ6Uf+1AksekQbBrKB5Zxlq10qVdy2Pgc/b
+B/ByMvR9QkcUhKX9IXuBF34FGq+zTMsDdug1z1HntCSMjPDPj0GQmv9g8pJZpen
1/2qi06jC7RzHYIJFgrJsqbPxpZeAObl7CsMmA75CLixxOXEMEPAAE3pNV/milUQ
umHC7mLY9O9IeT9N+WfAHIHI/ogeP42cfmFtUF6tKEhekhVtx/8D04v+QBIrQfLW
03K3M6D3Xyja2xmWxIt/tJM13pKgpoccrlVCw7XvGjsjnhL7l0Ywhv2etTvTNSMr
fgB8ejKpzSUtR2+SxLUDt0I6aOqCJEbnyppY7WOzfW1aJ4yHN/JRdn7aqUUFCE6d
7Wd9hQKVSSsWoMX9sB85kA==
`pragma protect end_protected
