// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i6dd6N0BEvz2vqrUMxOVR2dHBJJVGT03rKZMYnOywyB4RFWoCxajefkutlMzAEqN
v5PKq4VH5ujdOL0qXTxJraVDnNVIDDKwJqKu/Qf7QSaU4YPYaAyYDiR0h6ASYawd
fBOtdOUEHGSbiDW8zq0nbp7/fEFHqF3CJZaWsfEA/h0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2240)
zwguoxc2893JmeHUCvqs61xbQp7ebeev+X8iDJA9wczZJhwadpS9cE2rLo0EbqjT
mybI3/he7oGN75g8nnilXaLIUcnZlkC6I6n6spksgnnRHs2jho9BhrEnLE/6dweS
BSmfzRlRTmbOOuraCU7dOpFOrKVsPKsCr4pIrwBF5Kr5oTxRXRYtmye65VwxcAlj
8J5yw+g2tLe4FuK4+nD0ZRAmRZAjw5Dm1CXeO1zn379IByhX1TnHurGUPhs4jL+Z
9qxg9m9fwFrJFCgpMREJb5CZuxcnBRaYl2jBJfULwbS1TifnNPNGRrU0Cbn1yHj+
7jZOebZfP8Ch865ODJAmt3CopFN8p/Pl2KBRAml4flDoAF2mEZe1oH7lmcDXNxr8
X7WtX1LGvsbgjHANyuo2qdqShX5htN4Q5CDOEgMZa7sSLjKS0eASPnyWd4g/cQ8S
8x7s8YiWRipKzgQQR/EixaxHgBVBSEPRqvtxmHNEbGGJLeQBF+pixyjTimA06ex/
is8kewIaGYyMTz9gRrvWRTX0nRMVDo1CuiZ1pSBO81e9FdjCPD6bUFhY5VHf3isv
H1eBI95FNPYokDomzJ24z7yXt1IfJxLq3btPxOHPSkT6f9UWzRDHDBBGOCf3DGde
p+uiJG/R8TTx2vRp6qs1MWvwJikNXn1tjh83nGpDs9614Thivl1hG0RrAyHGCZYP
gwYghNbae9zBSQRmIhEBJPsCTe70pJ4wUi5J0zOKch1tRKZqoLQjbQMVO1g4Bup+
q6vfZDnOL3PTlS5Pp1zPK0+2HsnzudNElmN4WEtJiPwUW/6CtDUuEZdWiUUmmrZ2
j0m2LrNiOA4IEHXyYCvlzBDoy6KTB8dRrYmHgTmkDFY7ZFMypEtg3mafy5Uoq5PL
k3cHf6helGhc73/P+jPiYS0SvFaVkJFx3aJq2kQDm0NkF39tRGIQ5301mRDzQDBE
7wgZ1+awOkRiV1OewV6lg+U3FMPjE5pvtvwGFaySVNGRx95iNc4aWepWGIxegqrR
QMr3g4EETia2x3/g8fYfBDLDnsIOypOMvQP+QPaZQxwvx01wadn3gXuQie6B7kap
itUu6vbRwNrW6pw/Y74HVSJm1ZETgHAOUg4KUKwiPrkiOgN6kLXEAV6fTmsLQXGC
Th0gwx2cyuLC7L99ul52S6QtV6EkOKZhFKvNAxpLAvPOqCA2p/JXADuA52lt6VXE
GYCk2ddpnS7RJrgzEBBCOlQMco+G/1zfbxgzIQBdozPdW5XnMKlalU+dHo157WX1
W7x6ZQ6GR9SvZQh+XvfC95YlSZasZbfS5dDla1AYx4idQN8yAULJ3TAukAiSDtqr
lf1+AXe6xrbTtgqYvI3ySWVF5OWW5ZWG5BBvhXpa0NjWm4jf2oZN5Lin2oDemT7d
psFbmmwxXu0QeZQH2+k5VrxE6zI0iC9bb0YWIdOqfXFaXI90E7A9TaMMtjm/Uq4R
r3Hffa14UxM1q+WcU+mN3FKKKAld9IV3zOfm+VcJnK5vpy+I5yvzD/7Afo04LK9t
nYGUn5Eu3KsIRboLsDZIdXTT4HdAjpll3ZR+CKJ6yNwjaHprzmS928EgklXx3TmJ
r3Am9acGMeGIEm900hhii/b7nAL27/3ZU1zrc6v25JFkTyUKo3tSrmbljCsAQ+l7
H+wgvSU6hLbtvlYiz4LeNESb3MJe9vqm+7KOKjRwtXRp12xgldIC1JsAVmA6k9hj
J64HyFuQKdMGEE2tiikF9OJrAhuSIC1unGdFdtxoQiPvhm5RO2YjyOm4YQd+SPWL
I6Qh1Ty4rs/67t32vYuHJSxJkXN1R2n/zt3z3oJCHe1tWqiuMgjA0b33n+d8sjgD
ONE7T0IAIngHkZhnOQqVY+RlS6twveV/+u9+TgeRzfJl8lKj30PIlZV77e6CEnHj
MoJ/4H0tvD9L72P3DyLbf+zSqqmnS5sbvhRSyhJrllwLJ8wGTbMzeS9hX2hIHHY7
6E8VOljju6FiAH3jNTFNZOTmi1K2Cn7M95LUe/YjbaeCOgbf+DAOCWhswTCaaB/y
3WyluP/0WvcOgRO9a4iJhRsdIEBi7266K5bj7B5LhHNS5C0k0jj/ZmDRS9HudXJW
QEQr0j/vAUledxlcZwHFibkDGa5zTcRj5AUnT8bzHyXz0XPpW7ucXmSNpFKyZuRR
rJ4bMJEGBZi8itIWe7qlbSrt9C0m94SlIK3wqqfJKEe2czqU3nS3ed30NdqdYvP0
4rQmQCMVghck5YqkwGiiPI8v2CxtUHAmb4qK0LbW/mxOjDidZJEEW7phB/pmMxGN
5DTwMbtZ6W+9PjZlXVixbOF23WL/2V8YRJjIyBfG5aAXTQw1x6ZljNEPuqxyEkVd
05vodJWPoFv4H8xFybsRYV2ZoIQoBEOdiSntEvDIhBLvFk19X5iO4QvJJx9wKVnv
QhwHIdbTVH766Uxz7KeealLmBc97nb3Q7HYO5cXaHGFQ2cgZf4/5PLXMLNA9Lqs4
i3BNA6y0Ez5g7D53dBjTt0m/3em/kdv3xisss+xTwNpNCc50F3ofdt0wvU6rcWS1
LivMpO4ctju4BFVhhDFl1edgZop/Pp5XgDGaFeCUUFfFCLxW8lXEj3KgoA5JW4Ho
oYtigs0kZEsmDkSy78b25Qa+CtGWPHHu3uQYsfj//Sxa05dNrSiS0LOlZ2Ya0GKJ
MYCurCoSsohSiB6tXVmDciwrO8ZtQxx030+0BNE+jZ9fnVN2ZCNLya2Fg1ETySym
ENbC0IUVpSMcqAomDaSSVVJlYGYTUbEHoYWvxQ5aV4IzFqR6J12UmAs6xAdjTgJI
21oEfWyvUVhtCSeUgf4Sono4M7C+zrJihdT+zxyBcWDm0mKOOdWg3slIou9XWPAr
V0z7KGD45e+Cx/kgkHxyxvHZtO1/oILyTBdSz4UEQlLcXCku5VzKoG1EA58J5/iy
PV9Qn3mVDVNlFpczKmSlJyx6euO3mtk80hQ1RJ+9W2g=
`pragma protect end_protected
