// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:51 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Du9Od8twWUCxCF/ttCxZ5EntfBjWYC+o6vJDAbicbprXeyBjo21bR8mjR2IFTm/y
/tSrCuQviVFeJ2ewOx9xKb4V50fgscegRTVkYcpIUFRhFbkYb7fUuE0mPKuTreWp
j36AwnpCXqDuvnI+oCGLtPohaQuy0AP2g+4B95vwTlY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27680)
qpV/dE7OW4Ruz95L5XOV8oq46J4//sinaYxYMa5r3U1FEseFtt9aufCGT5WTW0LY
p1bCQLxBiLiPeqdAbDdfMLaQDwrqcXYgqLn4awnbjKEdziqUQDnSTuGiyKBB+klY
5AN3m0gG147JFbBoP56H9LiUt0YG76aphO7wlizs7rDExBs5WiUvUNOealrY5c41
8f8CwWKkp4Q5G5GTEDFiex75RZ0shFesGq+MxSHgSZBT8sKChz03MfWKj9hHlfIK
5G26Dag3fDWnBvW6oXGucnjelpeABNZzaLIr/Uk0o9ZCJJsavqQZJ/D5MTdlAhj2
+fiHsx5NUm0ScGUv1Wm8BbI8rFXvOtycv7If0kNHzJ1Mc/ArOChE5mVLTdGbOxMa
UTxDzdLp69Wlvimvsz3MOJT8vSsYvYjddc04RsYnoEeGabDyhFsqTaG/51qi833s
aNjMCXYg10ec+y9qxFzeDyhO0vg2IXbAmp0zBL61STQQJf5qIJGQ9rxms3nqeTOZ
BwPOlpSQU5FmlFGGwPN4uZQKOL1WNpoSyuATYlHmbKiOJbIomnKoirJcN6j9meOG
3ad1prue/yXEThelcYxrTXeGXym5yi9isevILKncPcC774ojpHIqtgfS7NAjTe7P
qwtoR7V2Ul9fh3/VDsAa01PGU0nw7qXaDH1dySqKcPL5F5qlR9fObr5ovejO+WGk
qvxSMQIXfcZ+hIWv2FKOKtzrQLUH/kB5ItDuYFUM74UhjXmi1+lvUP5mXAULEBqz
AYpVKopzhj+L760cE1FByGCt/Z82ykt1J//fCXE5gkzLibmb7xm1CNPYrXJ89+PC
emh4Aw3mXh8vEiH2Oi9CQd8M4Sw2mi7XNvC5mALq06Wx/jNlALSA2gSatCTr/E+a
beoBHBPrBf4kERaCWV13Fk1ni2iLzOlYlT5gi2JkUJJU4bSAUswkFsXm1W4QtVzy
1ACMf+lwgOXzBEiGqEoFdS+AgnAXtAmhBJFOCX+68jxcn7Pi2RuCk4se2zsz45rz
BxqtGYGv8dT+bDe5/u9DsLBNuT5fu2yVMAxSGPVvJbQPfYAs34zm4iVHwyf4dVFl
FeQHO9SPmuyBIqQyGafgIjLDHrBQqi217TbWkwsOkIUGMfR4LCW5GHhoc35rKYqZ
mSxMej58SjI/GQB5AqubHOLPZ0N3kGam/YECeb1IPFdB3dWBNju8JeuGedadhxOK
Vf1zDxJ9tbklTRQ42FL56Yx9uhNT5j6gCaEUe6YtHnLC8CTsVBsXJ09YgVKgeAac
4exISnAS1ZSikhenHZvXfulW21wLM2aiTmowHTbsJnpxcaJLIK1cHevWT07u+O/2
pzYIIE0Hl4lPbNpcY/+eT3hOb0gqt+CFU068SDX+F+l3kagpwWI/TQjaRaEfWQpQ
MIN9rvNyVeBpJFLEp04B3tHxC8SCM9AoYtZd/CXKfLugmW+BBFgfTvf+gjNypYD5
IGqZ+NWu69/k5UQaJRfEXWHk0RV49rPCQperDTRClW1G601qxKH32+xKTwWh+MP2
2pNE/VlcfoBsz7LRwiqRTTOuLAGp26atN1Or8GbWCL+uEkfQzV/w6KfORzRUGDDz
PNE4YZzkoquidofY1ZHFxsb+x2ijOO42Rbc1ZhpB7Vv7LQAVsxjWgh0D4boJEThm
tUcUY1LY+nrzbDo6lALtCU7u9Hjq6WEfXxI1jZEcg7127fyG7xo5rqzMS0JOe0Fz
0cl1xMpTXyAIrUK0LW8LnAF5zgRPVCf4XvMMZS4r6LgGqDDsS4vQNvTG2vEcnTmA
IhGQq1a58Dm5hF3DikNn7V7mPbmwlVCK914deA6Fl5XLnCt1lrYYDRsgCnsL6VIy
UwOsO4Ay4SSUzY8WWQ0ou7+Hw00v8xavsj+fUE1KEjrCgBvyMT097pLWPm/w5YCI
SQSBW7/eSBCb5bY282LudyjmZuGAoFVLb/gP9tlPRZi0DYzN63ZjR4+QONGgi4Is
C4rt6Bz2sSrSGxgVAS2RvFL+q5OgRszXgz2euHB4cT3sI9jdnYf+HvQ5Dorf9I9N
G8zN0CELYRWxititUv4/IMqOydOFeYJzHE/uLnZqsAODAU2l9lnAYgpHe6f54ohG
1FQWvwBTEkz/m7H5PGk1RWeWrHc4XWyRpovyyj4T12i4SonhnWq5kOTLniWNnKZk
N2W9qXrtWyQu6EgS1xM2WLvMdhqEL9Vy4JDHyuTLuk1pmbLOqdNN+kjdKI9wZOe4
Aum3xFkD4DgijFLN3a8x0vQVshwI/CW0f9vgEbdP+A9MjueagwjSTZd92LT3wsG7
g+Bl5qOs25VRjTd9NOFKiIdetg/piN10Bb/HBFiDVl9NhcpLy7ARz8mGvqK+Xnil
dhBWyH9eJ29BcDJjNrX36JBYV7JdSAaSgoIcJS2bQJpK9cLq0tX78vOYuhu0qrp7
ZZcaE+WGHTJr3K1MlkDH2hu9uAoOusElQxK7Y0CtuBLNlhL6m4Xf2KMtTMdcrKfs
FvGSp1okZWQqxksVaK4qb9mEnVXU8zTmxcgGB3tW1XyGPKKVZvjJZ4PvHy4WpuJ7
UXO+SsisXhtMUdnmEdAfoHmIoGC9IBgSvmxCGUJ/gRvn+RXawthNtBnVWJZeXvdB
zpVvEQ22uFw4MWCIr44Pf0OrPh2RvwrzCF5VejYrqf+bJhLF7aq1lBlLhYY/meXS
m1mOOdrFCZtlsgomUWQ/dzRNxWjK+ONoUgw65WeKzeSyvFzVmMaSDJP52hqMsqvv
BWG4oiBIp2Cdc1Oqi4/w+imhbdwnO5n77s7+Qo6OIPWTg5ymWQFTYnS4yihCJTyr
eywxlWJmMFMr/GehgNtoKJImoWtK3SOYOMUXlK0AMrcUHpc1NV3tResIrD10eV9d
fEV7EbZaE+vb4tjmko1vL6C+9jHRP2EObaCKneVmuYKDzxPAxP6Tqf7aVihKNhof
rz4uFvDpmK6PULNskEXWP76sDodCY1ux2ZkVo/wfLmFndNtjuLOoIQ8DwreEu+4u
r/Y+YzF/Pw8ZxGaGu6L0GM/rEhWFUjT1Z8HmVpdj4ZEtUuNBw/TQw4SY7k8Vc3Te
WTWOPp7kzETyOwwgils2REJPUv2xygvlZw+kIIlrVLso3Nmuo7kkQ8SjLZeIg+eH
K4mikXQXN+agXjhufmKhXf/14zfV2ygAwHQFvvATIlUv4Er/zDwebJQoyxDYoc8e
t7WGAT7s9ozn5i3rMjrivxWPV6cbQWk6aiFvBddN1Y0dZ6K3jCAhICXELjwDenUd
uLao2sLJTdWWqql8w8wf5rMbWettHnOw4GD9iaBI8AurgM5ZmrMLJpIyu0ejoA7A
D3OEu+NcNEARYjtk94ZswjQ5glEs/vseEqd58uQFrFSluZDYNimnzfjjMp7+xQ4R
EAyzwN16WhX/qMphPf0tLOhC6h1AUmrNIqmfCCj+KFzx0yd1Zwl0tM1H3QhNJKKa
jlNpoIxnefIH6KgLwSw6MTHfxgXe0PqKGL6oFwG0ys2YFDS5KQ0PrSGwZpJNOBTh
MXKGP80aXhO6eu+28icwQkUosK0aBbIfi5lAImWY3gZPmNB5nBD9UGoOlj8kY4Dv
v6sOQz3XSNcR9S+QnSFq+wUmz10BEgEFtpiUTjWm9ox2U69GMDArVAej7QxABzEg
b39JPISk2yIyelZzUHYG7QzezAwbQ+JOvlpQqPnXuh+OELo8t2k7gbRaTYbjeHwo
GhRvpXyBxubFJiQqpHoi0R1UuVYnygh7fXdrv3MrxOEozBB4Ko3M935RJVwgCXic
1+De4JwapluW23TYdC5osNyRghRFuvQNMSAd3tqG31RnrRXyakAKOEOAnQenLDkH
c47tMkurR3+aB7YR38OBN5ROzVMyJdeDgingb5/FJ/ga6jW0XTtqqmjv0mMX09ma
D+0xeOsOvVBJYOznW+Hu38aU9RUPZZaUDo1P4E8VZ3K1mg9dIGvWSzNKU3lSyyrk
ti7Sj2hYOpnW+3zKcRx+bxIuDPDVcpSZI4ztEsr0NYQitQq6uPr5MIbe3NyF2W3l
VsmEFSEY2vPPX/tZcnCacet+wEhaoXqsBrYhn9Bhx5HCYZiMfUxxgmQTVeVKUL0E
3jE/TTzMVCo1nnhbFUvMs/NDNY7k+go3XLqvmkllRrwMmFrYCnfpJvbpPn5exb5Y
AdIND744hbGmZfKDKHFN24CAGwETkTZ8Ji2KVj0cWe5AJfFYSwoG9QIxLj7jp9je
jNRaJiAZmTx8KaK3FIoJOxbzYx8A8JJNMmF9HyzxHYK2Kz2l0EktW6+IlbnACvvj
vp2C8nQxLLcsyqHkTPhVwS2Ruxb9zIUfUFg+tKeZnDvIQiGJh+SIHAe9gzT5lGFh
yw/1CVdH2qvvDldazcspPh974+gRwnZ1BuyBUNXBvAdFNBG1MpuCp1Fv+AEIwwuy
Lc4xIP1ZcjfkeznETLO/5jGbKtNRXDofSK/LHOJnJncNLG7aN+lZfiJIOb+ayiIM
w+9fuDGWVRCmoILiCQ5+hX3eD9OJa8r/HOXZ4Uky5e5YbakI7/FQdGqv1SBsAmHo
kEv3QDyFwNafpyHlhApiC/x79ZSr6ghLPzwX1EMKnMozubuhzZEL2uYSchSIfkjH
zTn8Wzxrl/edIb5uHxEVbNxWGJMkN1yeMcAG4ViugcpvQxBrZdoYMiAd7lpKfNbr
Hm4FWKisKWWWCiyVGqDbGWUMmYEh8VFDGRU9qAoSigLjGVMTG0cqxaoC7OR9i+wr
ioc4xra5fLx55Fb1ybPbH72F0mC6OB4/YxLqmTzUZTlPkFgcNHpEOj2+DQFWza/S
suNiCg3fBiFJ/ia2zSX9SeFNSHhgAnCtWuHV9xHrCqvfaq4hrNm0c8AZQ1tVCzWY
Inylye0vDD8+plExbpiaiQxNdQVQN8ztI7tfXacI8/1M2SnXWZ8UHbMfpvfoHWCc
MwPz0+TxHVdVB1COaLGxveVuDhFWV8cIBzMR1dFQ0v/m3WK7wqqIWERZj+SptF81
/LleEL/03ShQt/HX3UFYBmPeRM5wE8+Atn72ojE1scIDwyuUw6isIDGvMnc5bWtE
35Obo4KzE5gK5Bhdlr+d+2PlNdF3wCSgAM1hAqTvKT4ePaNG2I7KayFK2RuCMnxF
ECmsbUTe5km1kQd3U/tG0U6dlAbiJ5/NwKtGuiHHjg0rp4yY2IlM+odPI8cm3drF
connDNrOYVU/FNQ6PnK7eE3xm/+IvCuy7s+QxhDNohJgpeGX43RvBG4kHFJ5Wq+P
u2SfAlAr+kQJJteKwArpi/xaZkHMFpVcIhkPvR98NAS1dcI+H3BQiB6ekztSwoHa
99tI6yqUxec0pNt6tMLuSwS6Z72LODHnh0b0hdkKTCck2j+JrZ4uOb47QM6I82zW
Zu+JQt16kq1Rt4WngS5Pr4Vxq8nqHABz/SIc0QmVCsyB9fXlPXcHP4HeA2uPyAGr
eL7dDoXRRAXPAI23G33LB2rhNQPJ7uupHN+ydeIWa4mCeSp9qaDQdn8Frh8R5/3w
4OcKb362HT8hLGJQezGm++uuftxE2UxY50uBYabvpfSuxlwggQtd8BUcgdpiHGR5
73UeCfePOjPo3l7NuLzVqQC6D6oBl8XWcTg9/XduU/I0iOPOyrXWpGU3Heu3FyZa
ReE4i88Xqd30csbgGzjI6LpRMD6xdLStpsT3pDPTCj5AG+0QxGLNbKvGEJwKJ7sk
jASAOKBLY1nhaU9nSbR0ytqHtHODT6A4JPnpT96qEg5Kk4XNUu4HXsn3s+846RKD
PsHWKEfr08zGX2b3ezH2Bm3lkPHO1gVMMqHj5e7T92/kPuGCUGg0WreByXwZ8H7w
uhCIlRiP5tdryxmIhriLDEsfKl8vSh4Qx3190D7ioYl4q/DUF105y1ptuV+MXDUn
V3XDhGSG5yNwA2ajfqI/uIUW9gSgBn/LLTZd8bP7fs0Sah/l8rDAnp97ZI9wQrFw
RuGWKgLFlMeqxnu2AKgLiaWWcKWAYvYo8mzO9whJD6OnPRTjEOjWYoJC7N6BqHzt
rAMG7k24jvfOsO+6hR3MJv3ieNTbw2iWhT8etmuEeCm1HgMb6xc6+y+cWN7ZbFFq
wdyKXSKxRq/3+czdcXPKRqUQJEAfbL52g4pWoIcTU8QawtnPJkCslBaSAXTmLXad
IBH6UJbxU2vZTZmz3P9VT9C8YNPR7xkWxcmXFd+KXsstROvMxOSBVh1C38EP94HI
fhbN7lxKmqU5NM/396hVAXyQQa+mCM9jutHPT0Sdc69SGY/4vrTdWUWOOCB+47wf
BfpaBVr8C8+BEYJrn2j6xHWWuwKrgxapOQCpT3E/XFJX5Flm0hn3mx5KNiTNnns4
Vl0/gaaHgAvEROZMk+RRZ8URzI1UVPZMEEzfKM6XCoOKwnTKHbFEPiBOT+8OCO7O
8JGlQRr+nbye8uHiUmwJXcw7f7nN280m9CpIOUdHOQSkgMjgjY8Qvd/nqsiFUzHc
Vtk7o2jO7I4VCusLw+oSyREYh7p7sfVSzW39KxPFfBE4uNisTR4VK/mQQQp233Rg
gh4BsixY0AJz6iRhlbwyJftVpqb70A4i+IKu/8Iab2RniQBCzmEZf/JvXt3jfHvh
sP911+XOAw9qCwReHiSPJ3B4g2Z00DrHgJw3vUqpHS3t6lN1ZhfVvc/9ETffeW+p
voNDk913zpm2DkLTm71xjAYG0XWYUvQ0Sp1Lz3jnTF2M+SrhfQJJyeueKCjst3gX
vUzy56KLIrJkkXoOmeHIgMs5kzeY9YslB4h6GDashHkq32Elkp81QnzM3HoCMKBp
IEJNxyeYP1JRyLnhmlAPoK9oGEl1b95vgI6qYeX4JpeNwlD0gW7L5KRlbNMnxBmv
pk/K7Rd7a4DELCwsB2jK5vVm4tsxeussgmaeTsBBXIQZ3mh6HXamQW3BOJl8ba7E
3WT+mC0GTKYWm1mHIybhS9kCEhNbEv92zyzLB7E0hWyKGLE+xwQ+DvfHpwhdeXrC
zP0zK2DGiTTwEJsPgMOsQQ6CZXCq6Mt1ABh5xCx7xoQDL1Lk4XBBBM/F/2XF/0VO
TSJZKhxpQQXbfBhxbqntwP+IFebWjOsRX8IYy8yKycRK54s7qg3xVSRWDs0nTwin
fNLy2f3TPGPG/D0Qz9RuASePViu+J8oPDjZT++iJnyIh++MXLjUj1fyveLsMFliR
9cDojyb8BjXGeT45i6u1AQAnGLkqc9QRCEuNfbUSJf+xeYPiJ2L7lfASrWEeQ9og
mx2y64Ub4/ciVIJmFasXzeZ4ZzqzxQV0dd6V6/gRRgks7n7H18HlGuLOfbR1QttV
NGPgGB2eu/0UPT8V6x7ZRbv4yupp07gOKFSxscePJrZMhD8ggXYKBe6N3hP+HZir
nw4ZmzrHiAuDXJP+iSzBBQ2TXhInI0hY//LsfgX2kr0PA/A2oQClSuoIaHmOVLOj
5iNQChv2KYrj+HkOnxjQBrO76tWSSVO90djotMGC69nLNu9PBq5CzDh2G60abvzz
ic9C+eyrVrxfmkzlIJREdrZhQk/oY7IGv62+uROyJqfiiHFGf5yPS5ERRFVBphUR
GFUajQ45L1L8OmD9zMGKiX7nKhDYyksOnhblrzLeRiYHMC9DqGLgl9ILagIBbLlz
GyyyiOwp5bspVUMUJbZyJSQgRDbpy9JeMEm+Omkf4IkWo8ypypgWZlBL5Xa21V7g
IRDduzHeba5jO8rAS5tbVcHAIlH1b7TIRFNntUrl/c22FoOVwY0/pwmO9kVEjXOQ
qFJsSQPvo14aw4g4Xar9qpC6b4Yw83V6a9QaRNIVMLsik5BDWMwdVjYtgcVWfrfO
KsAKGZ/9P1fa/5gMvCSU5eGl0C+ioOBNAI6GyYWK/KXafeHQGI+mJt/X9Y5frJTB
/l5Fhk2qDkPCdjT/vFFeek1vHvtstQeYSx0plYb/WfP+Dj8lPK+uF3XuiPJ8UXHW
YGD6wpA4jBHp1OTZ+OaSa20beaDYK6/lEbbn7BrOvl2fu0ElMyNTaCK07uqpbr1y
UMoj9YPBfVwxmYvFNM8ZBnkplTeejzIW8JiHgWje18i19yf2qITX0MaE+bjTk6jZ
3u4rNJ1VFoEccdAyo+Io4YBn1qatDLpzi4CQG0112iwwRfftHiFc4UdHa/Y5IgIl
tf7ac1cD2G7qmQt9WcUeDA/+7QJHsjmT5r209R3T8NuUf+uiYe70+L2QirgPfmLg
UysSRr63D64LRaXUN8j7w7J7YK4XcWkXwV4fqMmjKODvre4SKoDYTEtDbYEmATKA
R7rR3v3t9moFHhV4Qfa4CnVnmiSCGWJNQlPhDKbGH31/QcHOmsWc3MSN42Jf/tWq
W5BkuVGNfkVd5VQU99AOg+FuruWfCP8Q52IB/s0TBPTaVnq60APcFNXz0+5vWXFK
pNwCEK3AT1o4/3LRJhR4CKJmyBWFgyAueYndh39SpVpDuPCZfWxPmeV42RVqvTD0
7w8gVCZP11jXgPr1FmUwvq+PYxwX4iSVDjr3fZXfyLeLtMFRrrJKjn8T9UA8JCAl
MqXh107d4o1KdS2r2P/k6nKetOYV1JdLn6ytdxCjtzfCYo6jV9UkFvRvwZOjwXg6
ExpkikfFG2HWJBwhxz4AM1HhALBMq7GRRzexT3QQxB2oegJWOvMZgXnKtc88hKYi
W9Q1x51jzjChZ6KyZCdhDQPZZmyjdhE+fpmhN5yJIILPeFiV3fTAc1s6URlePjYI
07tLXCx/Ft233LwHmdEODww2Saigix3sa6a/xG/07V9HbjlrK9xXACgUX+Wa74n0
os2FOiC0D6VvqnnvULzatJgIrHU7r7jujbGLzMprpcYkyfOe1lfY93ZiZyEE0OLs
J1YldERYisd5/nUE6v16Jg4LL+BTsn2qtbqPrD1CtdY8vcaIHg+QNLN7yREd1sd7
wik0aq0Km3VPKohO9z9wZfSdwkivl7RDS6qbE+yp/dODA6QEW6nIBb7FOnhZCeSs
8sSVUgxm0kDewrC1L16ELXgu7JbSpgj3gukLOGGKTadyyYxuLf1ydOcWblMGuZbg
iLK4Z0cmkcKjRGNYZ2ATkdzh7suWtAmctZJdy7Z4+cVONnA5wNiktMazaWtzX74p
aild/jTWqAdAqPcYQVBZ4efiIh1YWrV+lpc/O9cwE2KT2QzKE+eO1cFC+ZB/i5Bd
bvGBsgkavSjeaxek1lMXUbs4sSJvt7zpLn3TyVaiYrdT0a95ViAihe8clLdxxWCk
WXLuuI+k9cZCRKQ2poomXBraRAisxybITDRj+cAaMVdmrdn5tL1kvt0nMwVSORtO
cbg9hD8tUJ4RA/qZsIsFYVc+G4P/d+/ZAb64Pkx+UoRtxmEBA4mXrzujHEB9cITE
OCfD8ZuTIIiNC4iRkHQugDa2YBKMqCO7xv2NmjLWMg3eT5TlhYo31Q/p0LKOlskg
Z/tQDrXVK4MraN3RbKA1/7sMSdF0O97UI1+P5LIUQ4eVDSfMeCgo5jOUNzYDWjaR
jVtv/YoxyjAiokAFvu/dx3YOjAuAuBHUF416wC4LIHE8Xs83L6E2Zzsoi+EBUS97
CJklSK44MzUnq+5kh3rrmNz7htVehOHjsxpzTofxEdhwtFkI9I4BkKDa5Ejr18bv
R43STusOFQnLd+AKfuSDiJ7DROH/9NVnmOSu2rcwqs7el5poISxWwzWc2sp0K4gc
rE5j3Odbdt4qzAa5sh7jwnaGNQGyin9dKI/TZZpS+32mFA6m86VMPkdGnixiIs8q
T/QlcggXSilpVdPjhVlqOAVu6gb6jsNTwVaKUaWizL/WGZG/l1sdg+3H0UCPAMui
2YOk94VNHghcIjxtZdsz9Hsh5y8uRMdy+7xD3fdy5Y3pSoVcvAqwaVa+baeVJi5V
jhmlifS9nuDFL+MPWkY4lHuA8j+avwZfqIvsBwyIESZi8cdgQZuNe2+B94YGlRlD
BGuE0sRI2v39OKf4DX5NztWogUjPXkaBrRnDOExxEzSSreviA+lpBiUzPs97LgkW
X5NetaEXZhI59KFhORzhqnWbUtHxorD0oWxl5kpVOdEmH7aksxHHEJN4PETAqmPS
4y5Vw/7wJOlIbAcsq4td86iXNooLhFy6ET8JrpYXhYq90GZodLYKIw1JX+lQ9VIi
Zk0HaGIf/vEZAVkacMls+BnFbboX5+ove3kCj5GZVVsUE9LM8AJoEaaOgzA4+Qqz
cjOQLgg4BN5BZtkAqVS2BV78IJN0X+BD+78AorPapY8UJ7lHocBbWmhUERMIv/kC
5sIXWaTfX6M9Vhg/IhyOF2c42cM3QkxoWduABCySdXsmgPSF23Agk3w9gVk+aALj
shcGDmcQoeawPKnXgaF4ZZgWcuORQ7CsFxL+25r0avvu6Zh2caCMEx2F4iYn7Ki8
2ds8bDoAEvvYT5KnuAlQN5K3qbrK/jq4aaUxo0zbOjBfklhbS6A6FLK5Cl6BRD9z
IQmF8VtuBrrIA2CRJOgEjtWjS61PTfDk8LQ3/f3JvrOyViskC00/BwHw83DVv6Sg
LhuH4YwG+p531cEMAURUZKIaX+Qj5rtoCLkp0011shA4Sj+nUmocWMUq9bu/coE+
10TT8hjr67bOF5QQssEHAMMpHbRubo7Xu5oHxC3va8z60WMJqtiAE8uR3Yjnezk4
1J/mtsYOqEMZzRSEhQvpjOv0idoKjPvkRUyZMROkbVUYgAH7xgMmvcpCJ8sx4CmU
6hRrNJhAdFCqXQAWHVUbaiqm5s4l5bS/lhgHhcFvQebJxcpNGjMFVaEqB90ILS7F
6OnUOpzPnmyR0iVtbTlTlWA5Bva46OOzolf2y3LUsWphqJULOFv5Uw9tOqttTyYt
O55Bc9rio89+m8Lf8wOXpkZdYlMvmNoPpD+bKtdM/7rY7yuEdFhO5lr5aO8J4OVG
8vyg0you6jAwoyieHVYyzryJvQu6wrapXQV+wnjGLJ7oMTQZcY2FBupEfpBoIgrA
DF4xICQEEjdIpQasf2oZqf3YblpZ+Gft4jwuTjN6q5jA/bBvnyO8QMGXoGtO8ZoQ
mY/+Ak4VEDY3dNu922VWNzSB6MuvZtmE9yr0EnYUSdnYtvuwMI0RCHdcKYq8ePWI
qkepqcvmVt/ue8ClkoXEHzRHLG2evp4ZZ44SZN8vUrYbV/idB+4aQZyeT9yCRlgK
euUNRcaT4L7pCDl4olRIspDQJlGDEHEKwm5y0hsP4/jVnY9VzTuVWo+9fUM0mjqf
brHivJqpc75gd0GqHRZziEA+BWKDjUcW/8/YjiahbIUYjoFa7JHFpDIP9y5lOuMI
1gySyzosQRc6UrQWxOrZ1K1n9qzOaRDzxd4qSjRPY27nKLlhdgCdYEq9D8iQe3zF
+zlBXlb2DKosncU7IAVP3iakM8uImknmuSVjnhTx4QH+vwaJzDqf0bCPJwiUi9Re
m2YI6FLDZl1snjeWt4VRWAWSrwr/C+8OS0aN5eI6bNXJnHfoJLsu7r2XC2mVLTxA
fwZrUfQz29k1L6d8xNRkiODfkp94DWUZCy+ib39KdBMNA6qIJYmzW0NzMf/mODol
uqiwNxA91oMU0h3LWxbjfwwEe7Ufg3uki0kRhYaR8DalDiyRZHa4wIBkBJHk5dwQ
AGGwMZZIurJgv7C3mfid/GfqcIdc9JRTftNX56yZKmaK5pyVN1yysaYIpdHIUn6H
1khZnl2+r8mq0JSnPKdfOltATUHdBGPcXwfax0vZSJgMjCRvusV9lLrir0fT8BRY
BJxpDKsRjOZ8q+K3DpGmkPdMZvnDc06N0x+5vdt4C9Xo7H6pWVTKzersOXyLOHrv
bE8qRExiKkU3lrVJuVgTB2KvEsstR0r49dLsfgMeTlZ/dDTrUa32FwclxebMJ4Je
0eMM7GpzXcc2lTHtFoQamDHjNdlhWBQuN3jDRSYdraOuajfVw8iusM5of/3xnS0a
hig7Nj3KCw0YwX6NJYk4M9lsElI284RJJ46Tt5RNu8WedIc2iLglkwswWKoVzjOZ
tfAM/R7r/vOQ/kKuIsFg+PFflAV1eSj4SlurceXRrpiBUms1DPOaq0IIenIfmAjf
gD3A0NDvA8sWT0PL8DeCRig0B2A3Lpmpp0j17Fh88M6uVI0LYpK/rxWa9/kUbBnX
zEedzBepY/Vv6G582TZIw5IKMNMLDWGWWAYyRLvk5Up9tIme31FnMNedkFXGGz4A
2kEoiBO4Os6DIReDmiuJG1Eq3FEYHImrRHGuu1nLUUjglLqgq9Ccqub4EICkHuDn
y3FUl35Yz8jt6VAYsLx7c5P2SKXyWjJ2vdwn6+8nGKlHXMGFhYA6s/3/XfXOjvWK
gS9ovN30gJCnZOPYTiB4qZVsyOLXAj/+jaOtwt/wK15VrWMrJP2hBhldsRk9Kx8s
sslGHoCwKhlfr56pc+u/FO952dqndXUd0pQ6JGVwhF1o66iA3oQyRQUUbuYiygfO
KdcZzExcb0D1rmsDQBNFz6966UiZMFda4YGsoWXqbT40WpOGn0/ox68fnPLMdFfn
UnA1/MUVPTTjUIRSlsrJ2Q73KQ0y5M5fwtgGwIlASeKmHfJ2mROKzn/aW8QQTJrX
Nt5GgLL1rwPDXE4PEyEgC69n24mYVcKgkOkyu3Xi3NWSa2sGJ/jCq0nQMKGWr/am
l5IK1tZITcGRxRT6FJfcyNzqCuABMEQwuX21+X28G2Rsnrx1qjQxF7VAgMAXFUpE
R0SB6KSyjq+hW72hW/AvnIdYIykxtRis205yeXZq/0sw8olOJjIr+cCezJWEKfoI
VviP1QeS5aZKg0d1LP5/aNjLcezCRreCu+bBw/BTbwOAAIiKtV3GuptnffJQl/RF
JNyTdtIlKJHdYOnQBs/UKZjhtgfT4QWFe5A7gS09Ci2Herhk8lUDH6Qbu1x/K8FK
jMHcFaxNwxzj/CXoRWdroouEJrQft6tHU072JWO3ALgbZIVD8TE5iOAHPmWdFAS9
9LA3Ekm7RsKZRnIl39GYRCpA1ii3fbWTN7u4NsQd2cNqujwbLIZpVYAGpiwMmGlG
tGIDq0VLluuTZPTI8B6XGvS9Mg4V5wbFJLnaCKeqqv6u8Cd0DM0WTfzv7UaYq6i9
IW9opml6K8HYO/qIGUpS3LUbeBDfVjaCsMp/Lmoob6U5ovdq5Nk0kEipbXH8Ak6o
/PiOdBjzSalABRH3ATlKiCxsBsxZWuJi7thFAK1PYEw2QcZkdzIqeJGGACgHo3s4
fAHMZZrWpaOmTzrbh+V2ySat363mMu+0VIye4HMoLAGo2HxyBSF0fpNmZAYjsnbO
qI0KxKnQAeMKWMnG0HsB8qoWTNOk8ktQ746mVrGiw1n8htS2wVIg0RP8GrFknD+B
DjQSO2hf3eoa8mqcU9/0lkMec8HmoRgH6XO6s+AWHq3Fkmp2MUJUx8IvvnfWbgTB
8SX30IdNK/7JevU3l9RkIzq09ww03ylqous/6g4W9PjftwkZNopAR5b+c7MWjCe0
crd0agWqPgF07o2FtY6IHKSAgE4AB6RX3OboeFG0wo52ZwMx2RCYVkFUdTpk0oYN
9vWS51kE0K3IVopTub9V7Lo45akn7/FcVHDdEC4nfOHDWSPmYaTpo/0xGcCnzlKl
xLZfc6a05kxowriWUJ+Q20g2Cs0ae6O7NlJWHfHotFeB2asEDc45cQydrSJTQrG+
pxSvujYr9XtymA95KpPBRIETRIeoPhEh2jLzUD2ROtJuQyumr4d0ehl/5Lus7meo
CtzvFOBgB4kPvx1edWeA3FCRcEcW4MmNBPpZu8fgG7QiCKyC/mGwobQL+6sGGnvt
atdndU9gMs6wLPPVLlszrmo8ZDZTlbZ5GRvm1ZEmoUIcq/KrNfo7aSh2Xq7im9EL
Ktq/SLi5lpLrOL5+8xMrde630ToERY4LI/b7e+LvGZ/csOUu2O9HAo19EexLT451
ds9X+mITaiEWpBd0lZ0RKin83AWbctpQr5d7Td8d+6AW84EkyoXZlx346TMFJRgh
dTBhd4Ue44GFe8uBvSmadpLv5egp/Cf3mzSkja3ehzgESYmtm2Uayu/nxYmiiqJC
Ypenrud3Pec7+mVLXxo/lJb4Kz7tmCmZJ00YGp1hxAtcIZCMf1NgI6TXEuf/UiUC
aFhtiCSfLSsizp4rsFAlWQx98wOf8TUca3EO+XG6A/3E6t/x6xENj6uyL7GwiSBn
T1PX0k7huY5PlUMUrRfjqUK9LNVyC6arzITpMrPJLselGsh9r/OY1Y9cCv5Y5Lr2
8cV8dsN7FSFVfZ7iHei199fWq1NkPoagtolGX4FOCHyMV0FDyrTdHJpBQv3jdQhS
Ox5MONW09Gwo8qqzX6dRiF1zDyHxkKmSXF8HoKxzwsvv5vyPVi3idXY987OrOUok
jYWE3z6YnD4Sm5W4T/FT0ByAMH3mv4niVxXnn3VMz/AROda6p0WhXmf8H60Iu8v9
bJ1sshJrJ8lUM9kU3S7JDAvGPdH8ftBYsPsxiAHQKesMfeE0zMmJn9OSg0O0avye
gFggRKUXAWtKA7UPYCrg7hWRE21saVFQ7xj3MM32emCkrK3kyyyP/R99S6uVGfpm
qHNwq8JUmt6b01s45YtNqnxRmH4HOwBT4SAYeuE97cpSJ8dpi9nlIlr6c0PUUGPW
i25ELB+/Fz1eZlfRWgO0/PtVr2o9MQ+nSb1T08TBnerOK/05aZfgbVJDu3UCKlJT
eNQAEtIL15qnNZHG6HybhiSUCqxBiXZIN/Sp1mBAY+CZrVNJzcwn0pXAgRsss76o
U0hvpmqhmMX4ORuzjHppLbPKch5a4gu0dr1fl0hOsDI8Qa9bFZGRlLWuxY3SfhHI
Pb71R3tk+YR+AZHbhxGbV00GpqJDD5HMBS5RO/T7DxnsJC/qE451eowyD1VEpI4M
8OifHbWmEh2OvzdCTrchrEGQ+r6d/StPPvL0tHcj39kECFJRS6CxAwFviiLIYVzW
P0CTcvSGoPgvKmOqyYAEuUs7b9EMXQx7WYIWfuVzks8NhPO4UIF3oyzJOiOMrg1r
B4wn8sxqg1ajGka/QQjansso6bSjeTJpAa/hGJYiILLY/pTnhj1oK1H7W0aU3y7m
hVha3oA1Eo+VvXQmjvgiKxtMXJreuQ0q+vJvZuysiW/e6X+EpwCmvuL9VgCCKFZO
+yRS4CVeFOGI8UMH+ViIq5/m0YbZ7yeU67e1Hv3OOJZa5NYJGqplhFxKcIqXEaGO
adVXdFr0jxkcxyVTYllfVrunoBbK5JV+joIb5k3rlWAshHCaxIfELktCjLwz0eN5
g8EEg/9SyE8cOvaboPSHL4vqu8a33oOT8spiP8O9bCw4ud2YZNHZ99CjSi9PCCVw
Ek/yok3SCrzgPjHhESV/TmzPape6sAZij2qRpiXFxib/uQ8cyP2kFhQnowoIYrFH
CIXKv6Nes7ALrtp1JpXLcgjLBEMUBdo3aRL6NQMZsyjHdtGM2fEMpIyJHIwzo9w/
lj4JD/qzgE7QpQpl23T3yi+TZFgGnXUYD3GLCyr/SP5X9LnbtW73DWdyHrMwfHKH
2QLNINlft1fvkoGyX/XASXXnf6KGnaU4//csTuajH7JbI7rKEcDIQy5KWjubXOIp
6JH0Mm/gXdMIp26/tygI/enX+SIN8pEQfLT3UP+bD/jvuWoqNuqK5C2y8i7D9alL
luglMJTT5MTwI53+ecBT03P4DyHOuNYd9wYyQyXtWOIu1tbWmufkSoU/XQ9xtu1h
yFGK5kjyQgVC+C6l7IrYyFOYsF2fmLCqrrRAF9HUAmrMAUkKf/UQz896K/nZ6zyQ
8TRqPVdOzGDgpNCuQW2GSFqZ5a6OEp6RTgUZlWcHhyewn+5TMKpYUuUkekqv1lje
zjB4l8NxnRABZx3tiQGZxeeSg5/qrnCEkk/oiu6O5Sya+IcM+sawUFUF2Fezxzm8
0Yk50n8ZehGSW7SLOESIGmrJxNWqXho/DBAN0sSDwyPqbcn49+fskURj4CHhzaFK
jqp9FI7905hCodNdoVNtXthmySqds9TNMHhqxGnjEjJEwR5BwqNrEHexH7m1kHP2
u36xR2UoaA8/QxiNJwylbbdjC3/wYxoXSHAWmVMoFYULSftxx/GWdI6U8j7gYFAV
tMJYT7r2JPmZvGTHP+kubSr+JbyDgihUraESTyMgHQ/XiX3H4o+xsh2UkvLPOb70
zE2LiVjlJhpTMglgdgVeqpVfk9HMP5ljo7STEa+GHalVrF0zlsqW7D2eQzOHWgN4
NC5wyOxwqOg/+wH4n84gandhJRGLGw6k281rFAjKsXQifXMHvEmw7a/We0bFN0jv
ww7JrjU9qrikyJzRTHwFFINizFCUH6oyJI/U9RNhEFrxLv8MmWcPUpp8n1Pguo0C
UaqK9+9wUYGnlorFFiUkX+2vMhuEWfW36pzIkuFyqhguaEc9zrVS3PR2XLeBw0Uw
nKeTDYk8DkG0Gllt9ryKIZrVCwijCppGYusEGnm/gbFw/cqhPQIvjWwaWqdSFhUq
oO4mQgu5h3S7bsS+izIO6+v8n0bsnH4JFOJyI2XWiK9QGfMNuDANkfcGEEGQ5aDB
+M15vbK8hDS8yN3O77vwXw2q6HKFyqzsHW1w/oF8EQsShPFfLR6m83/30ZIkpKyF
3+qA6GJp3f7qbTT6YDnGncuFUXsBY57am1TXR+UCd8qQSSdGNOimpSIFP6BI8piU
99kVzkJGEtyKE5dj1IERfIHBMjLU+9AsbigIOGd5GTnqbjVJDKhYBBGxY2W4B0tP
axGpPAE08Y1aFAEaEWeGok/nPNpatntTgSQftUH0Bf4ePqpUD7Jq4uYSYa9ePPz4
XjIRftL1ZcL2/OgfQWfAoBKcyeU0U3OXByHGKVy3RYCUGBM/1hjGUcZ4q73pxcIL
Zfuoj/ChVhlMtxpeO7wMx6J+DWIFkpzy6uHyXlbuuuf/1Z/PygcfQDhIMNvUatMK
rcJLmKdSmATZ9uXh6OA0dmiVjBAgZE5OVWcarJ3NnOF6WxCuV3J9alNvutuFuNRo
h7gl7kDx01gqSaKaL5LZRp5bATs4w8i+MPVL4ne7m184StILKXu6mDJblsSRdeLj
TI0h9CZ2dX8QCNvwVPtzhzaA0+6uHFtIDXKQaXq8+o/Kuq9lNGsqFyqGxEoKnFnq
QUEjH6K27F3fGbvioARXkrGdOuctj7WcMeGkluLmbfSEknmCN26zTV+bMKbdC+VM
+//UVPpCOpOVJzoNxmoyymP/F6LBv0ToeYij9Lc7NE43WDeETUCNqyrfFnfXy+zL
ZEjn7ucYhGpZnp7m5aXvFraKvbJSZOzDGxEqcKbJG4F6YwYt/Z4NmIWYRb52WG1S
JWyhzZzeKxA8iNoop/XrqZkfOrXsDsKWhxUpSvXbc4LK6JojDh7G0f+pUaEgoalE
2kBTGyuAL3dLxpUfJQ4lMP11G77wxQ/ywKrbziVLEiyaK/aDicgv3OyJQkN0NwdG
2nhRgFCVMDhRZ89kNAf0jy4Kavd+rJ8aE+Vo7VEZ4+wIKwJ3HArqKJnmd+znDtj2
I2KfsB19jd65mdnW8sxghJ29ZztXkP55qU3QwQOrCZrU+SP9b2k7uR5ZEyKxHMrX
tFZaZUtCnYufI7HVYLC2USBjKaO8pAwm24m4qQb9tUhDO6hMB/PF1DgQDej2cMwX
dIKyaMNFxnGyPZa7hh47bMOar4g4VZ+XuRUNKmK6jrUMNoJhyK2Zg3SFoiv+wTP/
VJvGEwkTPNBCM4nV2kAswRRnkqIhvHaUE6i8O2WYtx5eLYajnu4dLTuD2taBwdKB
Jq5KYSZsj/nSCp58CaEqybDd25crVXgYGpGS8uuOL3dlW6rw4/ymPwM7eS2l3I+s
22ZY0poI/ORy/532dgYYybLUWGKNDAGdIJltdz+ULwit76xyuIgX2K88vboisxJx
Qq4y/yu3EheNBVZH2+CzhT83WUTYvRl1Ijbh4z3iuJ2jxhOAYs9vyHkbHoWg2k08
qDFeQKeaBFVFi7jJo7sSVRLS3PkPvXXkia8rhafqoKfg0++eZcxbDdb39Kpd6T87
cpvjBii5eEx6Z/myaHF+c9pWcA34JYubjGFUalEM6Xq17odnylf9+xDiBhLUe4S1
ZWV4MtRUslSy5jTQo97HgtCjXR6p8KDcwfgxZSdEHOS1b4Qtm0ROq47gvOJRkqI4
NZn3HKXyhFhZSa/ufkuX4/+L7GxLQ9iPME1gwZjmzl3btpJh4yk+NUGmM+Yz2Mon
QSIwI+Qt6QaNWZtA6JB6F6cqy1zCvOpkmQv+dvwHq99N5F4cd3RFrNHaeuSgpE90
6GbvgDOmT5YBTgwJvkDmw9Axazl1gk0AUTT+Vq6N6506sSNqZmC0ti+T3qZJZdzo
oG5htsXYB6Hig1WaClZ2C4CJ+KIYSIDykS7aI5ilyu2UBxLwC/6UcOH4Hal9EPnM
nVfrN7t7nBU2FVMQ8xos+zUEzxJKtI6bIMbjVyqzRvZ+jr/HK7EExKaAO/lcaKOh
CtyHW2gTN6AadjK5IucWT6PPIAzfnAUwndscJSPDcLjwytuQnfhSmh0Dc66H9jSC
zbhwveaoAL7ENQ8RTsP9mX75smv6V8+VHi1mBaEh+U3OTPdQJ/30CIZjWQTyX5Lg
ihKg8XvaAlx1cgrTyCR4b9wHWVyKtasCTL67jWvhz2X+dCjjM5oCtIgqdD5nX5MO
VidmR7QAWidUigrrPL3pYwqfrS4JOIJQK0eLiCE72TJKUoVGCftXREY/YAJkeaZ5
YUWIj8mmw3a1pcnOFTVEG9ghZ3IwKBJBqaFBMXsKitFmVWW06mwqvZxBe4DJadiV
Oc93D+qaeNW0oqM094GCVpoJ2vBMdrEKoayTHI7Q/uLSh0itx2G+81aYUTmf3QaF
g4Y6FbiSuYc/Xl8w0kjryoEOLvI2IQFwPtDA+iqE4x7KIKyY0Ifr5vDFNEKwVkzF
4j+3jQVTJOf5l+H9ZxaldDAMn5iyrqk//K+MXMZYTh4Bs5S7pkAzEjHzN6TWI8YA
rPWbIqEWikDYIgQ4Q4wShGzyd4thnu6cyCqvfc4e6X1/IE6Y+Rl8ese2VNgn/XAw
jx543Su34jSBJbv4ixcuY8AWfDp0XKpUY5FCT3fFYQyt8vRXZTWqMNGiHF/Qv+G0
KmTphrpOzA3qXUVxOyPq7NDCzSS/t9fi4CLh3e10dvpKzNeyOBtkWE70VdklbIWB
U9KbDZwu+iwDo+qoGB9ECpPDedCrclbOXniSfMxdjdOnhIJFKEJ0wdkd84QJQQmT
9nOLn6pz36JSpMtk91kt9F8C89Usf3sNwvT8Ljdib39A6lY6Pp7nOnaXPmyHSPNi
uJPXZt7YUxy4fVqiCBa60VQa45qOFzjRHEo/PX67kmDGyYmtnG0xn89Xg33Kvrz8
dJWHVUhKwm4hn4MKyxphXXYdwg7d9vzMyuDXY4zYYUZRtc31bHKVg42EZfynMe8+
5f8fFDnckWXfs52aK1HkVoKD0NhH+uNLhr40BqB0bYcPPGeBePOgZ80kitTmhFlz
TQGs2vKQJPOP9MRlxZGEgtIbNLEhSj3aT1Zw8lrnAFza1lu71Wo7wylY6bPI0PA+
BWtFmO1AWx7G4qqPO5j3luHFF3gmyWhCX87RAZhIKoiR55pMxNI975CcZhxco3RN
ena+XEj4BjmyG28yXD16opXXP5IlWIihrOr1tNetLlfET33DHGwb9Ng6hMDWJbdk
/b1usLe7vl+PrlVZP3a9Vp0Xkvub6aY5Iry9e5Jg3XSC6DjJht5CtNSzOWDGXxEJ
KZAKcblwJao8Uv2ZOSQTBG+t8QbGXCCBWrMTOlX5CudKu7xzkuvM0EQJSP4rehZ4
HaKjwHSrubGSwL6XgcCGSlw5tNSkjzXP9/BCqIxVtT/v4HRlSKsNkBydSM5KJ9nl
pu2X2Vd2HpPlI4mc43izRI7fT21YXvbyiqiblukxnZQI0/5onES2HUlEGKy/yFG5
u+Dl4AaFqupLGomNBW9I7Hm4he3yG1NRkI2d2eChIxi3EFCm5+qUV4Lbj8gjORc7
FI4gx8TGMn9uSqr/MLxXRD+m8JJ0zjMlZoeFM9zW0Mx6FHtvi7An7rQwWqEKr0U9
LkIXe8efuu1vBhLYN4orY0jIvJL3OgGF1z5m223FFSFugRToluGCQOcB3oaJhX69
2uqpyp7bWoiryCKhJbawcIPWTwo5giqdzRjRYOcv31QCCwGJrg3iWK7hrk/j4LTJ
yb7Et4+Hp34rSrPom92BKffDU44rMcbo3D6p9uUHK4Jn+I0WhLUN2kUxJgCmTxFO
9u5HCQR6B9AkwL7M/abCWMUzYVX2mMn4M/DoKM57ltN0Gw7OJP3z+X449fmvn+U5
8tuUuA+0/2wBVSnZHSrw6A5T5v1Fxlyg9vfOX8PsJQ0ymJcCW/UbAjugPl4WhpfH
biwD0yb89TGdGgB/P1tdRDxlVCq/wD5HpdSdPUlFcrQfVCPkGPbk84kRZfnpOWMR
CpKC3mUwNIBpi5GSZRPg54z52TSxrhPZJe2fjZUNsSvl6t7VhQT3FFMn3ieSn44d
qq9egdyBaXExrI+fR+rhuajyrQz72nwbJn5BCFsXdUP/Dyr0SJ/CVEgyxZ+eyMLf
CXH9/wDlX+u4Z8tYhRhZC7simIBX9GLZlFMfiIaR8y24Mm4wgiTq9eiFCAwN12Sy
aNg/uW4tKc5W00Epq269aML8v4vh4yZA30pU47x51CEBexS9Rmh+HctROML+H02E
zlEYHiD0qQsj+NdBAcIxdCpyyPTdP7hia1H+djUqHSCnr7wbaltJYxHSxZUKnLqG
Hl5s9QJipqGK7KFvIzvSpszi8GPfICmR0/jIWK5GPKH1bpSFtdfa8VRPzTRhSHf7
ARpHzg4ap5OIkevXRbn2ETuO6uLO2QOVxwWf5JBA2S2mOFQWo1eNjDgppJdatkCW
7kxHCWIZ/VbD9pVeOhOYwwYhHwwQKqiKF1akUbPzZP4buqw5KO2eBJkSUn4tOmcp
vZvWJBs8VMNulhTtSb9LmqB0sJNRy1/Pzfhoe7b56NHJTJjzj4yY9l4oOpDJrAhW
muQ7rLR0SbA7pECd2ekxln/FTAswbf7sN9/3kgvpa0AqjDP99I+CgoMmw/Ra5P2v
cWhikzMIJRv4jdywxDHukP/tEvDDq+PM+8ss4JKwUDDryVVwVp0u94MKwqP+RMAv
L9hCYj+z0GH9ekxSJIkkBFvrRkboKE5Y48//9B5UGsCLgY0nH3z9FVEWCCdNWNPn
cQi97r6f5aC5ooyiHvsUXAYW/pxE9ycZ7PYUH/1YaqCAf53UX6eZHG36fih0eCWy
AyQUnta6z+c5XIohPvi7Un8R7V77Fa4ln6BIUXFej7pKxHDP+2GTiyfO86VjG/bH
nyDtpGq34dbfBdS+OApTjwXLZoSPBMClo46by2PCimLrxHjaWRK5PwcaRsMpVxoH
wheyh8wpdM+Uf9gZqzVP1Sn8CzueIb0lOWOlaNR20eTVB8mvF0Zu7OtuymL5uVjn
wMINHwaGvj8P5ieZ8b0+fOYNZPSVk7gf4AXP+Ob2gUNFZ3Tg069zX6L/NUUBdDOd
yxxUq6Xq9dki1ffW5/QK/PZFpnbtjO9ZsvJTX3ShDrX91BLx0oHuxOmqWGY8H4m9
7fIK1nqocQldboYrL3YWSGehurCI855VUc0C8twp63m4BA+6rdN+PsXz8Wz3bzuA
bNyl4mFigAu3yLwlHfUtNdlUxtzBzJeQ1OAcnbM78keZ4semil7s/xMuk1VFlKMe
B1eAgdgM26iMQtU0J31T6GhLH7aDFdHIqPzHphQ0Wo/yLBsG6C08IIDvHWeCYGlj
jF/fFsv1ME/szBJdXUH6rRnMiiMCBW0vXAGRsRnrv1YDF6Nwro0KmxsH87eikrVh
Ag7ayrl9EoVeyhN4qJ1t6ERaQiixD8+JMHHUor87nAsLfrjZcILbbpom7TZ8DmNT
1IaETEmVxsk0NLW7hG2g6oY6vhzi5Xfz7IRkhhxztF0DWygcPjCeCdGEJFkiIUFN
m4FlbSpZog9xm5JMJ+rE9q1mnbsHToS0foJ+xvajNstWC9tLgRw7cqjT/HRoneC3
H0JCzGhyIyklHQZgGqZ2dGZyrqRLtVeBWplsQjI0N/uK1dpNXUd4oAWRaetVcaVs
5dp3ChIiqnayos6JvUZambN2mISc2wJAYU0sdZGyV/QziW4mruduLq5WWaOiJB61
WOAbX/HCRkBzl28hsoPgDUR6Lg217HomW+zNBZ7LSAj79mW//j+OzhnwR+0rHvaX
85PtpsG+tPwU+eCOREsFikiVpl8wkTpLYbyVsmPxPxkVzgcm0z75ak3xMUQTAxYK
8qb05OgleDjwCjx2dVpKUXlQ6K6ry9OICfk7j/HH1AkLfgo22vtBtX+/Mc1r+yIB
5Mrzd0rfJ9akCn8nO4chGldGGCbcH8qBbrMHJ877PliaSIW/y/jQ28SZVlRboAAo
EpcTh8zB2Vg1gp8WbUrC23df/JkWhcT/5Ulnp48ivYbeMH4gYq1MCl3iNsHGOOgL
FD5SpDlidNAcK7C3dn5O9PxAg5pQX+GtJPke70AoJY4woI3n3UL/q0V0/E+EA5+7
1BdTcG4tsjgUOsFGHg5iAKdNZLXiRCq9hO7KA44YYYjzCJgGBGPZWo1bWCwf68pw
wKcKHY0uGQFZD0/ibtroNI8ZL2oRSMovahORwVXEPWkGdjwl9Qa6BPGtPZzlAU3z
8NIPKrpiP+6Z9FjwNGHffiuuhNgB1MMZh0DyCyqHhMf+cRaps/oL4sIGWg9Z8gyD
ZTkdd2FP19DUORkDdo3m7OLRjGQGRUSZQ1+YbLAtt5syh+r7ImKWWb3o47rHK5x+
dNuyuitpIdImE4Ekw9FQ4k7E6uqQOAYvtIAMsr7dq+dkQFHMY7Pip6irZIrJaK3L
GpAeXgNUtiYXBKiX70xkHjLfv7WwYX4lL/cifH1JlwT5K90RefT2nDB97VsWbz/G
ACEGN2L++j1AOe+f4ca/XC3tONLk2y/JHLFfxJ7iho5rkWGHF+OBQ5LaQPsy6WmA
U2xd93nLxAEkIlQM7jO7naC7t3xAYQObkvNPZEGyWxe65MuRe/efsFa3atke86Qw
tv2Z9JvuLIRK25z7rEkEjlMvPSNCAyJI2IhgIaPWAYZQvCZJ4SlJOVRvFYnewz+k
g19coqSihX36e8/GpaORhIyZK8b9LLBWmAm6OTnCfeujsdfw/iimEkQ5qbIOhQK0
sJTz01AxP65J/Pl8+AtCS92IFNXikRp7+YeJWFbcLLu2sci3smELbx7obvE7IzMI
hEj+nEMPSXJCUFEPZKRhZoRIAcN+VsCDLQMRtZQaIhUyBTnvy4YGvx+/YAAIuH6G
le+tOfD9v6UanmWLdMDDdK/QFr3/k54Q5YZ2zmmWKU4WqTiBLqyBqWXdq9dX1q0S
zynALCnjWu7PPKSC4tDbBnL7ZzI7NZeHV8E7PCKJTySUD1XXKZlr7RJOs+gTjuZ/
+GWK/YMWsUAj/Q6BnGOzyZiUI4x1SNyRU5jrFS+dT0mtuH456NBPM0ro6B7Q2ekz
C5dYfqW1d7AH/RedMY2mHhWdHGZdwP/D6X2wHHSB22eFWc+P1L2apGBV5LQtLOSK
AJTnnOHLfX4fI9OxZIyHUMOmwZ/FAbv0NXHQKl+GdP2phHEnm53B72NGr/qOFqq/
RzJOwiTtcPbCay0p/C3wzJh/69xmrFenwmQ5bHQR8VLZdHoLf2GNYcKUCuOtT8ZJ
FHSLfRoxAXWfuUHgapSLGN3TOqPc8IoWcI3Mhu3zcYZR0EuvgKrRDyZRS3W/wRmy
6BnXZTKAxMMPyR9CiWkIL5MVehw1b8c5ISEATjIt5IBB4ACJtBAwnAHrQV5QFF+T
uLygM/unPl4uMy4VjR5IY7DsJeHS9gBNHAe5qbytmVjGneTN4vE2MveJWzCPhY2c
ZWhCwd1LbrJqx7jPny72pFEf4ZTwNjcfrTTLeglkv75CYpZ57wyr7TNOQSneLwdN
lTqIgo1RSaxix14OkCHzdnN52TQ1mxar9KKvzgBQqYSNJ5XWqNCopljvQVXNqZnT
zSMAGNIwkYgF+i+dI1ukiUhKasp67aobUym0RPV7pVniQ6ol0a08sqoo4ys1/qck
LQGAcoOWZXsqnY8oRNuo78Owp4Qcu/Y1C3HqiTLvEJTtsJLTVq3JAtO33qgHztyt
3E2B1y6bGmkiXjtauAXAoCtClKlOHMFBfWTPkGSCUDxw0q53g3SMFYh2YfRZnyqV
uaPfEch4nI/iYKYE7pdy9KNJcCnBoYx0YZTv9S/ata07EuTF799ZmztOEAPuIC1h
J3w2kTCQPndBqNvnIys8p/AVggAzyGdhADNtYu2LQojrjqyRUX6MIc8FUx+D8yHi
lPcKrlgi3xRWf62AUc55NDFIuhy7yRthAJjx/UEyAeRrCaFa7IlYyDk1LzhJtC3s
+bYpusy6n4cw33fGvxmQEbWNDAJ+Ta+Ur/gupCJ+ESqRAo+MOSb9QcNmLVTSG2LP
zye9/eOlutd+E//zyZnqNuMH48eNraxKzzrK9wcdOjcySX0QsDCajQouuQLl4Ktn
GlAYCHx+4QAMcEoztPKk9uaHPY2B0OWjPQhoTO5hdeJU3PJAvZbpfqg+GgTDzMEo
vSkKV/6HbxChaDc9GcLLppJehatO1pKB/XsBhaJpeplCSqNvb38CTH6nqmbQ812F
PVLdGQc3MlRaKj9jjKBA3r7qQW/xoPi7DjjT27TqBqqEDYmzA7zDGnrRg7DHoNoW
DOau8GchspwxUylBEgqKpqOgWw3BgKqdpG1ThUr3ZZskpel/96fjPqEAflTDXv+C
TrUncbz5ncf4fHq9ErjhmEDPLutzIVAlmJUbu0+Zan1bJvw/bDNugZxGG2z5I5Da
QuL0gaOuDVFbrrZScha9XKiiXuW/dtmg5XWnrTjvlXEqrk1AlaG4XXJ1/Aiky2ig
A4WeDK2NhEQtY6F5pt8TAgZQcLaoEWax0PtDmEJH/gQF23GilQd3gqRnrOvaiPLq
rtYmgqhJzX1MQeKHkyINz4Oc8kvFDKlrVKJ72dN/PxUPT/IP3s0rHSCG2uZzv58I
Mo6IMktBF6/mtPwWjbC7JOaUFV5OPCLqYShQcCrl3S3/268p5O2KSnGM0Szz02OM
moVT+UStd0cEFiGO1OLvN8IplerhoE0Bu989M+aEdre8LRgpBM1RlryKp3fsKzMk
FGtkviXWQya3GFnWzPAT8mmSgQoXzq3vfKMoI1pSMk/CRZAqSxE5hNgCWsF4EWBd
5OWQKeeEy3bj80q+rJylQjYt9iO7kZfx5lo8TAKg/yu/ThcIqdc9KsRxUz76/f/U
Ei9OTxc+IA2D4eD4J+WEro1zD2L7dr/Lg8FPsQQrWRQSNx+CQPJXWlPv2SurcFiR
ci7gHPKC1KA335qC+j0tf+2XcznlKlNHdEBJQ4r0jxoNSDhneOVkW0ovrVCgGbrs
otxihNwdjvZNjJSgKpQD0S4KJlux9FEOIXdE2hF0WkHaXt/yHuQd68GqhhQ+jbFM
zrxbCGE5e1ifA85dv7WUtefuzGAbxKATRUPyZ69hXTZF40tXA0KTTF89RlKDDldU
feQNLm8bTtNPB3W+d8uI10jc9Poq72XQ2kY+X4WRyl47X8k/6a7ukCRPJ865mkbp
o3NIjjLREHsejFL1yLws7OCiWT5NBRF8dyJwRI8bT0tO3a0a3v80ss905KlZpyLX
58bQiy1lCN4FFp6hZ1qyANIIYopjezLkkBw9zYeE/j6PbbXSKJCvRDgNjkaVh+WL
hFBrDMjlXGd9raXCeQ9VIN3WKmi6juu+Zn611pba5+aON79+Cr4MtfuzNbBbGk7H
A/3EynHfiO1SkxVnsA1lU98jvbGe/I5YYVVbJXSuBUNXeKiFup3lg7u5HOawUHSI
ngQS8hVAfe7++B+wJq4Cq752Pq+bdz4WDDLu9NJV3yULOPR4s6wXpRuetlafw2yB
3lfcnY06L0gU11nrHH6bH8MWpo3eImgCt+Z2fCD9cV1fBkQCAp/Cmr+1LxPm1aB0
CVyt3e8ZGA9Me2EuhZSnNVkiPNT2Ymni0UKu0bBMF8kEC2aHJYoCy1QLPbYQp/uI
Yma3UuD8YW569v7aEM8eliWxiLB8DBjF80kDQGqq7zpT+RvQ0Z1WxAgzyZJTfSVr
30lHjQeg0hDOAUDI6cjZuSBIUWVU64Hz5ajrOIbdvHxqJUlpnNGKgm+5m5O9HPAH
hLLptvTJRbseGATQVDEUXAsPjIA9IXLVd7hJiu10qMpz/w+rKpgBvJIh/94KYlmX
GdY18ScsMQFcky7crx3Bih83VTMUUWRiZ0HKfLw5gB5w5vhczwGBtxsKSE60GTh3
JUH5kDFn7s6/eJPtL5WzjFMmdqmTqI91VhLQs46AfXof0McptqmKBwAbfV0naulu
B+hWJGdyDwe/xvzjovHjiHp7WKjbUrQOMH2MTO2/TqZBX0aHRkTQISbNxY4CTStX
ZdTDWCdw2Njze6Ai2VXxMaJKrgXDGAXjEo+8LbcdhPMbCuLCsFYeBSqgzAQXFi9P
PsxEZ7vBgleqeF6fAoPbhvFsIGhhu/OEvq1xmuiYXIkokPbVNiNgw5NRUqYqYvRm
S/90Wfe9NoKRdXZEDPzojsn6R6rA/roeaMWcarrZY2fA7S+lvO+g5pjfwipqLTCv
Ukwl8yor2kUQI9h9sVSnrSHaBwEeRcvCdmEBwJuILsVAKM/TFeyQxp9fogcYnuxn
tmnu6yVGLvjWHDnWO5Z60JqK5RSRO78pA9cTzM0CeZjMuB1CFmHCB+0F00vUaPk4
VET+azJlZj7AZH0DkP3ZtVgvwh71g/FFdZajUOpV4InAG4c30MsMWav0X7lqhnE+
xaQXnfTfogvWSSToemdVaJre9BXaYCJKJ1U5VOkx+wEjTQd+lUjOSqF05MpICobM
mlCWRaH+xiGQNQ5B7rSsw4uFFUfeZwpprswFsAStA1ADoEYKAte3cG6vC0SYK4O4
h5u8emw/1oeuyRtHnBP3kBdL1kzzeo64Evq6t2tEHmpdRwnhENppo/BV/XLE+Ku6
g0gg4chN4RzeNFHeyZoT99qR89fzHBuwECrYD5eotl0xvln180aQf5yjT+3k5n2m
lwLhh9SrVl4FZQKA1qBNfLH0ZuCx5vEb+irJjzok7Ke8ULMqYk6qLDe5mdjcQVqh
3enz3GW7OrHyN3lK8ZEB96gW/QhBysbny8agHd/URzoZbEHXBosIvZUAQ7CqmGMT
vIkQ5oEJDKDpPfceJCBA1qiLyuZI1ErUfeUwoema56C9IazmEbju3/Y5DBbpOuID
mErh5qJA904BxkW8vW9Cm+eEdNagg3a++lgijuWYdfyVY63KNWTsQ+1PX9TumviH
4ifHwem4MSilK1DppDyHku/KTTeh9nUezfhhefUeRJ0q+xC8dJGUQTQmEQmauBpf
scLF2hp5vYdTky/GipYVTMOTNIAq5CgjYnbm66fiZx66IOr649Yi6yrn/cVdVaAB
xSisH0HeM7uQBJVpLw2MtAJldUmhyXWpypZyHtQkd2zamtZHXW4OnIZcLtBEsEBN
Zxio1Az6Ob6vCmcqo1rANB8Y0vl9zlZI3CNYtb7uhWjWwaJGX5dOMBpTeNj7y18K
0/1mJhCTT0d/UP3Y/8xGVj8KfTpDlVYp2/2WLmEGPoCpjpfMfWQI6khqa4A0aI7l
wyIXb1dXw4thYOe1BhhLn+Uwduag4mwzc6foPw0jhCfa2u/W374LhKtmdOGhd4Wd
hgAfMvtbw8mRvqHo2AA9TlFZUkMV34cic6guVZqhc2sYen9Wjk19idL75fqFtgNw
RwQVEoaTuIDqh98Lu0mFowERTjKExnn9PiH91Ib6RR30t00LluqqgNgXhRZ4Ny0W
mE3WikkZhvt9dUI5ytpOiznqQFzQgvVn14/hyEY1pVpSz5ab99a/uam9pJkucbWW
bBBsS+nQkHid5OJxTOr6wD0CkkOHtn6Pm3Um+F0hcovicf1wNyFCYopX5CzDjrHO
EIu/EEK4s8O1HcOJDOIm05LHOiWI8GfAvYH2xrBy0edlxRDJfILjgEnwmgjvVGTq
Xa+yVUUeIFbbepQMn+PgvAVl3fRj8uEi+i2YO973FNyfjHmwsAZVSuBhUQYCOe09
Q8lHHdj6u2E8ukdZWs8Jfjf0MPz48olJ0i+HxWbiQfcYdH/q9udA09566zFqznZd
tphH5L/AmOSo165t35rUzDd4/AMbC4EQ02H1bAoeo+q0CwfF3TmB/0L2Yf2IwHBm
EPTAYDq+EoMuvu4XT/MXWMUWwFi60+t6KvXJAPwXKAmeVkhjATlLUhETgkO44J4u
mOiLRz4+yXCEYW3KK7aIpv9i9ZR+PlHjrzl2nqOQY/bPsGRAYD3SqlNdxMUHj/De
ayyNbQ+2NyYqz2i7YXjKckt98dboDHOW90YzeUh+Qc5TTwRvQoMKhWs/+9DnXVyo
3HwxXPuLc3+6phui1QEfituxeIaf0PiT28YUyr24qiZe4isHsq3cNgEnfaZ/Z84w
v4hnsGDN1BOlPTqM/2i1q+o+L77zZBkdarTC3b/5uOyHabqDlVdsrr0IV6rzXDY4
YYxSUtJyqD9LdJAEX/iEUq40FK0KK0peXwzycvocFFrK1CJdbT+RM3noGfLfBOsi
kB5PI4rEsxTdgIAywfLLlV/xKQrX9Cx3l0YPTn5JopZqnfmOLIY9da7uIHuK7Brz
sUf9y3HGJiRnA9soVQW05O/wQ6qQzhhoDF7Q8ptYRHu2r6g6wQwlHAxmZOgRnzBe
f4CRPhU1aKN0uskkjZBl0RyB47ik52Px/+d6do58HXzAk+0lcH3yACx9RQ5/bgwR
IQKKKatRpTNZHuMZDwjEFhk3lV6zXbiL23psHEbaVkm+xfvVhxRgvaRtsDzP1zaa
1hkIdIM8r/Yq14+aViguCxjzXu43x2P3ClHQizEfBF4xXSZ0s4/E7r+nWJTjleZQ
y+6CUS+WraRRLBsOCw3Xa24KXDLYX+rmPPhDazKZz1xuLL8A8JqVe3m5ypk21UVh
iAj+wAqRh5lO9o/TJldlLyreWRvNNvhiQd+ATLJngTnLe10uHWKUga0gCx9m9OZx
su2mCXKNDOCnuA0SrTmUo0v6KItVZ8nEFeVsEBjHhgbcI9Bz3HTuio5XzVxLZs4T
9ZhiezdyFmVzDY6HYj6a6jhyCAvKl8wo648PJMm9YDK6DFXQa8QPpVf1r68uAb9N
gdUbH7KOnHhJVSfWgw3ynEXRCn7Tvd44Rd2I6cbYdTzxnWEQDaS19RUEDf192CKH
xHHaY1fBsxb/ApeawGxERRa5A2baJ1Qzfq6VgyrR/IyGRoTO1Tnbw+sgCj6l9J3O
MqHeEdG3HLz85jWHUXkhMNwtm5dRAJ9FMqSxNSQgE2R9UgtZGnM3kQUdzjn8AmDc
Fui9kf6FlCvCCylClp6pJF82iwhb3ewGor8mck0Yw7QqDUEkDaXZHR4bB/+P0M9r
BtKMj6AAho99oQrGzFYyxBMca0Q1lNfr/BGUVwpsCGiYYaaskZlRt2jAVtKoBfAF
R4HiKT0B2+ION9sQGm/mDCcYV5IGtRNnvUr7vdDEgFJ6NFcwhwIxq3Jt8VmYRk4b
PMWTQEzSrCb7b5nOVUC+uSy4N0ZKeiX6O8in1+CGmIv12U8KABHWatZzfhJeKYYV
uZJXaNvJSH6kYh+CurWbaQRZJCUQ0cEy6ftHUBrmmd6VYP2x9jpZFXto5AGiiJ2g
PFgTKCnRquBbmiAWtKjpCllrRIPkaGE+DRCAGJthKlTnoHk2aZRv7DhielY95czg
0kMLOIawqceMbTO3K4OQGl3nLPCsPFTcW4YAa9Cf2i+7aTU3hh3KetSsSXXqFGvY
ZTDYjyY0u0UwjE1OSJbode1ZhKc6Fs29jMdAMZSFS8pP1i6rV07tjDRKunMPQWav
G51TnIcJbvPJdz2anNgwN0WhwF9gTvw1H+ZxhoIKxHW4jwfWnIH8UzHmXOKPhmyH
PW9q+KWcJzaMH7z7aqwSZtqjcyQU5e9pZMlN+GdYzHY02zTug66qsRK3kEN1Mn/o
37Yo/srRKj3LwJ8gMX5Uqt5A9LmQ4hxt3JMYM1gg43oFSPTT5veW6UQY/MjIFk7x
WnGRC2JwnVWXKo9F9N9hd2lMXt/NmQlQVapC9Wbh8fLLEOw6wN5KRZhiY2y6upRv
6FQKn0Mo7ZwO/Y375c1a/wlAyu/rhlIdMP8H34ZUvFm9gE1EWtuspI3lr9XovOAW
cNy3SKC+LHAJjTFPRbq5U5Jmq0RrelRngRDSrH6NfSCwiKP3kctn3IhwuB05JM0G
Qjn6UBJEJ/F+UPus9lRamywuSr3Ssx5PKwMFYQFXA8buRff/+lpCPyqBzJMQxM+4
Kjp5198emTtHZog0ytJziRb3xQUuz59J0p74944urIXZu4MSyfiRYtUx6gMR2GYO
Tb8i52QRRi5q16EdVjne8eiaEYIzZY+p+nAuMcjU+a0AfeSiA000NK8vOOBwPhIL
9XGIrcEqyfMpkUMOvkTMKmr+ra/AQoyqsXcoIf8LbuXm0+9NLTaHG7h0sA0td4e1
Eg2ouzZvnnKXABsq1v0gb0NRMMcN/wmqjWnyxVBH0yz69Uz0n4snKG0aJaWdkqxZ
QVKBUoIYq4lLCAARhWJmnDJMUNZ4f9Foggl6l1uyd1YXl1LzNYuh3sl0mIiV9uuv
Iz1x2NKUZqkwN0ZcPJupFHjjKx5G1tFj4r0InQD5a6AE5clY2eaRnacqxKha0r1b
PzcFBvt8OI9fHCk6Qik4fZkMi8JYPL24RXJVsY8XDH5EqcMAaxNg9nibYxd2ctZa
4RSz1BZOLbqvKv/iwE65j3Xwip9DufPDZwHYy1SLXTxxQhf/2BrW3hY+zpPFFQqH
mcXiQUDAFCUB/sPN9IX7aGQZQVCDe3Z8To9z0hKQguzm2bgKhcdUdtG8FYnQbk99
tHG2T3TAJcGURBx5Tqg3bd1BdKROb8aZ5Sz2aPKB6xtstKA9l5jhLbssx5sOt8Ts
8uXr9x6D0UdGuEYxJx83nQE5vgpmJuD6G35cSmDljaAwpRMGr+SaMToAD3rVFO/L
BVdq6NoWIZNSohN1RpGvcrGOyPjyZxzPyAtkvtuLwQ69TcwzVaPUrQsgGCrTBlxv
rfooXVGiaCwC921YoTkdhoPNnTe4a6PnkTnFKSnXffCFJigmfzA9pQgvGM/1PPVF
boutfjRAXIFuVGDF/PVDHYOY4KyI39ylLKYzR3xWyqKiDlou5MR3SkjNA1+IrKW8
QtFiRSyxKJtgJuzCiE2uVg3EJ+Dzraau589X1I4gpzxI7qfvJaPtCTIuUlyeR7wn
o8evZpB9uhLNw2iZrSCQlPgSua/5nxw0sZnyPeF0y9XCTEbwXQFnzz8eGa2ItFxe
rgLfABEBn1aY/zSnlOWTjvEuO4YeuPRbVxqt2A2L+Cglwjp56eBHcBSr8AP03idt
L9OQaMmfTmMQyFsV+PSFHUy0ox7KDYYU91Np8QNvfACmgWTcEEGIDPnhAmbyXBXf
YqJj4L1CnXLpo1Lpmd+icjq9e85+pUAwAHCZ3LXysVCWo7ZuuxIByGZDlsi8/VnE
ynYMlbpJITzm94l+QWawR9KcnW17+iZ6aJv9Vk9h+DMhTSmpmzdpoKSlnyIrVSev
ypZe5x7+2dtAfpx4j0F/Zg0zhh964WV8h9KTVSyc8RSm4FYjifsSNuSiLL0RLeVA
X2xVZ/RAVMU+kubq0LGQtmPboPuzFpliLdD7+O5sEHZqM0fKO8PbEUrkt4HqS2vI
ws0+hliru0fVrBWtWqQvd6p4/RDj6PdpzUhRoEekKDGZdGRvUbPXIMNOjm23+i2M
e5DL5vena0qqWQ+8Yac21XXzQJ85rz48nByzUDHsIdKiGlHSoiZq1RCoHF5TirDI
IiHGyPpoIrOph5yDpfgifVxi1PBaC+VXewBL1xmgzunZm9lHuEBw0SisLe0Txo8V
VdBuXuFDovKF/+vp4rJis5bubbIdFi06OJqsPgm1cQXRFFaUu4B8TEX9MSJZH87T
hkByEVvNIX63Uq580B14m+bfPcv2t9Rl7pRWf1GyxiPYzTEHs1FG3HLXX9vbANMh
g9reqr8A9a0CZNGcHa44kDuCx5GAUpJy+FMS6xhllMqS5R5CaXgJNA10rX6GBEUW
zBzpddMaKfQnS3UT19eqvmsa2V2TxyXG3p5HARaj8PyhaQOtcPPxrX/i7ZvICKAw
vg5Es64nqeQFkfvP0y0GwQP38yleJtBF6cdlF+ERop72q6Hnnldag2vYXboyXMvU
Tl8SuFSN+6ie8lbzjoHq+XjcXqAHikxy/pA0eHgTwwut8fQ7kSa+9zeTyWolweFB
VyyaI3i2sqiEXO7ct8tzFJb4mkqDPbmL6ZanfWTGwLmdwpg22qSSJIxSfPnQvXSv
fADQSptMi9sv0tdQPOh7noJozhso5+sCR2unNnPUugwm9ZqYHX6+eICEzHN/tKcf
r+K0243tLqak0uSTplrTgKumb8VaKscfCj0dnHOxTqWuFEoPrMYrPvDCkmvrSrRV
LXRa7oaBFOSFQZukLDm/kLxttD4Kpe+myldirdgeiCncs5JnoVFgTEsvWSC0CBpY
94vnZ7F3BD5pK27q2S+Kc1W7kD3uv7KxGEBTADxk91gw1VlsAFibQHe0yC/1nf/f
MO8CWZnkvMhP+tLJfW9skyfxn8Hvi0RBkcz0Tfon4hmMM1rlJb9cRnXZwiEeeUhe
VCtoZp1OBOimIN3UdNGo9PcV+d3IJ9drDObv4IM6fjyiqO+4g0BzePIYb6bHNMk2
Dy6ABh0GwKvfCdGMOKd7UU0hwyg1ppjvRqne4YbTRD7ipVS0jdRGMdJfUj1UdH5T
LjQ6liJ4dX6UzY4/+TuD5qSqOWgyZV/A8s0knEViB6HK6VY3Dr3+B1py4ZW8oOLF
4duIbv1d09mZqEOgFkdBHRwIfyhHv8aiuED/OZRMzQFNjAZSt6C8+rRp7LYcOGJv
yQ+lKIjYcU4tnqWSGYOgcZff6dHUK3fqTePkR5uvbAA523RN8eWiSg0RsbWr53lB
3qatG68Zy68qQb1RbGJvHUdIbuKik+l/c5IUYBd/sEYAVZn//bzJlJTMyWQGEiy6
7lfU7U2fs2MecAd0Kqbi6DhvEQFQmKJMynqG8on+9+qIRlugXLRFZ92XXoTtffZ9
zzXH9QdjQbkruxBj6x5iVaBAMfV+WDYlwIe2ucZ2YE0tWqytvb7VJQlsOYqnrUhL
07M3BhdJrQ+hK2oVgDHIR/UGr9StU4FG+tkzq2o2F8ozjHFpVRy1A/dOivdu1OlL
i6CQa6vJB5zo8PDHa1QDXFuHLwRklh/NEiyLTP1kPYvR3E2e7FDn/DQ6NmG20AtQ
OTpRkls8W5f6tWNHHGfA/wtp03vJFyCyGc64BsgSqgx11uZmSSv53vtKlhNCeMzp
1rZX5VyAl8ZOfQMDRQPNHsdeLvUkN9WN2Aw6AAr2EHjiZ73uKDmUhqU6p8zyeuwP
D7MjepVQQYRfpoDBO1feobAez3jIKIByiG3UbtgKOY4W5Dd7EEub77yThxaJkhSs
vSirFjN6FXlIwRMMeRIj9mQifNBGIHxjAnI7mXQtOVZD31Q2kMB8mYVUP/og6kqp
d9+wpNV2AaxeRBiL5dBp/JAVSvFFWlZcGb6yi8tYPJd4T8xK81QRqAUiyQy8ok5n
4iW6zjaPtteqk1rtfLbfmwCGRZvQUeyqzy6FIhxDFGl46S8Ia+PVFaDk1sxaOBjp
cFv7xrvk9Z8ZI6ZC61CEq2ozR43OluayEL6OMfEnjL6ns9LCzx3c817EjS5QuGya
BenoBfK7mYgW0R+U0mLpaUDnZ5MMckxVEjcuG5FG8VW6OrFny5B0U0SC4yZCGn1o
OAeDe+bAmYawFlJGKXeOvAmEtVRE+ddA+7zrUfH85rKIZ5MoHlDSk9ugZCXkVwO9
BbmHxsN87Dbxp2XawO8Ol3NZhPkHNPOT2rjR2bekmNkEa0eAUWkTD1JIrm7ZDZiz
OIQD0/2Ddfjm4yb29Nf3Il1tXTQWPWVRbnumm7OamN4Cd2qM5AO4ucyEhUJCGIfa
lN3JkLuoNdV7k41ZSDXq9RtlAAvGenCdEFgsNOsp0RKWIYFlgLjpR85/tcfwjX2L
uS3K4SjGfUB/jCHYzHvA9XM9cd1dkm0ldeO7uAY2wQ4F342/ZD/el3r6RhJoVHQm
+FnwOjPoH/xNmgwgQk3cHv8HGEBvXBfK2wmGGVOAa74cdxQiJVlLuA/t/hXFr2qt
LTs8nTQ8ylNIcrE19PpNrckTr8pCU5JRDd53n9n3q1QyrVZxAw2jfcF3kg/bB6ZC
XsY28ppvp16jUfchln+cRwAZT96q8XnsIwH1ssIageTiQ+wkpz1fYQNc39olH3jQ
kHslUNHtYJZvA3zAZ1MDZdLM5SUc9WyF2g6BTtnRmfdj3o9vGlkUxXmVFZkonOYD
KXb6tBdbrFWO8tXf6ZjwE5B9iA3R7NcGZ+Ceh3lOQ5c/sJiFTQks1OoCSa5iFgNJ
kqdybxAXbtOqOmQqmmeTDBzeRuwDMCskT/wk3UUiqYbtxA2L/aeYDKcvsUp3gX6x
fgjqOOgphWFOuZZPK+GhLNGpmrHX9JzwsiNntLb4nGhmvrPgppt7sGPc+z48PAMm
D5qDCotD2HP1nQ0zg9QOEUEjNoAW1CU1iXskpJd67FgzWmXcAPL/Lo0FqnrUXs6T
6VTOI459CzZNbBpJal2DrynCH3pxHr+KiaKOTcAG2PK1sMcgjBUe00v2pDJBKHw7
w59LzxGwXW6XmP8ToKjQBc/cawduYl8ube1Hd5j/04f8iwMaYlYhpg1bi6a7b31L
2TM0Bcbk4xaBhSIAQBpSy/FZ0vRRI8RRc7wVYiv5apNGIYRgJFN7Ra3e3X5+QeMw
7j8QT750e03HE8srvySDxOR57p5JA94KfLIDscBhFfxO4PTR/SPpj/4poisJ1FkA
B/py/E9//edSbp85z2ih3WZvfRx1ZVy5NdY9Zhyr3pBs4GsHzSg02O3BvsA6xmzw
ZNROJjNAdzSachaJ6NW4iE3osGeeIFm5q7gZIekjWOcMO+2nsvtYM3Z9u2h7xX5A
EAuM0l9FqTPT13VXdK8Lp3ZXFn28mcaOdByHuNXbV63BmsnwsOT8UI5lxDWYtmCw
dGKQaTsN7ETK7Dguwy16mrQc2EoExzUyZoTwDkjFF9tEXCbRGl42yMO06iTxYF8C
RV7TNtACXufy+oCNGKx9Fj6CX49QUPcpS1bl/4vXiEmC7uIQSSHPRHuOav4tIpD6
tJG7OZM5iZMgR3kAJObUn+jiG+034kUugZdfirdwAMlhUZVbcalWUAhkIIi9BZ2+
ENJjy3VLx+2piodtsBfgTeJUDofQdZUsHyIXYwFUxGbuUS9JaDLge916sbhJAo1k
m83a0/HkFzb9KxcwggphL5w58OvRaJK75npRUK6ratGicuzV2hZIthZv0dMvGJVF
cRVCD9WixNDcEDxA3IPHOAstEZwRIFr31JfUbXhJbttnrMpHdZjv/5aKSC/4DkzW
afrgG1zaWsRcen/LI3i41ffa46+PfEsbhGeRjlDPUjv0FTb58qp1pJ4+Au42aakL
8tih1AHQVmU4/k5dg3vVzZI1gnpzCfrsX2QAqmSFQ507GdM/r9AvjUJYfvOebag3
LLcsrGFbH3SARkUSoMQZi/kOY8akBdq+rfud6GTr8O6exPfXB9JSrkAmolTt36mi
PvOIOmXxpZ2SkhIaMB/aQ/RscC8A5LZPbuA3rURYJnQH7ru1exiPAhPNEmFKBoLP
t133B7PkhCgWoqfQ8zOiEOUiOp/wUq4566QdRz2C7uU3omLIEHfVroIZXfJZrB1K
VaFORQrmyRSvNRQXGpPx7iU8kVymaq2KX/jpYB7B/9Hpyja61KNElk3pcn8ZR6g9
OVC8AVNMdRhAXyU/8sJGKmYQhfZF31n051I6E6zqL0ziCXfa6L9KebBWMCKtza9P
K2CqMqdKEx0SSeHzbJ4Iuwml1WLbtqbIZ60+ujpTi6kS3WungK4oc2LpifqRXY4m
y09n9XCX+KUVaQKN/0XbzbNCsB9u5spj6nnmE0Cl+FxFoEiC+IeI8x0Z1Yw6vQcG
8PXxtUyCV/rtiexU4uAiEGKpFTM20vMVF1pPfnQwf/PEwSJfwFJNo1VLQuKGzTy8
zFm2n0KalPEm90kmsbO/rhSYAg9Dl0tWtUJXLSF1+3Q+AfAzVtBerRF+QWxS+P19
23NxsT0YIMiYQQav+bFZe31QvIQt8eFPC/pu/Fn4wB8YyGCvGeaWTLf6sHPkR5Em
dqB9O6/yGnR+n7MthZNBqK8HaSjoQeNhqwP9ITpW/Tk/1T8dAF5V89JRMo8NXbBG
cbUYxbHfbRuQRWHSBlWTf867ObAZEePh0SQqzkQJE7fFnF9XsDHyVYDvW+Vwle8b
RFYG8aylBPuUUPdFjDcjgpzshJaAD+qnPcOWcEpPbEAN9/TfrnY6nmYxXYdny0Oc
KSMDx8cP6CFGHUPS/RiVPZYWk/RMJOnOBbSbu1UMdQ3viEiVWl4IDduk3K27SjcJ
LBagFdvseY8hLuqPB9zzwAzkzVrJwTOwIEI6hai8WBElk7Ui0ZrBo/rj2po3Kd0B
CX/8BwHrvyEE3i5LYMfYJTUv8IExnGZhRj56+unE/n4DI953pmHAPQkll7V/cbLZ
qjG2oBWnaoCcQTQC7o/TkshVwQSIb4ISwKMOHapUXpKLrudiChfVOdps/7TQfGci
Ki3bbTNCdVAv1JcQq8RgGc/eK1Bs+AIDc2hIirC3F/wL7rwZTksUqK90SGLXSbC5
b04QH7XVMW17tMzCS7W48FNYcMtOVeLWEFeUlZGLzTfXU243GEZK2/vFLNdcnV+j
2AyGufqHt+nkA83hDDbsSMTNW79Ixrq9kFaC61Uts8w=
`pragma protect end_protected
