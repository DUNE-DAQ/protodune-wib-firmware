// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C2kcCLEAcmdsT0ouMH8WDc7icx7eXHKQ8gsL6/WYQ0NwOG8UUKvBrjoqVf/wKbjC
pctse2M/bK/oqlQs/YCrhSc5ZywJ0+IVcQ0bRIRE80O65jTIjOIuGVPw6kX4tNu2
iNotFcPR+8LCXwF6pFLLLhru83x3OUrW1X1y3jvpQ1U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3232)
mnWKWaSb2cyzuOBPmT13EgmiyiFhkMR9TS9bMwz+HB2xIkcxSH0aAEskIOPERSl4
ypGNfXmqalMpvLRUJMGKYuMWEq1q+zncu73WTLVC9gbzwgOEE/4PURgnONXqGh3W
YDLEW/X2WEuN1wveUYqZVXffcVpG2J8ThZmwZziu/pWD+bBGmOrxhwpq3sLtKsb/
I+bdxrj8LtO7OopQX0zu5p80RvoZMn3QS2mqpe5cXwiUPQRUu6QmMssxVzXDCw0H
WmWGfWCf7IFDP8Z6uryOVhispuo7CIbbrTgUT01ps3dJvMRwqZj2pLjR1P8B7nyV
tYn+YwIlBEPijmggqRzzLW3ugpVM8VLbq4wdMz5zkUCIKr0cVnBz64HupXQ7yN+g
HjUFtZnQGY/KIAreICAwYCzXaoviuhni/UMsBojC1WfZ2z2SVgY9k8osc1/tv4qz
UjHsa6m/92Vuc74GpQ9sN2ndZsK0m+y7NtYpvCC5X1ftladJ5/GvfgunToAed8UA
tU0z1RBRJAsFb6fD+b51tgvrkTKA2Uw7/GkCXlVGtDepwuaYLdqw9c2h4yWu/tp5
EKEB1Hx+CeXsnBeI7z770Pppfq4KhWYTsO6JBneSsZYyePijS0nYXJnz+GEstz/Q
Vfg1CUtdOEOMRTaZ0YADJdiWsWVeWMm8VM1mHCJ+mJGyNC1N5IuRNGdVHPl8OKx4
cVxEbgW+dyGm70Kxy/E+5ghkctuHJRj2w7Npb74XdeOCXWaKAXTGNWYMexGX6Lvf
5VxtT6kbQVs/ba56++BnAVbM0Q8/FnAvVaWUoD3pmMUvSyXXP5mjQrLo3tuaZTjK
wFX/AUoLP4wKLlU6DxWZMB5GuxDT3LXVyo6bOKF3Ohe18RTNLiPr88A2wNfBpyo0
2Kx83lDCcB7KWovSt3FhFy3t1jolD3k8iQzjwfj7eAUk08y65EdGHLgBnCLVj4fD
6aW/heYR4+V+tfpkNEmb+kpZCU3KOCOPWbLQnPeJxi2UpXP8XZGXBabIFBp8sQrw
fZ8CW6LMEj4Fl1EBJJ5jrJbqeId69//8dRG4IBXewFV2jr1IR6DTavSDCX8KP1to
0g9u6rM33hO69koV764dM3fZAFJMSp4zJwtkLG/krl+jIfyAqjE2kRdkuGz24wOU
qH4BekVG7EhiweE3vtemruStv5SkCojP/KefHV6jyp7UsuUfaVmn4FkA9l4wxYgA
xJOU4UcSXgMRTEnt6iRrEnFZSg9u2aZlJPsWU1MPoWC7qnmfFVjuIg/Xl8ZshGGP
fbMuIEK1FJi9MQWRPTCNL2leAskWyXlQljmVaMwaySbH1LtysNs51ohvq3xjyh7J
6Dcj6rZDTyiQR7V7hZ78QXoYSQZJT1QEN5N3nPuQs6wkUzao1r5kmhs0ya1jEEs7
/XrGT8y9t8DPI44Seqi4yh5RM9T8lSmimfdox6cOv8SihygmkZ07Z1nrE8CeQ9dL
zHIrq40cX66lEunGk0r/rwosgApz6dfKbSiI6jc5wYf+X5/nTuwPgVrjHRPJCYl1
WGRi5z1cUkPPaRfdjBt+w3VV8EM1CuWIphkjK+efYpeFCu2UTVRjafQzbnrELdnP
y+ZSnEhUboSLDBoTciioXdyzJU7QbEWvZEtj9VxyHYlHeKF61aV/mxpW5IqDMHVY
My8I7iGUv7gH1pbC6ROx9NQ7OrELr7AHHWDPrxbgDT0nOtZucnyRte6JnQhl2Qho
crmiIgOy9DAZxO1CO0C37PfCa2lG+pGummgNaRJC7nqtnantBsr0C9CxTf2c4L0C
vA0FIR/v5f3oNCqcJoEs8GA/KcEBBXdhahJl9DwWJrHAsmuqihEvuUjySZLP2kMe
TEXiCjMesKt7ys8jtkvzx11vrzuD7HW3qsdHxOiJW8QEIeIkZGXZ+aW1f0+gd+kQ
/vWOud4j3lCfFoeSTm4p/6zjBtuRvvJfTf/taD5XrK6SKdnDBAkFAkMFb8UR802Y
iqVsMcxotOCp62zE/yTvZExksd1xO6b0ammF1M4aMXFSnTlUywx0WJpzTdwzhi7e
pHpxJ6pwBSaQNggRoGEgO9eaqz6eOihjGhaJQGxWeKjKLiV7ggynHYdYYSt3F7GA
K1pJ04JmBdN6Vj1IANVwNulfHktyU7hoPOtLPAF7iJr64lSt/RbnbAWPeWjeLcnn
WqZbsLkxl1k26FQZEcX3hXDmocCIU+voRaZeknx6+iMi0kTnR+XriQ7mxQD+VY/x
ITXHE7dqt/yNJJLtAqQOV8NzkMLKAnHhQ8HIMuvJS6eLt0yfgVAPrNtJnAkAA9FM
rldCBCAtrJyIl0KxS7Y1j5Z1D0JzjolfcrPVBS7obNWoYhC46A3HdYJ32o/1O8Dj
VLwYuGM11wRzrAu4+yfgtptKeY79PuJz8NzxRSzcYC1yOCvL1UnBeFKkzLewLTis
j+L+tCD81wBgk4E7Uubn4Oe4TsU4jcyepR6HfdM39b5tzt+cZQNoV1NjsW2Upt3G
Tgq0pVZTmbFV86hpKINV592mrgQnJGnJeQV+ZN5KjaO6Z0/jJDltcfLSmy3/dl3Y
DyZJN2QNyxoni3O9VXvRJ7MQV9fYl/t4erk/fOlSojgFAq/RJSMQCoUG/NcVNMQc
9+k+pXgcj28g+Hz3dolJZ8InVlh3lq8pr1SGoreceUi3pMLqzweeW7PmIK7aLoy2
tIbJBYqGKa3Gn7GLDJt7ALgT5NZsW3tILY7dvPvGyBypQHlyoF+HR4zhN/wq53gh
ZdHqzGKxU5zUdRtr5AfzQ8fa1pdBW3j3huvetsGITsRSIGFa2GXJlKP3KugOXCyX
+lMaFG9V5WTlbQPT5FML5ED51WpaYAqCtCz8g+7MQ/EXQlX9kDqD3yWDopuzLB1K
DIuaderueo5oMkIhhlDXeDXlZ8swHCd+ienAxmcd1aa+/h6dVYSftGh5reVpKBqb
7bDBeljW3Rcg/mS9wdrZK1634t8cXsm6/2WHIMrFrkwOe6kU/84dQZIQtp1bhy3B
c2XdKLhqXCJ/c6bNVq78BHDK/p8h8CAmMuR1ulkC8yaRW96a5I+uFEiggPLJTkG1
k384dUus7uZzuhgw6smmVp39NVO8FTL4BUWczTEj/ZfhGQp+lgKyciNyexw5eou2
NN3vTmgL8B85gWW8A1m9ufm+JWpz6tpBngvwTz5lK7gznM1rcuu0A8PtDzCVP1Yc
MhzM2ydR6nvFIFZHW4T7TNwW2tHCediD018KyOFbSy1iOsZN0TQVltaXI7OB14HM
eEN2zbtI1+Xv04KSrn6UPx5lxqY+ZClVNyrqsqL8vEX4oIsyVh24xY88pdjo9XtL
CSP28IsOK/BvJMGi2sKgXmMEmnOHvm1wEMQNUe90wE5Q2U4ypBwhGn11SXkD37WA
S6/32/CrX2jsT04w3MK4VEczV0XfBeHoClHbUxOPR7Jb2rknFFicYXBX8S4lFYAL
9ZxwEOEcvAXEIHGPnjLeLUXbtDkmIxFbnupimQQB1vSXdwwSH1DYbe/6a1Vwjsef
IW9DAOyy7MxoK8xRdDfDeUYD8efQ9Hfnjk1w7bPrRn5gGyaJtchrhDTfOCugEAvd
mc6v2UCJ+gu+UgBk5bJoIu/dTJv/h+Ce3rcHDhye5Q8uCXz/CHIOK8qmMfci+uZ+
xdEL6pdKrzYw1ndj2rK/c1lwsl5TH21+BIaofFvNMn1XSYT0C5YSbc9WLIDnHn8Z
UNbQzlKLuxzPQkh2jFQ9mRHHozE+3OUVFm0Ybs76u11quZq2BW5g4lLWGUi9e1/k
kGRlKc5xh/2EjpeFlrA43C4g1VUHKctr1iYyE+N5MW8tZcuGp7rW6aA4ighuCAvG
KHj1InzeaPhU2TuRa1lD3P8CbKrryiZuZVZ5WHSTcTubkoAznWUl3Aaw0LgtZLwo
RWl+7B/FfqN5qjXeVnmKE2XPTSPv53ThtEM4rpiP7K4bRM0tBvlAnOIMKu0Vvctv
mOQ61Ho6coAMNTiUvkafozw0M0Wdou2YHG6ROYiK+xewUDpK4dgui/XfQhDe9ck8
F6aQTBQERCJm7VWMh8Vsn5IQ48eqDyPdjdazOQK9m6SFOMlnRv2N8RdIwTHp+SGG
BxXddatXDkfxiU8vqwks/IMZyAAVRP+VsMnzBCMVmcKr5NTUg1JwNLVJI6SnnCKw
X4hnN3uDFV0yOL97tS9vFixNVPNqAyLxyZbYpjnmMX55nWX9bS4D5Kzuq1sBBtgP
XjOa14feqUwV7X/gfBAhf81mhPf7ApNkXEOGm0R+qml8ClL9Uur+gFVHYAESNDaU
ePZKbMgd6V2fOHPb4jnLFw==
`pragma protect end_protected
