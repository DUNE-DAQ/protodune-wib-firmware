// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mOy8C1QfPU+uhpj97isccwndjNiLz3EoA6h4HkTYR5CIFL7bk6593vmKmgntDez0
VAI2dhP5eeUzziqjHa+txIgBdpXkPwUYNtkUSQwKou/7yINkcYpCRjSO2wK7Jw1a
NcNCSys16DDJtEy1+DW9MCXB+yH9QohDULunxByG188=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 174144)
QRQStJd1+MuVhD0HzxcBqfYB4RmSQXXqjpSD+B6jH+xlrxZulErl7hr+fqTerBt2
uATA2nfM/+lRoIRnkMpX7GD7nX6z6CYfDwA3u73jjv4QfRow49jToAJLlz3Hj3Yn
hP6T2YE5Ibp0lCFhprnaQf1yAAiokDfgsd2g1zCWeik43puQKa2VuOkOg5Gftkvw
4JYDPUUM8Vf0eTR2HE+WNJEtQxBziwdXkjKVp3tyqPcEDWdZW1NgCMtTZAGtBiAT
R8EzWsYdaaaUzMnJMN+/Sf2kjRpaDdNFLt+e01TVh8Gflg+QLiUFMIt8frya7mg+
eLjSh0X5csNm+BzOmHqyFUjezXGVmgLn5wOVBYCpM9qpdbX+pJ56qhBq4E5FGwHx
T3V/VgNbCT+CmuopsqO7P5Ya0tnntAJJ2ZymMpBlOzxg9NNayQKulbM6a+JGCFCE
wtCHV4/MKkMj8YDl8eb2aNhC4W111SwznXlQZv7WREJJbIwXPQ2WZPD3QE0xnCpp
4XGvwfXxwBOp0UI50NY1/AfCN3Rw7FLTz5OSNZtwWi5MkgsSGn9yJrmRl5FKucod
ZDAuDdciGcRjzBPMcxNRuAxMsJt93eB2xu9A5MuFD717z2QySTbQ8hrV5AigQgbD
Qufy8nHipqznFLsqDlp456kEmXb/j7aP3RQhAEZ+jV/FWoqKDj1haDU5YGqK0NWM
YZzE//+JvmKpKDfbdEmRZkwOMqFf6EKzSSNH8XRyEcTyBfgqoefQNZGSzACD9dDx
VRi09vady0bqanNyVSnb1lksXIyUh2bnMzqBLs5oFLd+KjBiEd2XXrQ2ngqSh0TC
QypBugVegZ0lqMJ3FizMC0Y9a+yZ6D/UtuZGkF/e24OIZ1jDAxIX+1Hv8cspKWDK
LQOwyOF6QG/c5KA8cIiLF1FgL0FDJb0npIoIg+qB1eut3hCE54NXe4Sm75OI4ahJ
yCEWtIkAu0GY5FmKKJamDGEEXyf0K/ND3gJfWYDz0JcPmrdWYzXAigHwNM+lS65D
5wO0ZQwaJ+wjs1Yggta3BM71vVobRQvMfOwbXpPHiYowBMxvE78gqiwU9rJuN1+b
cMMafQjtOyBdmz/7vPQrdr/JKi3O5HUnAe3x92YIkqHMzj5oEaOANCCicU688ql/
Osp/7mrZ8xhFqM1/J3RWCCpMkuNnksGqcgG3Ah+uqHisGbCYAQ+R8fAJClQ8ihqv
RMcRjmDcocp+8aGn+DGDomGA2VLV/7VANlNtv5dMXbjLgLV6JnlvTuDvVZZ6UyiD
lF3u5yHcAKeySuwjtCQSUZWiM6pSn1r5QXpUGHOg9Tf5ziySrBeLNwTwUF1uJgLf
yd85EEBiJ7u2kPNohAQHM4q/gsdeKt9w3bHNU9JcIkJJuEQAFcqQ8sqL9FH4LkTT
210OdHQgm9ShpoURUry1flgAOd3kxe1YM+x4LeuOsAhrTLZJwV3VjL4pSB+UR25i
6xbKER8I3YqRYAMVfTf3eOQAw5gqO2KPx2f0wCh8h6TtUieVh671hfOMrXBMp/zB
kVRQidXCP38n188YfyAJPlN7dz8FaDTqdEtU+Vrew91XReU7OL2B1AYtKBYeFiRB
yjSR21gPJgBJU9G9z8GI6Z2myJty5/H/gCHxWKpDa+bzmh7U3aPgXtwM9uvBQXhu
hPDbhWf+GmO2Hyz5S9YWtIaBMn3VhnRrEZQ+WyK065SAzUdmahgcp7tf6DMjeIIw
m8iWurt0Bc4rvypOmHYBDAfWW/If5lGR0d6Remrj48alNswI1zI/EZTIw1mePtaf
GqZDW5zyKqpIL9oAF/6CIDNDKiN9QZckCNX7hiCky+R5zxvJp0x/uoee7bOGV7tE
gXiez1CEC/d5At+w8aE+EGcVMU82fQcihi1r5Rq5S7wUDyazjkRwVb7HGJqstvKg
yRv5YsomjfR2o9lUnViA7SEpksc4ByTRvWdvDdsq6P6emJnbQSfU2c+bj6pZnOFK
MoVVB8GjlHE5jSDJ5klUAt5DbVXadQL+lo4S9XFkZUvXoEVVLzaDp82QuSjNeDA/
Cp92Bm4rLqq6i+jBc5rDnJLSbd7faW8wM12Rtaet1Zd1GG4dC2QOd/9UZT+EJYnf
L5L9UNM7Wp4gd9PW0jiOXhEnbxOXBoStHHUIW5kbfXkIpZ76V7rFZDA4lMP+Tk9z
Z5E9ORmEi0dWwbuhsWhskkEW/8c08ARpL/7MVNo249T+pqJE37A1Cwi7bvBSTrjv
lHcxqImYoFsZyOHKYFk9lsZ6J7hj4U2ANxuH022/XUF+T/+AY1+GjYYWtQM3j3RF
zyHC8FgXtwiIUgalcTfIDx9AFiU7X0ZkecQ3jrNxdq4u5Puda4qSnUVCHUELIFwr
3VH1WYEF2xOBWYMnVkg1CUroURPV9BR+/t4Tsky7htZXoLi4cP66fSZmQlGXKmpp
qv+O9h59rLA16WLRo6If+mEJOtLnT0uBZY4uquqInhZuKn9G6mhyLWqlgFiId9pH
M9Ci/2ivBHjKxlnom02veVIaqqKU1TSZ/viNrIN9nCFnZL7SwoYQK1OWkHgUbHKG
znp6c7rAaCvmNJjbjzuy67ntsoQWc+AD7DT77vqW6wLm66xiDBU+1LSlCRaOzFb1
22saZZjWGlXHFvy8766uXxP1On+JxuHqkm9u+9egUg93topmrp/QmNZI5cOD8mYu
EEkh7q03Uws8Qrv18b7a7ZM5+YChUFnDWLGTQCurMoe8KFdsoGEefV7hJ1EJrzEw
Sdgg9IjspMaB6M3sJEMksN4UvoL26lX0Jg5AuDWdzkwgvO3wVKyMN3sZo7ZknDfT
AoCH+7Kn1tkRTqNPX076i2DgAn5fHWjdj5tqD2+hd/dsJOmxScogPLkiU56X6YC2
t9LbEV6UKTgPFepCx7rEf+GUSYrweWRWFwJZQDokXkpEED0nEpO+E2+Sks2F4Ikl
17tl9Lsn0PVOccCYzg7eQD1wwUyuiYQqBQbKNIk4W0vJu8lNuK60c/NngrG0Ul7Z
I4fZlMH9vhAf1gmrR0f9PvuvAhiB5MYfoeV7z9hUTNS3uxy9aG7Bbz5HFtS8/YO3
/aEOifO8pfo0fnhf/LPiiUlVdbEjPcWBTO+sCgj/LVYkbNT3P7dLE3cANy2UFLs8
//A2LRwKxpeJKcjXe36hUu3kASQcf6TvIUt91PLJf1wa5P/ARGg8fy3HLiMtjbOf
M2ucvrLdDHCm8uQ7CAU5ETSuT4utNeSTrCr/VY3ncuG7XJnNd2G9gN6S04sBtERT
/5lSwV0i90+iBlG+Y+xNZ5OrpdsPSqxKu56HU9E1kKoYBuaDcxbgnVd9EkvUUsHO
hinqEw74Z1wtjK+DC+UBKJgL7xvF4aToOyXUoqzv0gFAVpEmtLyemafOHfI+f3HT
pCf4VEYmKKuiYK3zdeetQaeqHoXgkDfL2LmOhfWG9u01qLaWWo+xKuxyTfM38nOj
lWeVfVT5ug+JrdGPqi1ondvuNpLxpAq3KZu4dNSqahPbEZXTYQmI0H0gyRa8QgMJ
GheSbcdPWPVQ6/Ogmp5YgLIXWgiwBwUrUnBFs893VH9Zs+0RX6LDV9sSgpY6JfD1
bx6PstJJsny7z7IyrNbexZjHHEbv27M//l6Q2SVZyIUDzxMMz2iue7VY9UfCOYZJ
z8fU2KT9st8Z1I3s401ovexsSwIK7nlPS3OnmZMphwXXbHhgbG6ofJLi+2tjPGpl
rkGIeTKBCYzT1CLHg0k+auJKikkyrzJPLEU0EAiW47/ugzwvrkLHbTKB2od5wLt2
FHJVr4M+tbCNh1iamKYbN2HKHzNuw739e0uBTDJGn94dVcsO5YPPlmTYkKJF00qB
ktojuOZg8DDLl1NCKvdDFwBu0iYRHhxqrPlGghrptgcQdPoNv8/7Gwhsg3WiiBZd
lrAmD3i0c8RGgskdg5q0w4BpUZSyIVR/He/T2vovhUCf1TLCQy7670SDuqksNIFX
1fmooCEQSq6oNK7v42/4ssmmxc+3FQx/HxBfa6SDpBUIKImZujiobOt5uxaZWGPN
Pilwgzig2YMM4CJvegKO/2bnqvQYkUN0aAIQcqNQ4aoB2TqLE9J9TdNuwqboDZgY
kcrDE695ajEA5iR+B3ogaArHVRwBwHLKhNsRfIYQcbQLgNUlPEw5VDvV0IMj8DC+
ITlbterUfNxlU9LtkXpDCyJWyoctgylVTD8t4HSCQFKfN/4IrHCCJCD8TdTRjLqo
FkhC692NaVIzTHUNvVyS4olMwd7Ud/uvs5EKA/iQ2Sr2vJzIvmSNUfX0kpeMVlnN
+205x0hd0A+UMIEzeUDiaDPZHE27fytjGzycwsTa+dCYT7KtsJZabwB0VEQThbRs
cPYAwxFaKGwlapFXpkkUj0vlAwVB7KNOkWXsmq8cCkv+rhCe1H6MInLtSWiLiUfd
cIi81e/Lz9YgbSZWvoy8ML/Teg+75rz3mxYmHw0FBx6vHIGBuUHHhJyv97Lj5zKK
6SAmak108XyESOt37La9sfiz3UPxmMfJ3ulFUkLcjEF0vVymIZc9ZGkwyxhdgoPl
XcYtW+YYKB153MnnhrgHZ2jJpo5k7+HdU2fNgzfm4q80AONTWrgW/RodspznFUTF
47U5rMh7BkJYvxqU8dHbmMcN+9k6Kcz40KRtecJmRLxDQB18G3oXvngNKLSPlags
i208C0N3kl66n0Naz8hMKV9JX1nKdFz/7DCzgytAhxHvbjsUzhAcWWyERaYkdHPH
qkJDTkEkdfmxmrpnVD7WNnl37Xrd59JcLFZ+Iypiu8Q+3iJSRDkUQyfm+fb/jvr/
oda2dfpEhGEyZWOLy8PHYxfE0zVrAIaU2IKvjm3Cn0cSeMpO8/3g2QB64G+3oNMR
ubSTJb8XzHprvlT2iLB8jaP9KgCyFX6TkWJjPFmglBn0Bd50E7a15fpFmoLJ4+ZR
BiYp1Yq6hHQ3RkNyOJoOkJEK6T26wA2ZbWjb+Rw+xKNhCf9iN354ONZRTy7fRmta
W4MNFbp2AEhXOzVrM0If44o9AohCEgGVkPtCXd/IIu1aARUPu7pEcF3fYG6gMO99
N3xFjSQ/8SfeNNuzNBwdbP2xcd6zMSpHe/rCDSvObADeoUmrQs+4nw0dT5RMdkkY
kI2z4F/mzk53LWcAYSkMCMZ9Ep6WrwjuK9LpvzN75gv2HSX8l9YKBZOqpol5qwow
bv77QzjzSsqQ1Zux6Rqp47PKS0Y/V6HDy0wkYMJNrvlFZYupcZEFHsExxOSb5xpC
lEFZDliSx8xvWkHxYIForZJAny+HVZC1w2qzVFhqLUHNiXCoW88dWLyQpMFsSfPc
Y0CTqTimvCfka04jp3FRj23knWhKzMwtyIdvnLt7lqNWXS1hR+zsOV7dMgAAbsUX
5kvIPJOYcUE+CwvZrxfPL+a2FozqOzgTsCWlQjwOxZad9BcORQFFh85j57rCWvwR
HQhJZQO9AGdQxTpC6+XCypYb7DTn5TzTlO1WT0Qirrh5NwhgajZ12iS09hCJ07gR
ci8AG2qwP5veW+fjVQ46Juee0xXl3771Jfw1L/kif9WSC8rL5lzpxnxHLTjKfyBQ
ued2Lp8go31/xqcNzfpcZNKKGuI+qWn3lmc3CRf0KKT7vTzjYeDjuHjh/YNMj34H
S0hhT1Y7GKPJ8Xg68HvYsdS/XQ4H7CPC9iKi4FxkPomFlypqz47alWvNcU8kaEZC
kJzghMRqbH8KrPxj6RFffVG2AcD7IwiJBeWtpo4A74kdEm3GO+GX6sU8VFTXFNst
ZWLlgV8YvDYn6SxND7l43nu0lBxI0Z+WO08ausCh/6qfoxudV13SZp/Foo3A2JMu
SH6UsRI5O1GgniO7S+vVp+KXQrYtVhDA0y0YQDjmB5q9+nW44wFLui1V/icHwuiH
znSkpf30h5kTU35J/q4bTjIpXdooHSHZcKkLjDEG8E4SGc9NAXx+lPrbN8BirQxQ
i9/gs37TFSPBVVaILiaXMP62/BaN+xeO7QQtafjQ+Ft/aJJE1fVYyjdtdWfLD128
n1zQ/x+rooG4zCFx50LdI33fDHMtY/iOSStWn62H8Rb32q0TsmQgJwTQQ3Tt4JQ/
xgEW3MfGE9WIK/BH0vDVTkrhe50E9EqRmnVbK0r4Mhbd38FFFqLf5mMB9kbo583A
r6zSf8dV/KYrO9LmMLnYpEMTfwGrJ7C0Vr7+nBSzcXVXLHKPf8spLniyUnLmPl4a
7MCOzHBPttAB8hGoYDmBOc2snb8uf96ntkZUyZGis180gTWIgWvMJkyI1OLPMQSu
G1CQozJWvHarTRDygYmTRsT5RmzTgxy5PrR90bUlNSN2gxH5FfDuQvUqKJ21rwTm
aj+qLmCULfNfqPiybytkgU7d/OHD9pUYk4cFTACaaY5cpdtZxzB6W/Y8uS+5lI3p
RdHc692cgSz/fp91xgVzctRYaTbx4pQRe3n7GGrLJu9q6JntgzjWT3OZnzD5B80m
6oXgZf4qvR/iZpHV8I+7jIp3BjWy8AlIaL4s1HDYC9iylmYDXqh/LMMWQ8pixaKp
aedOfiCq3cXZtI68qbCo+1vTRNFjJ0V6a/F0GDiIq57nUeTESXfMNezym8axYtUa
gDclcj4ssl70jn9S4a+1+OcH0FepErNKtlL4NpapQV9PFAGk2MBnB2kbZz/orCnw
SW8vEP1JVDfU+/dt77T88V3a1AVfyE4in5nL5IC0Qhqs2LBZ2V9zQ/a4sYHOjKB0
GHBiRLkzY5wCXOwMeyC25cKaMRBN7nxaaIcpE4y/IGzMxC4KpYwd5q5tsxWXIqs5
duHzWIzza0fj307BKrru958kMnHA1+tper98yeGpj/nFRu5HkzMc09ZWrlfNMB4g
QSMfgdQQDS5U1qcELILmZUK9n/M3C5QAakE3vSi4BOR9mBc92l7pZVZeJdaXDazY
f17dDDU6i29HdtIviHpGoeOH6vY3FDr2eNl3vZqhZotWoJLezrt5uJRI74yBYNmU
LYIhxrsQAcP5tepP/rgMViYijnfjgON11fzECN/b4SUEy2ZPWzuMfpT8N328pNxV
3xacF1tWwme2AZ9En1rkVlNC/ofUKH/MMv8MIFjB6Gy2QTgllsgtUnwM9SlBHJb8
mg474613jwXutbJSw8k8QjLcW9dG8kvhukM94P1D2M4Ltau4el8wRWUJ6rPC70Jx
L37W+mw+BgrJTXi+MV285HbBB2biXM32ymV+ZOFMo43TB2/Aamo+968nVFLsnT37
HMVgTWRwq3NHBQgkxS9/ByDRc1SYFEzyWc/rXYUWowz6wdcG5JcQuScQI+I4kRBd
P+O2hySKVYqRS6LCxMgzdwbQg90romsI1yh/iWfuKrCFXWkFpUQRLEkllg4cIgho
Aq3TPo75SHmUJBWc/+aGhht62IFCQ5cCmLvzJg5cITdswj7anV5tmLBMboHYLe12
WoR97vK4ihZ9ymGbaHT8jsAAEPie5b5VqiIWsyaHuRF5ho5DjtiZvBi6t+CHqUaq
dtNeSEbxhVScMmUZugipX0ubAf6pQ4BKVMhpnbLyeG7m261VxNWRNJ2ZxUhdO7nT
RGkeXOI2HMuBtEyJ61NtlLvH83qXt1x2vevkwO3ZTtP1/p5uFejTuP7ymp2jYkJl
A+4N+Eup5YOq4hveAf0enXiPyE9leO9WQqfF2mj+0pmm1Jvc1+FjohjcSl0CvbHM
JzVMiLnLZdllmNb21RNFICTYe0fxyEfXzojiEJJ8NaP3OvcJ8YYP3FVSAgkITqR3
Xt/4cc/NQC83ZSjm/dNxiq25n7q53CCU2jBIL6xjHK027ZWOZnEVRUnuhYuLGP5t
tswmEoWteSaO8JFlKiVfNKqbRJ8gR/ZCnpbl3BSQp1QpWoevD30H+SS+fE1362mV
8oLs1nPswSeAZCXR1E86Ig3F3JNbHX1NGudzxihFeWyGldv39QWPxZKKL0mrTL7k
uK+Pp9MLiHoYy3KPsv4cX+SGz8OZA5hkEaAQnynRZtGJXJPd6HGrQfPqv0wiH+cl
Env+f+7xSJsD206lL9vvgllT8bmZ/C1j9ON8ID8f9B738WmQFxNerk+acHcb5a4p
LYOUk20WrItk6SRGvkoSUaYqlDdePDhsSfD80yWQ5hx16sELMV1/AJn/tic7oBXm
aCXlZOa+uFZXC1qN4xUZ2obzdSGhXR8fSWmpQfmHWm3aO6h+iq8ibRBvB2ZaDJAp
hfFvRwAquvhpnXiza3592O8E4+UR4E3cqqt68t2Dg98tBNh3BPpzOyRiJVXoLF2J
ImIp6DpREg2Aqp5rFzqJFWhFdVh5AArriMDVf1EjY75mjYkv7kfuRB7yLhQQtoCW
MlZeVIRnx5JXlJMmMWyHOvCpzOqm96ruK6MFSnf8lAc9G0yXqLMXW2/bErCmQleH
8A2FMSHY/kGiFHsqZ8+funpAaezRM9UfjUxOgvp17RIwB1xbQsBMeXsNrGOr7TRL
7mHxDuS4TofJiS3yM5m04+/g3o5g+fQYl7eJK5rmyD+Ebqmsuoidb4YQVKczidYh
dOhc5EadGOlVLV9VjagJNr1p6PzAeUPmSFmZcXfWQ+cHifhkzsKTQRNISDtYYpOA
SMSaPWrCMJhOfkq59Xu+6q6SF2BOfthC8jvLDSHmgvzITg9hlJzkNJ/jhoVmNAVd
cgsDwso3gVtHVC8lKG66VgVGYSekz/cQKJNuYvbU2i9rEFvHBCLYiArxCITA6mvA
KW1nLRy6Lr4h7j2Zvl89Vx/wD9gsuYB6eQKNHnd+dJ7aoBsNGFkgM74aHlFB/dit
f3AcOBZhJBJbVv9w/QpIyWlhkgjjktXcKYtZROADHqZRd0RtCItBrxFM94MA99UG
GLtjO4jEp5k2+MD4rFcDPpKhSwDSQzsaKLMg/kAIGiQolojrzC1+Sl1Zf23R9o8p
q23y5+UuyESIG2okDTQxJ7ODCwLfoJ5nAHPcSyP85/978Trzjy2W6qCwwP4Jx3ZU
ecJvk1SoYpzAnsbd1tY+ks4ViCm8fOeqgwP0dsBbrsuKHzegEU5mZ0FzNNICwpMo
vrKjcMj0zqQF7VrOWHcUMlumCvNThvFizeeftiAqz9nFSIPVBD63EA7dSZJleCM4
i5MlQMNKImxR0/LCM1JXwWTWJFWf7DqEpLh8X5mV9bQuLOVbwJ9Xn6uWsJkD7kQo
H0DAr01oHp980h6ztIeyBMi8I96zehV3XuFmSGJHGKgW5cZ4pxshfbqb5gOwygLb
/JX4FdLT1m3xhOVvV4Cm7CEEjbh5adtsSsQ0dp8+cdf8x1ShhiMovWdfArFZGDjc
BHmvWZECnCdrPMiAaK0bFV/DXy1I8mNFTna0R9sXjoV5iqN50YBogBxvWoa8xZgx
v8K9E5M0ZhxAIRgLww8Od30amt99//HIWPMf47Zb+ULem+bkOD/baUKRu9IEovUl
sXZhvYu2Ukg+SHcXTYQPPsNy6opsbCO3O7nbVS1MzUwrjilzA7+vMrh6XQxfPWRG
7jJmu0ZY2aPD43PaAGIk1rIpDeMRxeHCnOoW8zvgtLm/XvdoYK1gJaHj1rgdCMUu
TK/822rORsLmiTp7HPIF1wCK/5spJAw4b50RDomJo8N6s/iZf4YDRwoWMRjSalKp
OcQ/lJVXJ3l+CWLQRvfwrpnHsHwrujVD89BuWxtW2s3KXeXPD8eT8EVPcSDTUkVU
sxAql0Hot79M4jAAL3aXYVAvL//heJ6o+o/9/hoTs9Bmi6mIcJ/YVTxuB6nClEwn
j5G92IERD5YWrr7ocIVbs3JZauSqOAeXkqA6xLlRC7cEERLs19++xTZ/IVayD/Zy
Ulj66SJL2b4YkQzIN5xHXqpizD62QTOGVxikGmgrY04cxX3G5FP1X1RvVtaw1y1K
A8XU+JIyUZrvj7iQbYDCzy2cdj5323XhdkOF1bNKn3tfqXuP6aTLNb0zdliuoAhm
RM7xRftcbNDjcMd25xA+/cCXd+WFvfU+rkCMXcRo6C2Cupl1PUoMEqtc9fNhWBnC
+eXhm5Bn6ikotuyUdphZOXD75PBxnj6FVRmWotVCdDxtS+OP0jq68bu8HhDwHd8d
NLyJVvV1RleqttF/dvc+qsXM4oeZc97pBgTudvnvWiwczZCzhMKuYDh3zNxWXAya
TPkmP56fYQJMb7Ibjr8hEaPY7tx6+i0W5be8OIeMM9lmm7Z91jCuQHC35mTOWNzS
c7bJ5YVTmxvqY4UlcUW6/QRRQdFejiZaQ8NCoWSQXA33ENaLQV+BlLWu/fBYiTNU
kVsYo1NoicbW2AlXyjJUXdelgPimHG/pq4+XlPvTXjgI5x3TtujLW+86zvRzDs07
tcYiVsypdiSv3tV/z4TqvPbi0YkxE+QVH6SLqhZXcy6ppvIDaNuf/i9amXhMiB+a
pyjBD/JfRADTRre+R0WD3GvAauRJ2MEM5JVyTbdZr+3akIinsNCa9dy6b2MP0xBi
vHqpReqF+ben6ycuO1l2cs3z1TNP8heXX5ln53i8Ihs53R/WAmzCJmyMbCkzXxZb
u2ZjO0JDGfiorRdie7svE62wEiFuFhq5ewwArjc4EiGKP07n+YRIJ1wCPz/uRqwR
fBOb0rnIowvzOWUtIUnQIfrXE9ST7u980kfZ63Hfp5fyIimvVkqZ5zkfggFxM8zI
0UPb0aoi5L71DnBTLollLCfdhlrj0f8jZJrkOjWfkO1jOEmPOB9nS/ex2XeAPhc8
xMVrk09n6CetqvshwsB2ma9OlVCbj3MNLl0tI681852Mj3XGUjC/N4eMTEZXzw0D
fD0el8BUjWAcMr+2vVwR2NTWSOA/m2e8cyYMA5kyrie7rK5qmhMasB/pDVAc8uQo
jIP/Igi0TYTtEyy98+CKG6tnBf2ZmYMxl9TyZIFlevYqCRXHKla31ajL3JGNcTlB
K4/xm1Ww6tecg1zw64RAT+EI3zjawevvroGnWnbwAhZ922cqWOcYz9ody8vthRWI
ra4P52vXptJj1bCUAv6V4aYk0KtTyu55/fIYCGFN8A6dRfxXbo8bPv9WpIdh8zmL
TISRFxtLyyVtjFujd2E9y+KJ7yLIL41oh2ZvrCGaI77B3IgKdbP1bMeabPtHsjtn
yXRXwKec/TJpoyV+izDF8bkbQQLpVJRLQiG79VCapOhCx31yGxmJYXifQlAL+b7q
kBpOcDdUp2FPFoDI9vJmnvnIu1PhZuf0W96yg52mclib+bzHJF/MO693eybDC/xW
fUhddBZPgr5J99I6T2Wl9EJiO3byWfZoAGszJfm4FM8h9YfTsUr9kvClQ6y2B1AX
54XODQENg+obPlG+dQeduIAk9R8kpG7iCSWrN04GPsWGf6vSUGvoAN9oAooQZfde
DMSD+H52BbnHm0I/az4eAFtpuP/82RtmRGLirwbMLczXthpsjlTMjkZaOGstw1Az
jrzDLBFJrJ6P/D62QaA2QifM9JmHOUs6IB15BCaxepu3FkPmygzx9tCXz1mNUKa8
ZzYDyX31F8c81+E9me8/cKpik/saKFSt1Ck0k2ZsL1wJTlBhMhyaxpxaZIiOq91a
FjAMLcvOh1MFgXKCHeA5jYvMY1XGTNXw9A5oKVqDPZh3fK/3SFJv3GTrBqdPtvGI
75hBihMbOIx9EpOjFuBVJCyKQLWdTfu3FQ1K3/jRlk42/842Ka6q7W6qKUAWuyPW
h4JCm5FWP76GEDsjYCtt9yCTkcYxSUfUhHSfC2f24sLCZeoekGBDdkRZIxssnhE2
BheLc4cJv7EZzHwA/enI6sxLPU8fGuqdAxWW5r2ZE3x0AFlDmbpppIfJ8xuWSspe
MpvfAVE0iCDr5MUDOSScGhzYW1APszfPAe0v9hTjuKI5zAP6fzKxlcqcJi+7Dbjy
4mscVUynPT1u87s47BCvY6azQCapss8JeeBrVHI4NwbdJCV8V/devCsLFNNJZs8w
OrctfdFuAM68N0Q1BDAAocPESY/I7/dap6qhS9tMe+YNuC2lN7c3NV+l2f1hhb9N
qTaRP8UuPlzBVlF2ProxIOJIzpZBIHvuSb7X/zanMMHUr6XZ6jGNHIqzk7mTFp2q
Xpf2e5hfAZY0s+JVGdK+V2usAH6mGX1TrIaLgfla2MdmKVm9OBEvRHwlucU0Ia8l
e35ZMjEDFZRZE/5VLaXbgRMzmaXExAepXfIwzVZ1h6kw/nlA8/YWnuT4eJFD3F5y
sV6VK3mumiT8HaNjyCN3hF62myP2WlpLINHAR/5uZDExeYCB6VOnULVpj307BvUP
22xXu8orAM3kCqJpNBDJj2c0j/qah2PEs4YxGVzVgfS92cPFNc8FOzMHD6GfkcCZ
wgs3sWfatajk+IDQKgrZVU2fjGSDqE4ehpKdP1iep5jOif9x7EM2RxLrSDDwBuQu
Uau3oxoY/+SutBAzcoe4mRljIS1dzAcAO04HG2E80Ks5+yICHsSiooCRMA8z/xXH
DzQnsENEittm4xWZd82azRCWag4171lzyYlcz/AH3b2xMM+eGWOK8sC5wzBjtADC
UfTnJRSN/RfB9feCnUn3vi7LaaLGLB3RbwA1yFJUdMRZCyd5AhhDaNiCNcmMrKNK
uKgQVkKRzHYiVatXGbXgmCom/kBYPnEAiUl3GMdvLxao+ZwHrZmm++Ip8GYI1qzh
yA+XVNVHm0yodn7WuVzoJknfsdi+JT6WdHmvFJxDQ/1oikvHgFfgOmdhIjFpD/cR
Bg0MPNJuBCmCRYwSef53GKb6CPKJQztkN2zx99j9wFey96EEZGugCW80WpjwFJNL
9MMaowhLIZXy7FKhiffwUpYp75A7n2Mv+TihtvBWuminB3SSTOZ/TKf15cdKeB53
7y2xooCDtZzgF4aqnW1qP3oBTyWBs9gJMyGZ+/h0Ic0z8OB9faMCPGFys/z/yBqT
6X3yahxI56rDM+8j4xKAq97LtNUDvZCqGeqTh+VN2ENdCi1E5LsFFk8/CnqISDj8
osET2Fe2MBLZ5PJaxnX+d+F+7/AODSRHYgqHFU+QKyKfYl8wyjHZ6df9Fc9FLbvk
d2wCZrcMZbVjLmMdPCoibIH3GFMTgInQfZgVjLh1NSrwXR5Sl2hm5yCKO1hyYeiS
uxuhQN/Po2PxrbJEyappEns4DY3ie5IW8CXBOxfEJJ4er2vKIfIRrNGgECGrG3hZ
TOrZm61LCcTpaBXPfmJS7gB/CciV8XtAf0EU2mWzZO/uPJi76Q+WwVG8hzmwIbWl
vKj8LHVlmFUWeOWa3FAmPFlp9COd78kWQCMEnfW7lDQTxsh4nZsqoNEYdXPQs4u7
2pYRZR1gyR4McQQwgdt2/XSML5Fc0kkNjUS0A5NZ3oc46hOL5SV6KY1iLLVg25+Z
caMs2XBZ5pQmf+5euyBnPBx8jJdknKnZvJNikqG9pn+ylZ1AuqpRJZiWRAaoxdLt
pLLlOGUqk/RsOVWcPTEGdHsSwFDYZpyv7H33x1zoLSP9TJcrpDXoodiFigDu3reJ
DjRiVgFmzjpOZCsqQEvEefTuEc6Csy8lsxYqhTHErEMrIZje57ffRskBU5F9cupc
BURBf7sqE/Q5KaV08jbPFXg1GeaCoQv47xN1FPS8Sc+RcEedf/DWEbgi5AeEidY9
+GcfwDBsULRfZxX9Qi62ENOnTHayC98jQHGinfSYb7/GK2m74J61rTCsbT9fR0Ev
/PWHuHz9AGsR4Lr9Xx1s8tu9dvWDiQEh5BP6wMi6EDIDdd+8aEz8fZowfvyvBkPk
7OvQciZT5dywOf8+RRpgghbrOHMFfet47SEsMLBbejIoKb4ALwBbsfBMXSa5VcOZ
o/PYRt4g4goHSPY5kLpcwldODindrGwXoEYqXHo8rVAJ8UWFdHkt/P8X8AkErpbk
VYEoa6orGyBXox5TDE7mNsfgKm5NA0VMUENvOp//UkGhVCzDKaxTE2ETXxfFxjWT
obA13KSn+PlDr81do2QE63sCcqM2VHUxbXBf6KqMrHxOctzh46zUqgX9jdppkxzo
JFkVP9rcEfJ+75+f5lQ5ab1yxsXDkvh00BzUjZYtRJjvru3uNQzdhov6zWDPVm2U
x57WI3HYTdxCkSve2SBL7K40jRZewmBgVW9XBk+2Sf9SC+4dsyw7FX+f2crWrMTV
Tg1Kp0QI8w2ORB5BhQu1yO340KkyGd3f+JZaWqS66XzY8AyDt+3kLvgwPUxhqFWT
fOisydvHRrFWNe/wpR3LYErXiuWnLcwBSVhsjpNK5UOs1zD4gxoWVFPtMVLFaUSa
J9qSoR7BJidrmX7BZ9nbd7JM7Hht5stlP+HA0h4t7bjoaIP4pHSju97l6pdwMj9U
X2nI6Glbcp4tVABM5kGkbnBZ+nI25iOw7Fd7NcPpNYETM/IInjxFwXWasMs1ryRC
W9wwBnRVrBdANIzWF5DCEjKYmj4gy2aQg3TrCULNtb4tKE59LuzSzgyCfO4948Xa
ktZ1QZz9V1x7Sj9wrbIG5K+X5p5sPFonsirmXYgVkJ2mr6dwA8KvmsU1oVRuR6NX
IwieoQhTyfvWklvSvDqcGF8FsUZW8Kmb4ZOSHqw0a8EQ+i6TR//kn+ym1RwhTTwi
aUckwo1RDdnOD9+YdSehqcdxFRSiBstJp7V/NF5sraXMpmTiIt+Hwssb5K99YKCD
4reqoOd1hXQ63muscisvwR6V0s+4FRckutlOx1KZuj3B2C1yj1wmYip6PFiPgJ2H
MsQRTZ4NyB3xBf2EmzvGcNrYhcWQimADqf4DPWiOtJrb+aS7WVjMZUsesjhdgesk
B3JeyqU/iNdu8HXtCs+t9Z8f+HFLWnQIZNcqZxXvlgAdC3Fza0YIUcCimllI6e56
0GdyVTlFasRy5b8qMMjkwD8UljGrvXggot1r61JzmAZQxmcPSlzdX/BqmLdVJAqJ
WrgnRRvNanONTtqyPTHwYH61Pp+1XgoQCjbAvdJiH59FgAmZRxauF2oZqMBs9oem
yve0wTCO7NGSGXZV2NuH8KO77jXFV2k0FEi1QA9bwWb+G0TdsVnSgAkDscRB6a4d
zlWbcnlcKPm/eFPToAa92RTVQGUkFwEkh8jF5ORj8hqZJbWkjWznA6lY8fhxN6v7
rIuZ26KODZK8xWlGMdu1d6T6QgbxjJKyvIILkBgG8Kzi5APHug1nnZAO+pAiEGYV
/JqWlK4Pizt96ttRcIY/Vu93p9HQj4+ncmH5zbJAE2mDp8EovwX2phAtbj8kyu9W
TV11H2UiTmGVzCal4YkEY6/jZfLw46BPBxJRxAelDG2F439IIuEh242bvWksSzAX
7MyqtSgYva18UOQOsMBgGCkCPZFxA7F6u3arDT7pWneiG4q9OCXci4TuZQDyUqaZ
7cv27zc62714s4FuBGnT5ftNn9pIRkrSFVsJFwJZuUC9eGL6jAc/pBZaV19nSeLK
KamOJYLDkWdVtQwx8RT5p0EtMPJLNaPxF+qM1GdAJaw8FoFohKfGMzYgSdIqdNge
HhEA23OmtATjfk6tBWXHG3+vBFLcq1hI0lglFeWCi7dy0pvik+oegdOsT/lv/iSb
Pw4Jd0Y0LyGohS6zYEuFXUA+y0PAwlrum5cuslxP5ULV6DIhC0rGptz0qUnbWAWq
S59lLPdbG13pvGpGOuLRlTRvxBdqpEE4T5BUv3c4HHN6AhM5wGC7x7wDr5yt07X7
y6s9QsztQ0HcyyfpSeBx+1ZT2y1GYQ0XwZ7gKX7TnfUXhp4psitAnxc+ObqV/wuk
69NiiUFFb/KR+VyBbBviP6tFFw/aTdVlyFBPDIg/7uAilGSLqQh1JbWLP4N/Nl0P
toBVdwsJGmx0BO1QWvmOam6lWvxFlTrAgz8KFiGTA2Pd4OaxHyuK5x9uuL402qw6
GaZhS7k6he+C3gDN9dWBnoBMaD8G3papdKB4KsC2B6/1LQwTUOK5Q6p4fVaftw2D
85Tuu2XLIatE/CYDa55LIgPf9VXvh/YquxKAXzRSv1pXOd07q4AyEY1gLmakjylt
5QncrBFoYS/0AS8Rm9HKnrjstCqOM2ZG6R+VLknllFi3v4PKqxTkYswo4Mm9M2El
g9BdFqYw6rIZFs5zeNKCgor+aVoAI81hGoCD0JhD5aMk2qqelgMmlkmbqPb6hlaN
K411xRBY+D6XkVVQVdQkyNplP/UrOIxv3KhZPiQeyY4Xh1Axw2JEWzXTjUhSONpM
eMYmHcZ54XSP6BgRYBwttd+LrS5IgXP8MoJHlkWt1c8BnIkjCpWMFAQU9cySPiHL
dThAvQicnnex6tAIjRe68sPf89lPHM8taHFjvk6lmiMPF/q+2Pum5W+l/BgcHfCW
JIQBbJlAiCax+stfk6BT3UPI4VLcgzXDbM05V/MEv0YgJmy+AjG18mN2bj0rkLpU
cOSdsp2Xatr1eGxwqMV7q2dMECVER29BPFVGv+vU4WqlBZDpOFOXxjVU2xhC7kBb
HYw62Wr+4dfL23GL1mFfXyShQ1f+DKrxBv+snxKonTUJ4jC0FZmQxGxFywL1QLpd
Cu6B1DTMqV2nFSgM8weIzazma0S/jYAQbZvLhTr8d+o5B2NvrtCk0wbwAg7SXfQc
iVEBG/cWOM/eCPJbY1MakO6YRX39T0kbwMbU4h8luKHUMe0HrXvIqqmsLGbD9+e2
xEbLtHKRr8qO6vsp5nvS++zyHcmj0uI5mmOzoj/YgBpFPjXlGwxqJD76pExo8Gsf
t6vt4AtB/DUWswXu1qsDTDYCMF8H/Pk5oyJCZ2N6T6yiYuqCYl6GyEi060P14Gcx
8P4KYqsqYbqd/+FGywVHKZvK4KofolwoQEJx163xAn/DdfK4kouyOEHUSTkUQpRP
5G7wn+DRCfi5+7/8BjmU75WYUw1HLvVRtb4lJqNNZlee0nuPl6ZieJGNnXzhko4c
SUrVtXlljGaJyEqJepY+VfuiKhbZrqqHE+tZWnBkIseDi5Z+uzN7KkGK6wOgjvO2
zgY6IgyMnlIfEm+Qhv/jC8DBHmu7BWXMHnsz/GGh4okd7tfyszt0wCKW87m+15rn
OjSgR7Ew+7z3JmK6tNmQl5wib3HuQfgGzIUsSn6SI1ptWrAN4m6cQC3wBYBY7oou
WeWDuG66U7fhCgWT3rFsWNiFAIbdrxNTS4X1+7MBrNv41/voC7GJwgMhNGdHlZcC
1T2uqhRWIMnaTsrGYJtZji6MveTXMqDoak9nGiTsKBqL5q80iwvbDNCM0bYhWGkZ
w4/AUg83gs24/45YRU0UN+DbSG0TUDmhYMRZ+YC8QOMjY1eaLRlw02GLpBtB5jpR
RW1Geol/5h9vIBl/61VuIDEb6kvxt4+BwyX5VBLWVa55ly0OqdABo2ta34wkrYKV
heuGqM2oggZpBQTNIMv0mYk9V5xYBtaMtwCVNVJaQ5K3GFj8Zm6mCKFFbCf+qMiq
Tbt09UqlNfgkpvgPACswk2uCTQ00wKT7ZRHIAD8uyGJE0kNKRGA58SSHniMHW322
k12QsQCTefQ4ZdAtMFCK5EFOO/Frw5I0dnJQj0NA605WKLg4WlKny36lA8ItmFiw
7Jw3CEbUTQ2w7cs+2k629rtbnLRK2LuczxMeEs4gCDcsl5eHYZUyroDdSI9EiXIn
fL5Zw5qc4iMl/4owFOs5FiyqwxUiGrfGldhcJvUnbPYEqRoZmaEQbhkDKfodqBVc
aDhLLHQ4KdbNKkxNeni9nGmlneu7qVy3y5wu8YyJwBkIUyG5F3bH+PKhnY/pdx8p
gXduXt0T7oLgYY27ou4LqhjUptyVR3RmmsF30mFKITUc8LDy0ngfZUj+2wZ+oFe3
EkxFy3HNlH839vPe1Fld1uA94Kv+mMe354t55GNqMDMsHRWQpkPhJw5pqiry0DsE
rcaOmtXhfkOPTnB829q8e1BEi+R57CyHuGZlRSZxEZ9X9qKMCeSoYWxWHsi11k8e
eTd4uJMwKfp7LwUHgYxeZkVyJPHCK91Xoi8Z+aXo9n+wEmPY1hU7/BHVnXtEsSvs
K6idDke0d4H5NV9ddP3WP7mnaBhNJbwoH1Avj7lhpYi4GoQPdFHFk1IlUrebjxIL
mWJhGTaYv1xPs0O1unMqamodw6J4jfgbw9kdPRp6hlV65ck+UpuUI6R6+RznAX1z
WLkaXEF7BQYh9xyfBKb8YzJa43YmG7Habovjv1dhqG+7HQL85OJS602M6oX2D4vJ
m7TuxYBGRXLsy4ySIsmsiN7Jp26dfZMhMwfsOY9+wPNwUfepi8d1VR7TxGqN5CVL
CKUE7U/wvZi4Y35AKy7GQ+dtLR+76DEiKZyh9lR4eWiJJZ5QCLmpK7g0oCu4pbra
qosPsXKpq6XRDavObpTlLeSMynH5GLk4vHgYQaQkBGETcXy+LY8Z9TRrfiASFE28
g37ynhvWfsMqRTpDcwbRe08isVCzTcy+fwtuFJd6O5XiFXvZIcdVnIc2FS7GAgm2
kbl4e/wNXaSg9yeQ+zumLKZm7huwzw1RVNwxaUPp+RzVDF46ya6pgvBpgVEgkLzX
zbOP+LXPytAro5wq/oaKVeruY0LYW5CfZPD/8gs1k5x1TInEG04wygwqWLsp0mz/
YGd04ITDaZsyn0AXLNVFfg8Px3l8uYYmReyzAulMMUsQWwIaK/7zDd2Ugqx8Ap7Z
z+JSFo09EL8XvJPL+ukvZj1w8WYDaoccOvwQgf/7BhEzKgkMrAQG22042ylcjV3V
ROOnNHmZVLbQ9mAnpB/uWQlBlP5fAPMpTy/siuTB9/5urBbn+1+FeAIBCgGJMSQw
M5P7NbFQFpSkFWOyT4QnRpXNQxj5l8Q5j3BnU8JEEAx6jU7MNYWlgapbND5XkBTh
2AiFohm9fkj7SXhClUeitUVoITo3B1rgFxbGvnhwwN5tpTWMMiGg4c4ndf07HJvs
+8M+TdOop4pxDcrKEeCB5+WQzJXd18lIYpnXzxRBO+O5IPFzr59qOwErIQCgnq8+
smLh4sL8xJf0+ilfM2mG+aHr3eqBP9Sa8kGucBp34JbMFhaNFw2sGs68PYSaJb/3
c8yREgMHy/ADTKV6UA+fbHLk3qKdS6u87VTvixSjvfQI+9hpg4GOf+owwpOn7W+b
tPq/ztmPogTSP03F3OmPxaBsVLBKUE8Ulhn3W2hrU2Ps4zUkMnSIXWSjDI596Evb
M99sJoraEzHGcB2AcGC2idW4ckRrF1US8BzXqK9Lv76LDkr0RIzFghyWzHp0p7X9
GkWpERRzI4FXloOMgAGCHW8APTx4E8v9p3V7bI24htSJDFNCnzHsRJug4wRBs2VX
tcy7mrV66aD+ys6PTgLWRX+PVVn8W1to0KZKswvHddxx7LLT1/9cATnSUUVzTeOO
bCHLrfYN01/8SY/YB4XZHXorwGHMuY31wS/dVgRSrrEiFqWjqhIBu0ZO0HOAouM5
yNWXTn5CTqDV3OW1lQrzJAIU9K08jZhUxPtHveToF3nBuTMknPxT/2RuaDRU+ULc
6UvZI7nQfdWmnzJXIfCWRJCHlPq0Bap+FS3zO2Kx+oFYd57ZV56OP7oKLl701LGM
vjlzBOczQCVlr9k0SWnmcqxzkopTw5FND2NioD06PbCVA/Mp6e13m5BhNDdxadYL
Xs0uAZv/KxOhcKjp4F20mE5JUaEeNHUxn7PzGdmtizcAgJFMlRiCrMA32edZW5le
IpsFlX9vsorqHHWmqhCd5IMjYRev9/94CFUg1D1Ll32K23JySKY5ARJtYjW4yoE5
cIll7syeOzDZAD2zIOWowcxIte3ys4nVvoG2j4moQl008IfMEfjp9jUBgm6TRZDt
TAzxmoNGnynhSb0EZQh2abXs7wHqeXBscOFnfvgJPEFOUCmXlySn2TesZHia9XtC
w85eMH2rtKHO1EiVQ6dGJ324Hy/ybfN7wnFQ8nSufL3eRhx2B13ih1TA+LU/LnUW
KJnlZuWAz/CWBRTncPyktxOFRIcNY++yJ525FFrlrEzxMlw3AbBQKrw5Mbe93l2e
lwvpidtWBKvR5elu5w6Vu+RPAnNAmhfwk5JxfZznKwSv8qmIxHx+IFI+jWa0rJ8R
1VC9S8ti70fOz9nGSA3AUZ9Wr+Vz0PwhZFNsWccaoEzXthEDRs1Lzh9ZzsUMX6iZ
44jnFkcQHZRPDrrNAE8wuKCSto4L+SOOtvWwk9OXWQ1I62JEO6dadxk91u8GMaqf
Oks0yKNltG5UkZ0UTKV6H5qrXfsMKMeh9/itVOhi2p55ZCKQcUJqLrQUw2Bo7IkO
5H8JTpEU2djuFXbTEi5Rd26RtVl1IDyl2UZZQcul2y56wfGbQIoRqTs92lZ19Hfx
QDR/HQyQavCLLdUGlnlbMxTuFmS5FJbpCv+CU+kJUPJ3Ty6Rkl+sMuRepuDBDIjv
h1fzdZxpbb+2kUkbbe2Deb+1fWF4+OMSn5TpVoJh8Z+MLMNOGx3Ovz0jwvdY9qpH
/sqqK4/gLkqLztcBNzReLsg4RuZOf/nXluds6Q39pMlQ9Pzy6srMopDeN6UQO4EZ
L5h3O5pnjoFtZOPZaEwta7vVaFRJfFrslGRDmei7Z1UmVkfn5UdbrxKqLJew9IOc
d2wpZQUywyPx6/ofHA8GgE+JG9YayVZYVAPKXzxfWaHBoZ4tTbOJ/1ZDZS+GxeyD
O18O8fPV0UmGZkT4akypfkD58giECYfK09Z0yPcM2PyF8b75E9ASOOgau9FBc+Eu
Y3WpCdMQU5uAvUqGS3cdtBP4eGirvF+moKEM7bv/HAlR0UFtoZVv6JoD53eN9zv1
UdOaCQDdtsnNXZscEF2/ZiV5eelfgQaao+SYfXkJ+bvJI/m+k1b33Q4RSpv91iRY
vwy6TXTj/Bfb9CWMZDz5iAAh9g/4jOhity796TyfZZ/Mbtp2yciM2s1Q0EXj8BTK
8gy/vIX/nP08BHDHR+bz9D2+sB6fnpwU4MQvubcjZ099ntGRifiFbFYrBp6hxZtf
WpA3jeVgHF/JnSt+vm8r1zQeyk76dSwOeWqsZ7/Vj7wrAkhwJEwGeMC0kJejY4zx
erMuWiTFEj6eqaMRxqLRj4eXpw6u662hahn1RP0q8YV/8+xHH+gSiLp/mx0HHlky
dWAYx9e1A6H4wee36kKF+iRPh8CUh5Ce9rWsSN3HllTe6e+dHWO1wAH0jPiexp8L
GCbvSj3CJ7s7SPPn/5MLFRgvV8BSF/yd9JhLzWUOdfN2Dl8F53SjrK9OLms7Zfd7
ypCqS2RbulzZCYra/HQEaSNquWms+oZTT72ZOJDeKPEsWpas7CSJnp3V5X5hgIgl
XLwo1tTZ102FVL2/OLjZ+eko92CDcoJ2Nf+8Pt68NwkVTjM8hMGrP30qzmUJoGO9
FnvAQP3IXeia0I8cVc4GmHrtQMb42r3r/FmtvERzkAoGAE7CXY2M7vtVwpDG/bRY
f2szjx0HSHVIbsjdoh1EuYjaMid6HvpmgkAORpXxUCSN332mLIuL58UgoSyz67bS
qGeaBu9cicfG4u+HODuXBy2bCHK/dpffTrQ55H7EwQxX81gIOCCoiRZdy/ekarT1
TupX3Cp7SdIcOl20uxbquvHEA/6e9neL7flpdybg3ohqkJn9twmMEFnKjQYqVSU8
4GkgnVNbywkos4eTZKbd199cQN0GDhCt9FPwVQephD7yfLCEVYs4OSE81V2P9QJA
Ut0XXurgjPswQCX1oVpgsreN3P5s0CloXmvfE8O1IPvZ7J0UxCjdfScZky/9QE3s
d+6U3zuPdJAtHGtCfeN0Td+S5V4BNi7xd3idj8pXhrGG+SvQX/pjQXT7bCiUb0HQ
MiqlX3KoX6+b7fg6mRLKvbIYJYKMMC4hFSmlFVfe3C7KKvIq/sl51x9+TmI7gC5f
YznSDWUMeGKn6SWQask02t4Y1HA+2310pEWcL1bFuQ/FanzJqF3yfkROzahmlGQ9
+xmoFO+3voPFZ13gYuC8hU4UEAUgPXVvEYqT1S63FX52qDC9N8Y/ijXq2GH7IvmG
RgJ0LbJUOwUAVvEXHahS2AfDcI6MpaV8Imsaxq3h1GOeLFohcDWF0QC34Gw+WmNQ
vk1m5Yh1J7BICLEzaNPQBBIm6XW5d9CNEPi8hjrPvr/xvdwbiAAMLS6gJ3VuKHgy
TVjcrGaLQjrF0+0/PFpnjRPKubqXlHJBwL+ol2i5bjSLXlF6XhEp2hg2tloZOIQ/
1K1KFwSuOMSYBDpuFHwhg4yuVIXjwPj2p7USxOY0aL5F5wc7vxdqqxDD8R8sL4yf
cEK43b7wYOYrbOPLMfT5u/89IeVzPtIoZEN5J8LFhBDH01GHY9bKRZ9LiI/EJ6L7
dvNA3mjJUeDqEGj9xZB1z1BLnxZZML0yzmhiCLc+DeyXN10vt/2FqBsXtRlXxK+U
AKpbklOijmr7lmGHLwMPw4SmNI+w2XCyD1uPBInRuo/zGhFyoJFsTGYzT5yezmRn
RD+8U3EjjhuvOxLlpuq6I9TjC+hXQLRpnJEDVq+EonmRiA/CleAWylatR+bNsfVD
jYbqd8hVVKUIBCfCfzixKJt14Zi8HF2QIZHyDfr7jV2E9qQviK0vVphSm9NlGNpe
iI+5Js/X5nBsWHjqQLF9f2TPqKU9vyFFmli2KYUlVqVJWZelE13h7ceJcytlUGBC
P5WFMQwxVLjPoPJvvhtJ6FtMH4h1/FVpHEs6aKkuRtgZzDf4pfueIGTA+oJtO2iF
fPmEzl644etj5eluIK2B/3mEDjbYUlEZO12UCNVk7x5es/FVmL9DS22ytjO5fsuy
APlfpF/ArRXDjieY3n2b6FilQNH8B8UWxoYQ6ou7kVp71yv3y/IAWd6BFwB1+U1b
hefMHHba7Gzw3TF/K1fdyAPnWl2evwlrQh1rRNIvAgBS/IOumPbpwxBEKxFsQJ9h
vz4KKD0pj79f2mCycC44TJbsxpSbzRT0k15YKAtE0bUJ/c2xn/PrOJa4DfjNzo0k
R+s2OQwV7YeDQ38RBRnghJF6BG9fp07v1MMjIo5nS+Q7AfFEnPcmIRpDFFNbGVm0
spgQYwFQC8KrEfsWsiIw4nryuNtlESQFN/GE+QYR/VOETqJIbjaa7Fbs3yqQ0nkv
dX2LEQe+EnnrXK+9eiwSG47HtjhERKB6s5z8papFUR9JwMJMKPctqsD8twbwqlKq
MSchXn95Qo/OxG3qwtjnML+tGMIbpVccdM3kmftLORk5O8D2lyDgvPu3aZSNU4Ga
Tz8cT5uP6cJrIz/f1I/5qvh4k7VOHyNvAiLNNyHqXJGLQaXEyf/pFZQwEPRy+PaM
xBvp+6ysszGZ673sEmkeQlE1fJBdJTqUNgRSDOQzKzxoCeSuaWCpRyO2Dpbxosbn
taHl3nBFwQB/uLZNdIt4ZftHEGgZu7wV7kakKmO8pwMb+05x+zPrtVHPrydSK+Lt
3kF+dztdxPC4iJCVYHbNbtZXh7FmOsNzJX0Xn67GRWKnoFMEVmZFMxdoCUFmo/2f
Ct0CJfFydyTORdtZKPKfep6kvwvaMVVbILwMz12ejq1LlcLzT4WEp7ZVjcCi0oVx
viVR4CQjP7JoaRI2/8E/iPB0Emlx4/zzR4zOyIpAZQTiOMRzmHZv+H6AgiyZyCw5
ijYFtZdMwBFX9pBOd7P5HQMAvFHi363vC4wOCl7z6dxWwl4uv3gKPLHhfqP+gLx5
Uo7AhcmMgaxW5S7seHRaMYOou3A3gQaqILcwajrJJyRw2Ln4aLAE8g4J/xr+op9o
yB+C2V6zyKZDODu7qV4uHQi6plIclIqpjFf8lHjP6G5ridTrA6gkxnKCmRZOlda0
QfFBPGXyuNjyah2tUFyIZoXZMHHuWQRvEibH3bSSZuI4QMRslBP5HOWYAIWnfGcR
M7RxR+wlnbYuZAU0XYBAMS4ihiMUY2bRF7LiD7aDNNl9Rcjii2MDuup95mm2tKnz
Pjyq/NSaSvR9UdV5EUuU8LTAQSP1BRmNMo9yFSxoSv2jSVx+rMlGJ6pdhNVgpwQF
DU/suNN4EQfR6pbkvImSNJ6q47+/9hfPFLlJFdlhFw6dGYyDokEBnEiUx/F0PMP3
dqpZyO/z/VbB6zrMK1kr3FGN8FOrU44oZ4Y+M5XZ9qr+9xkL3XDRh+owX7EDC9kf
71Memp7DNHrtuS1ifhqaGziS3Q4OYnLwDYklThUO+gec3MKaW7dU9EAF5M4VjYW7
lgqTrOfw0TS308hhSYFq5dRarCDG8rghbuWeKp0k6uSxZd7jOGoP1KoH+zvRFLJc
jTnXz7hdmDmgk9HRoxqtEtSd0kF9mmrMhaKwaq+REd4SA0XMgrFRRmDwyH3EAdZY
got5931DLI+//6xes4wb94hyydZVngp6RyOKFejRXjtk7cFsVKT23vce8UUOziyN
gjyFAtn4dsO2hOyZM3BSpP4VbObOJg7HEO9zunXMwncIqHKX+cM5+QTJHtsstbQZ
yIm1/QkUqmtqIFpqgPghdoamHheN1m31hKBhpRw1e8XD3lLBuRRic5Xq8p8EWU/J
zPL7o7dsfdZ9WbasRSUej281huo25uSVm1L/35XmfYChYUaDoobihpD48u0fqWw0
bhHVjb9gh8LGgQQlGQ3Bj+bNe3ZKVFtSdhjxAYzYxT7wXf/RUoe1YdAyEov5bqz6
lP7MKk204SL8SSPv2hFuyT5jhMZ6m5LER/Yp0rCaYrklyNMtefraeu3mXRqx0QzJ
P4thiajsBwlKjJFNOJA7cekjf/UJwsow0TMkU99MMizzs8fodakdDUPjWBrDbReR
pAZdFYbJ1Rndb1ZA3fBYX1cZUapKLKwXOKld4yQaWd17TJMDHjcPIuZPkb9EbtLA
AVOYhtLk4vjjeqXj0jrxGSDoMIqVg4MDgUDhnRTRKDozpc5RApVSvQ2d9KJzSiOw
HihRvTITYJq0lIf1o8pbvG7a1QuLBcVxq6I5IXZr2tK+2IuJZ9xhnavPnJUWss3f
Sh9tlEuLB62WiSWHeVd4AvGx7bh8BYj3RP9489DRjx+b61fSRH5nXfmFG3AGnuff
Nubn14J91/45p45Zar5WDqEUNCyix874tmWUteAa9qvaW349tKURNEZiofd4XMLq
Mi5i1iL8TkOW0kitLZOqZpGcdJwcmaWu5Je3Eg1e1sxDsK7GS28I0F7DpF10Altg
sLRSuizStDvdyZbnY2GjQsTlnFyjn+ir42BmtIW7pe+vkm/lqX1FXbWbRxWovYd8
VUvPRk0UpHshtuIPtRSA3KOeHYQfGQ1gKGwrj4UnM95TOfLO8ftG86NGnUlRfj4V
z5cE+tCM6VUuFnf5B32HLozdpENbX00SevV7+t7UtCEZO/kuR9+pnZakThL/cYy6
dKlM1EE7JqCbjQRe1JJhtCOflC5orTC6k9pUD7nVOwx/q+37MdhZsQPMRIrvaZn9
EfC8DjFNEi7QbvCRLg9V5OCBrg/kKQE0s9fyJfSm8lL9CG8vIjq1RGWPv8VER1RK
CWytCZ3zje9YkctlbGea5n0ExzwiK1rkrIL+cm6zMD5J5HBe3VPuQPcbWmOm8gRb
5ulkTR8r2aKyK2a4DzJcrcAtsXI1a5Jg5CgnwMxiN2h6V73lb4FAA1z26j8ceW0H
YNVpnTo6/StUJb71VlHD8kO0Vp149zgirNBbhNZ3Tuj46wvUEY9GndTclGG+nknx
nc2MeB793vHsvIdYxJovgCu4+vmsYhFLiClePkXkLFX9wyP0q1P0G6xuZGG0ugXs
a6wbz8AnMd28gdO+BYoluU7dRg9UwX0a/uM1/CJkbjn8BXVnd/pYVNYTo7cd1ptq
dGmCttl3VwxZUHLuJ+w/64LRStIZnVJ12oxVO7Pz0nBTSg+lzAqb415AzgRpdCKT
TmPCqtF6QzyXobYw3ieDcPePiV0WjviSFw7++e1G3DAGYzDha1WABwa2CwhDFQou
KKJYV6i3PKFWK8ZhzyHSi+qmfFn+n2PfkE5BL+EBAWLWZVX37C9pS/UIEbeSalXv
715TioST1IZlklwmcNkesPr5HEhkmj3rN0tAktyvqHrsztpO7GYwr1PbRQ18x/DN
CX/3Dk39l3aaaeOkHX3TTgcxuxaW4vpiGk06xfs5IytSHN1OKuvimPTKQuTwBMDw
HkEVLpMnAKCtErAP4ivnWZZRhdTZ7wYv3SsEjuqPbquA7xBm1+luIodIigZgTpth
Kmrkp11GRIgWcCAX/ktgqyiB/hrelDMVXP+JNP2ljSoVEyMVnVpyZCYtGo3Ztfyc
iont7g+5elOPA0ePyVSy2Hxp8KImEmbtmwWVHk0nmz3j6wA/err0Mv9sIU70yA/x
DQZmzuS10rR1KMwjMa4zVZpfstVvJE3kf4WXL9vAcHMfSRyH2OHOaRccvGnq3sbW
8N7DKNcSFdo+90icPK6Xd1DDLNom5/F3F/3iVtxUf+NVoQ1crKlm03H+Ow9qqoIN
/GRtxJrtCzb4soJ7A13tk8Okk9gUtNGu/ZD2mn2IQ1WIT+tGkSMuArhZawNNFbYe
ZKAecsv1iPISsjwG2zdmM4ntBMdl5eUKx/Ph4349Vbp0vDwusa84L2w3XovaHfmd
pH1osmprhEB1rbu7UNVKQ2YeXaslYjhBld/oGfiHmaFeRBUayEtQOw3VfIRutSpq
7rI1sBYEScHUD6LKAltGHFPWo5a/++ZZidHW8IurKW21dxPdcrdKanxTvt8tOLDm
hPmmfrakH3djMg5csaL7kmb4h6j7dVXaaQ/bG9FBkUKiRHfbBJSFuvT02Oh6Y8RV
XhW2hXYZh4iIMpim4CLXb17nRPbEVUzfK35vmOz3ngO2aVvHtJKYcWAV03cWYOv5
NT9bhHB871c27u5Ll7yktKTvQP1hN0YFQ9YU0BjYZU5cWTCgChYY7UCLhMK9VwIs
XXzIHJHWo69vx4mIgozMPcBHoisowPrSaay2k7DgfOzq/RjVRoqBl8PBhSOCJB2y
RihNDPqRFMfdpVm/zf71Gbl7Wvp1T4Rti+aVzEnKrQHL6EIstTjuRVjzE11sC/6J
s2l3NrmPzKMYbw26uQrS7uxAnBX8xytwIh59LdnWdAJpl104RMFt7fg4XyiBsPZU
U2ZcDiMGwmgfcKhmD2Klq/d2BTvoe/lTY4QMhoYW0AozlxT5OnoH8icJJPxOwxEd
fM2h+SHc7EzXdfpycb5Zoq1WlwZ0THLt6/X2Rk427mYY79V7myXT/MAVxMPAZCzP
t1kE/Zqy2ifDxpbpnwekai9fEjycuzf9+PEVu68NKRlMlAXXOHeGFs8b/cE4vQTE
5X7PiZi1TwXFPohMwANfc4YJO3eztBQv7rgiJ/ie05x0aF23KPtrXum/PYjmIAKy
FqHChu+NOslpmUCZFWKhOImjmzpZiTuLVISrKrVCfZb6wuXIjuzzHjG3yhCjurTh
fCGpJmKgYdgaQ+SeXxoV4yAqM20Yu+qXb0282dd77p5WP15NfZ4v6TFeiZV6xAF5
wbG6NRCD4vQQPTQF+J5oyK8Jolwcgs4ATqB3kRFYIymoG544g1U/GZfx2j7Lch6p
eFA/2ElNLiHlkcpolh0EYUeJVfRrEt6scx6lTCIizXS7mAJlGWHYtMQZn+7uFVbY
24t3URBmzwLW4fsEal2IDMfpsgZVaJHcSN1OXZoiQBlX70CnPlUQJTMQXlEugOiF
DKJHsQhWBfdC5l8W+c63wD0/AB4t6oIVc5LdsiLBc/K2R7pxbd8/kGlQeJwlY6QE
kH9OlfWxHlVczpvkl3c+yIWYCfQS1EP3AwsvVZmxLINph1sQYCU9RDprM8tu6uJM
1/bipGIylZ29eCxVtXPxt/5oBFzDMdj8wxz3ZpUBOr61/g1CLDbxMosv8N/vjP4P
pScFFWe8D4PmL4YT8lZThg9BrKubYFemAbm3ma8msCHAJs/yA7vtnxBssLdm2B4+
0VCrXqK2U0CVhAwGrscI4EBXgi+0p5n87XG7Xr5SOWYnTHFOkS7Nzp4G/QlCygA/
Xn9FGZKAUIJMR2RfzPe2nsOZsnI2AHA+gtvlDfu8f/ODkRNa1mL2o+3yGkoWVsfj
h0SFQXCrRd7j7fHB8WtLMvrtaovMhXn4Goyejh4drR+pewkgB3oKBvCldAtHIz93
sLKcyMMBmwur/98Ho94Y3l6MtWrTDId2f8FAt4mmico3UcozVNQbjIVDMIYCAjxA
/UFq8NriZvTDryRj5FESGpER18iy1Nh/OvN0/yTkxwNRdTQ7tluCpju0mi9ct+Cl
6bTsaRfEGTjbFbAjTmR2LEwstWOKr1lQPCaN52wRW+n5HCKyLdeKmbSQgbLXoIzl
wm9Eee0VsU/r3V4R4TwM/L6aadE07vwOzP7qXRIkEmtDPuZ1UBTnQzQhBUHBlWBF
QFss0o0VciwhBrB/QwsDCowoSo2Bq10cBK44fnOoSI5KQ6DkwzYyZ5WkzcRHTDI6
BYjooHhr4naHH/K6p0HI1djz5ILhK+kcMbZMyo9AhaGTZpR7tOv+Iz8wuCd+v76f
3h1VQ1AZwI0v1/GbjIyU1guDYmvia0K8jszt3AitnksjiK4R0E2RiFw1JUmblMML
OKzb1VaxLgVtJgmHFCjCypslise9nI0u2JJVmjfnaYE3JpE+oKrCsRjz/XEfs8Sk
FJnt3E/NoOG1oatJpad8spQjKxpQOSzal2++D8hxs2O/ZhsZh9pfuoS0ZK7v4Msj
C7uYZHwSSsYqKbLSG+EjX0fBFQC7xa3vvIezmmbugzeAUHEYUts92MVm8ytSQDhD
pd9RGPavyIYAZJypJ0rwvppmc0JILLJhtMu98UK+ejcYDVjF7WySsGD/EZCxLQOt
8bpv1Q2oLE9FsSgM2BTVcszk76ojdUsiYG2pnLb9jvT6aSNAIrqWz4zvQYoufFsk
x6p5BaTJmNsN7XIqBXcYKL9ahpjJcUNnimZQk1Gfz3PxPqaz5QLWUHMQ8eAHoKf1
Gl4HyamG6z08i6kIX+jcnS6yB6DitppSNfO02elXovGgFXsyealJlHUWcjuCU2Kg
PkWgOVNUzKshf/xVZBmnvlSKj1wKggGiGCKSFjftIE3RJdExxO7BMEI1cRwUG0m4
FuqHMzKxtOjgRCoXP6h/pHGv1DVRLiZ5Iyw2kA4/HQwXtmCxW9ATka8XmKCmZb4L
LHTtQeDgJvbwAyZEhBoiVwZj1OeRT+11IoyCKhlJ+KBys+b7dVI7fYhNdD53NDgZ
98IEKi4poeOE1ishf4YiEoj/K26+z3FD6wHAUpb+wsh5Q+10lzyzbrMGMGoeQ8Dc
0qn8G5eH51ICVy5ZSY7UUph7Yw04HxvLhpX63EUPX/0+c+2ghgqveUkaeWXU9Aps
p0dU2e1GczXsN4AaYtZTQIYAMtWGQzzpnym8pi/l8wtuwW0wkJx7hf54UqI6wTGj
WIyh4fPxek3iQpI5AV1ledEhOfbBiOfDXpAm6SqldxXVptlinW7TB6pIcGsqhzb8
Cg+kHp6Loq5ncKkPKCRdT8Pj6OFOcY1sqOtQD/uzcKL1/ZSl1FZav1JbiS9P8Kie
5hW3pXpUDuMZg/NNlWT7VE/7F//DJtHLyC+GsnnIJbTn0NRBtK4aRG0r+DRceqpD
a6Bk6TM7HwiPDd0AOC1I3djbDUN5JS313WfXDNxj4t2focLwvHEYvju7RoWcrdaG
LucTxf0j/2/3gBmvO2KraV8wAA5ULm/kOt5d/SAaKC+/cNUjJN8LKmmSrqJJqRR+
G4/3MRBtzsGCwiIxDCDTuKnzJR4/JbdB4Y0o0HHquCGXn0JvUIOpNreb+0LfLANB
oFyNx1IVjN3rHdreSiFaBifl1xkEKWy2zHaUb2jsGUOgZSy2Kym+pakYUo1BqB/M
zcRaiQtB29Rj8rJ/9S6FHlFsgDIi6ea55Ny3OtJuIw82s5nCthDAVYUkL3qqQ5IP
IXvF2ao/sRJqrV0W52rpbMrQpuEUAqiIFbhApbxy+r77eMh7/whiQ2m3IHOkgMy2
N3FZdzec1X1ecW9h9V7yAjkAK22cCjIIoDzQRYSKuXw8qtzxbgtjPut8h8Kaz2WV
/XVcnHn1Zxkq+pvbw+ce6ed1t97IQdfOCy64c2cYPT/SPJ+W7cD4tqyh6RWQnLfC
tsIfM9KKqJ1t/M4JLpSsu4SE2Ay2eflQyIW6ZX75hesjEtXRB5UiBQxeJjJ/O/EN
9aoV9f3MDnL6KYHhc250Qx/4LFgjWTyltFtYfTz4IKWu6zBD3b5V3VjWsJRj3tlJ
R/+qmUBQwFUQWJxwtO/D/nr+puc3wE4VtoibIoIzU38fgSYmW65Wrh+W7shPE1rc
cu+XnNEp6GJdfCkAlil1+aLxFptotqwemXogomucrEtKCqZmSR2T7GClcc23Ggka
nFiFTFAIGSrxQ1UxU8nibVqc2ZBFmoPK53VQeRJ5Xo4ZomUHzBE6hRXdbFzLPcCL
B3AAFdtwnbQCBshi+arDBARjzLPr9pe0hOZ/YGfdTOi3mjMQ/x4WPjZxHLyZfsG0
Qvlu5CI/qRBBi3VzuS7fPxhTzIJ4HHhMZIXwkRUtZVwH8GEVTxAwuVDrq8vsQPzC
VgjS8uCjyXebDQKHV4JrRDcmanrAYkyhr7fPRYnPK7EU5fuMW5+p7ssVpVp7CsoH
T8+lYcXkIGlyfQE/REA9iiEqGfuCtmmP1KtG+J27tSANIGUkacqoV5hLMNkLcTD+
nbewoCmox5bvJp+aaj9rCx+tVRN0wG+o8fefL9FgZm88ABug7Ixi8N72E5p+Q+VI
qKzfcFMal3Zlh06EgLDUVmQZxStyUOkaCDpyUvCdOuijmmeRRnd8wXntmWMXq3xN
Yamyl4i0XS9Lwc5zUvssufMn8vXRnO7LCdnVXFgovK4XD5AOiD9CtCjrcd52Os8w
uorJEoOqEDbtiHOtlZfh9t+3QLlFUn0Cl5QhjTjQcdW/yPFkMnK9TvJ//jDvJ7Z8
ShQl1pVWaWd54AWIJQVlMlB7nfOBGrYcT9cse8eJKFzdMQT1zqRV8yN5+eGhUefW
uOEBLm9d2wccTssutcCRTvapmPiLhFkZWCAh5I//HiHSNXVEU4pIpiMwercURFAz
il9hT0aprneNu1CsI+G1h/bjRRz4PYcY9ndDZRVaHhA36oZwMQGj8+UG+kT9wCXK
N6ZGDBMy5yixpjcIqfcVFx77IWS84NMqJcp1nQ27gBqwAiI2Td7hegN5f8ecWDuT
0+5DJ/PtbX5+jFzHMC3ICttXKKt3lFvWLNyPVo2n/PZ7QcUKLl5kBDvXWeqDRIaU
Kstww9PeyCrSXbjiPzbfPatiUvmTY4gdFp3sdnS1YY/1eyklfyV90Evfd6E0B/YF
sVAqv0YkNTd2/KdZQXJSEa4lNOsfGmhpNZA/zrATbNcSIXOatbP4dDk/f9c2t8jo
uOSdq2TxFJsNANhD51ReNuLeTW+VBpAf3tMAbHZmh9DKQAIzJuFZMrR4ovlcNy2q
Z3A4SrOlq9BAN0riy13LVJa645NaSSRCry3O2JZlafY3D/gl2M10zna6rthNwvAE
sgwLvs+izo7Gxko2B0NU5K6/o7LMCMN+UttMCuxwKYefbkzTssZuD1agAbi4NLdy
2goKQeEku+KPpdM7YBvU9beRrmsNxcAGAPlIYXncxliogXntBhf8RiT2gDz2zcBH
hh9cNKaG04kgAuJhWiRszzcB5OPvWHC6iOR4HZaTi/DYm8ykT41ApGhvIVgo1lHb
KGuOjCMFNc4f2EUKqIXcc1snLepjb6mpSSvnX1dZPba08IwdP/GVjE6hMLhtR5Co
ztbZj2hakZqlReljm2cC/KnbDim41BRMbtn9xdZp2CYBLy9OSguu6lwiMipHlhqE
hSKHDgOQ8nPM8io0yWebYkWYncbKQgos0AfM2Y8T7hPSBEIFTV4xWXv7ILKRON4S
UB9c6VbdZTaKyI+ZQM2rAJaGx0EkDao7Au9uBr5y4Npu94jhA+uGFtXsOVmGffDK
3EgWGb6sWnoJGBo6NMu3MSj+F5ZttvFF0NrTeQ9v8gpY6baJc2kGvjFimcahsgt3
olTv4B6l6y72uURTBlacu3jb4dmlBpzWQs0Lz+xYd8bIvMFwkxgCc/MNc+bstIP5
dkFtFozOEsF/lQH8/GWG9ZnsDnpL/ncXDDIY33lv8ieh/oAUQbwFyFeyr+X6p6tp
ASJ9aTKidWJGwtoba7s056n3zazOKypWlheaRXc9Luv67J6REU7f9XvhbMXEEo8y
GCBDoY0qUweBs3jS0VFxparjfvczuguwjbK8VH8LQddfJLvH50EmY+aZTbUB3vyn
O+PtZ8u9T2WVi58UW6zkVYczPfnhkXNfAWP0lp9YEVvb4SHVz0+EwBSC8X694cDA
RQdQRaaA3qFB4Msoy7ikazcWWcE23Sn/1xvbt1MdRIfOt3A6LgEpQTpUMFQmV6L1
m7oqjDkrClgrrqqREZsjNXA5PQO7SaIgkoQMH38lEWuiOxytg6AI9k3JIj9CxpJr
Mx9AUk5XVxH/rR1oTiJb1YTne4mPDS3U19Ia/tP8HOkvuEJv1uBOh8HNmqnBiY3J
DjuqEhgRcxNXdIhPxwvhsYTsPFwQ6mTz4qPIg6YRtXW8ydMm4xKd/Uw0RCdQYSBc
QcomEMIabYoi4M6hYStK+IXE0EQsobCS2kpYeOSKl8JGbl4gdcUdgyqRecehiDDn
PXQ4zOcilizSD69tGoARjykFNy5v4trZLOZb3x/hxDC84jQF+oQOKnD8+bt7p/L7
4H9NUhlru2KzRSJfXRA/pituLIYs91NcgIGcaeNzjKSZHoRlfQyRm9WR9DV5R5e1
fMOQRBGiGqfdItIepfzXWkR80ZmyGi+6SCcEriiS8fObEkLwVOMzLHPRtgt69r2J
O98KvLRgWpK7bKF879z/JDLlQ9+E0G/49UNuF8XE2iBt4oR1c5TabS6hcIxvvWeX
ZzHJZPwmY5VZxSSf+NLeTSSnGBRN1I4FZU05xJ4VCWstX6dvfdIolk43a0E39z8s
RP/YsrSuy4jJ2mjJrRbDJ5d5t9ZFs8jXfFN7f46/K9HkIGDKJ0TZB2Nj+h4YJQTA
cfDFcH6bno65lkkNGbLfss1//y14Nali92nNw8QpIcOEmftBuf75CqDJq6me91N0
JxvbKzmlAdNv8HhUIHkr4v3bNjbFniuiUTI4/1ekF66oe/aFPesHffumxOJiTipT
oBE+hHiPCONOH+GRbzcGk21mCQMMx8YGdWWnERa0mCEoyTeh+QhywipwLJ+DgStt
4WTSy/NWi+ICMJsE/s907wDMy4trvmaUtTU334ddnF82z4QwCurh2i96KfODY04M
f3AOveGa9oCEnlRpP7UycMOJQ38xnxAAX6+J6Qtb9KfPJHnh/gkRLu/6o2nqTb+e
OM9+IcKOGCCrWS69/pSaQg4OGveajAqsBo+2IOyYo2BQTC6XZ3j7aNR9DBLtWbcO
mzxgMSoI+x4NlUgfXX8sLpYVmB58mwWl8sj1ZSHfRyjoBWylBE1XH0O+3vbwyZmk
z5lU3RotxgljQcJ3nIK1wnLNBIfPq5IoATkptopSESSJz3kzAz1GUZpt4ukEtjXf
xnhH1dpwgbQ6X6IvAYnk7VqCjBtlLf9qUaEs0PsAXCb0KsON51RqZIDNXFZJQcCp
6mX5/KsjRdeULTaLDN7Itvk/Kl6BX+ybUZZKgI8C8hHToSEd9D1qfEvH1LjHQvXK
O7wnMy2JYeFj7FveXM1KIlu3uzGWJnumR5/7/U1IcyCz0mBXsYA3xcvwYJLd2+4R
e9XeB4yPDWGGhxG8QRhM3Ts2FhrhKuhvWLPL1kQGHoc58eQRODQWgiepI++quJIL
JirxJTria/5BGtZQ92cOjG0vCBtZwNKEZ1SP5u4aPeqzfCyWml2ip8PFetggppmG
d6yL8uJ3/4Zs0TsilM0/vDuBGgQr/Q6avBilPOnNaugAvDdBaQEc4uRzGbCQMTp9
hAJNzVp/4UB4j+nF3WCHGRmSi0loxbNCh5twp1UJRYjFRpKAAnUP0L9A8RjbbOpq
g/EOAFjwT5rYoZWfEs4DcVjT6mQZ5Oklr5p0dRMjnGGoVuG/g8vZNBcin1ts3Ko1
2/sm1kJfaXU2CCO73LZCwfzElv0y6/LkOTSjTkBQuGAShwkdrq5ulRHxVCmIBhPN
oFpx53x+IXMtTngFR9UmIS596wJh99VjGzikCHGw34TKv14b9JhdFBjJZaFP4Sbg
8dUfe9n/sopY7df+UMFn7AksgfKcxuFNhJ6mzz6i9PqPdLz5YXock21XSZf5Qdnx
gLReA4epa/3pqo98MdfGcC3OU6mSVCiyUfu+3NZktVs8baZJkrXm3KT8JfzPedwU
hl1u4LGNsflF3ki9AIh4H9tiE90xz1WZJJXVn/62l95QY2NgviY6BiDOf6Ied50a
l7FHU2aA4tTYUt90vnmMwlKpYKMhVqskdGMqrP6kDq7k/8uB1Vg9cii4XT7uBWAZ
frc6rx8nYRLUI7GFjMIhVh6ftiJS3CcLL0e9JM5qbcZ49fFqZhSZ+O320yh1KQwM
sfdWYF5xSqrroGc4NFvWQ3MCio0vSl9F1+8Y4RVIII550cVLAufaXjRmsCmXRAGF
Hd6n/1iF/MrnVqQ+16+rzCXgeRzr0olqIEQcr1cr9eHDCCo50pUuA7NgTL6YZAWu
a7KBO00nhFn4XuIgkzAfag3Q8F9FYbS1NYCEMFMk83k6IpiE+gwutcFnt0CUZOx9
nEXfAWifbGLEKbFjThVLTa3Kx9fU3U3+sNLGhr1hukSzns/PQO0O9RPqdzkMjBf1
HwolbRJ/wA4yW1LdJhVj5vc9ggPP7WZuXpTMaCnHU7f65C5hZGRYSyVXd5Az2DIJ
iAR4+oaaN/GLOfDIGmvIop6kF/g6f6/k2exIeuh+6z5pytEhkElo6sre/x9wr9TS
RPapvWzs8OaaIhLSUjS2p7RAQZLxkaKO1g2o3LyTz31BLKiHZSCl4DNeAZyjzpEV
NZTDT8Hvqn2xYtCCDtVtab/yvxVaSa2IOJLk2VNzlYPjWjQC4nD8MlBZGyq3kwc/
uJFglkYY7zZVvAUPhqDLBaT9yVOPdlL+87tGjxnw9Cn6nPl1Eh5k9EVWo0Fjlni9
zwXk7mnOwqFxYL4TKcjyWJvHmS8GqKpJeDsNWif1CLtjOOGsm9KisPdyx+I1ucen
pWugO8uDiRxiywL7d6gw5X6apWmlPEMQmCT0FQo/1r/wimkq+fL7EsZvPj9Du0dN
5Iej8lnGpj+TDtF16fJNXrkVP6V2IytmyQd6df6ATodEBvOLM4nzTL84crL+fMRU
x/GPiGeiAWBhYVhPQREGf9f7u8t3jSHnDlcIj9UuSCr4Wm9Q6VONfiizdVpdgB3F
ToHxWALwCDf6PIPKjAmJx2yR+xoz3pyqOuvo5rKwfE4VWjekaEQ+eWtrgR8oL029
RSHwOAaEC8XgGFTEuHB/Zov3hEwe4/uf6a/r6hsDY3ofhqSm/CbuN1NYZoYIVhv8
44o6OHCIICDbQo0U4ozNwdjZUa2fK3wCrCeCn3fXj7a83qC9+LrijH0m0JuBFJ27
hz+crnRxupSXBEJariaCxsjjQDyxkzpX4mnD1opxDsedApda8myPJ7SIJDUl4N0P
iOehjwqx80XX6Xj0jUQNk8sNvK2SeZBzxSSdoIxfyrYEOGof2h98mdlD42iuCfBB
QhH9svCTfokSpG8lfh6h1W5fdtIZoecwJa4RG8KCVewP1WFLrLFwFiS2wA+z6/ys
fry+cOknk/vDIjics8qqtyUkooquLIQai0nquTpJqWR9ly1ek2T31NHDOo94c7L1
hYZXYlWg1DD0YEFl1zD2la/VdJtXH58M07I15C4AnNh0+Xxn3KSnNMlT08A8VZCV
e94hfpl1jkeeoqWFlJXktCp7gBMizGU8Jg8kEQxdH6rNeflS0H3wYd3l12LKwF+p
T//lF7BPXMuTcvLSrRaLMZahu44QM0GyHpqyQsaLMDCPL2xoIsWcdroCbsCAgk8A
zo1uilf6AHV4WusR1aUm2kQfS4We+Xr/ebP04pKLC6zq9F1aQm9F4KbS+zv/s/tE
QdCnmNxyKF44m9W9IczvbVFWAx8ebh9U2jKCrML4Y/qBWOAdQqyhDdFO6VVO4HQH
7U95WxR1boEHByFiUFELhqqRj1FZ0LgmXZC2MO9xzh9U11scz63uzzcel6u8WAJs
4u7IBykJHyxWGdShSBAiTHMMCFQnHRdMNQTXWhwq1LuW/oviY9qbHSZ+h9rQsdQz
+k2s8ro86vFW8td31dYfOz40SSCY5aGZ5WkPt3YKmwh4Xp9aiKKy8XNQ6Fe/EA1L
8o5t1sHxTIaPgd4C+/hNeYD8drHUkCL8DZBDbaFWO8meIeiioX4zwbvxH3D3EMcz
gD7+EmosniHfmt8P6WH8EYYv9iKG+R5jMefX7fvNHFjMmRPXtrai13HJ0xuhJCEz
u3Ztacl5rrd5kwmMOcZuXidVEuOEsZqURfobwmSeAoGIL+GWy1qJOnw5EYCjNoBU
sKHBEcIepJRZvd4lqn/PNEDnsrNwT/JldOWbI68L2PhbiT5rSfKmLiaoFUu7OWT+
c/KFeuMwVeK3VhkMKb1CO5cGMyBoJBqD7CqfK49/RUDOfyaCpXCJZSX/gXTo+gqT
0wmIx1QCQs6t6am8IZahOnUEGGTYswKIB9N2TioitCeRo2jnGo9cheRIZVWxUVyr
dP/Axat7TkSbKIG1fDqv38KhI0zgnwSv3shixTS7MHSJv1cmbc9xtdy3hFcDn/+z
G0uDaLXecPeudGEjtTdN/wAA3R1xTUY+HAUYM7xmaZHIyT41aAFMXrYC5vd+IDkE
VQU5ad28UcbOWwFuIlrUycxjlsnEQVIWMKyS14O/5ZIKnPv8QRI2+PkVVVXDG9fY
rB/UEX3SiElQoVLc4UOpQ5QhsopIjP6Sl3E3r9UbmCnjvTFqRH/lWkawNA0qAAUX
3gf50/A3hWAVjmgtjLFUSg+gMszvJTROPyR0H0TuH8uBVCciS0iXuHZSIaBP/c85
AAqkSWhyN8TWJOomzZhI9sKbrP5CBlG6f/UcZ/r8iYA0KLzCwt/g/elVFWL4KxAq
vFS3qBBwdxebDP57VW2keQSZunHz3dGDO1GPbW8RRhda/LKDUDQwaYwZiFyf5Z5k
J3dCSNAgyZvS8w7odhh4lK1mfloZnfWQdSCUThnoo3JTG0fl9kgNX7sEPXCVry9F
JO5Zd+HN5FP6mRqueQjDAHWSRO/hbNZ8uyiYIoMqFbTR2BNMqwe4VUelmD67ta+2
sGD9E+tteTCf4tPsfMoJ6hGN2CdEknNfB57fnzM9sufNUkwN/xR5Jp1YbETaV4dc
mP1yPSIRiNKneJTfGAubZz7p8lNRDwrIp8Mwwg4g4rQ3ry1MIK+7Zw6AFNRrnbUq
dMlZy9W0/0wvpra5BtEr2bRKjZaKrfACAgJrBMj4SPn4TkD38GKP++MWnYEtwNuA
Ku+AytmFUArD/zIVNviukaCjhfirUXMVfZ5whXm1e4p/tJjH7ASOgt3/Hya7ZMDq
tLGL5y2BboEKz3rVuh8aSw/Cyh0CoSH8bfPyHUjWQ7U0f2FdSuQD++0TSzCHIb8F
jYMfDR4+U3Yy9cNt5UcJLWNyWdgqaiXB3O+S8XsLy6LisuU1MnXG4KMkEqTLvrBu
s/H9FwiUvJ9PyyBWgMaIp1n9r58e5UGvvOD1gb8Rs8O69ejq2lO2SJqF+RUrmC2l
l3ut+TmHLkUcgRcYk8WL8EMcTeEdM6LvTEJJy2pVzVpf4WdaAx8dUnp5wEe5LB9n
eteWNbchSNgQTUbzFO8C6Lr3/yQPOkts8bEhkxlhfu6ByQVv6ob5+6mxJ84Mg+Hf
Jn1u+GknsT2txd2eZFZM7uUeDKgrQFQC1NvpJjsuCU+z6oYhD/Iyt7v6HV3+hXmL
AkDtpK0n2jYbRWlXxmehkMCKFryGodmL626/IJjhNeCnzERNiwWyXnNg29Xa8noq
HhCyKe/bfzzAZ8xdUfZ57hnoO7Hb/FgatnqLgJbgGtaIfWp9958cod3UTrpxcQOj
ULPlEPIIxWM9/cmgkEtQRM0t+WFdb+N1hqwsJ6r904pPy0kuB8s7Sr2s2ZM5I24l
knioGEZ4i/AHKhLxhwtnY4t4xocw3+lxGltYCIuBariMSNahfiTkPPnemhkz9sfi
DgUxSi93oTXTP/75zm7dCQcI9NffsY5stIU7EdHPTtSuPFi75DiO6a13eLousRDN
04CDdtf6oI6SvfusYEMVal38+zCgJWzk9AF7KJdtZlOM0h0T7+DllZ/y6vlZjSyL
vTgubMfulkB3SV1ZqkU/kYkpHp3P1LKhA6SMDJSUQa0aHueVFp0LAWJom8BAStkM
3Kd5HXENDU8rJu7AvSgu3p2az17EP45d7RgVMOxGLKFso20+OaQ3G2sPcoXoSXzt
WTP1W5qLYU9sWKQVSOrUKYQzEOHEnc027gRdQLOobczmwybTslVmLgphJuC9sFco
VVzbedERzNDpjtoKL9TME51UN9PT7oN9JsPawr4Sb8uBmi9C1KYyqVaHB6Gj9HkY
vz8m9EGw6xp9Vs7ydMJppSGHIZCFCOwjMVlgmhYT67ab6CZJXMkaEDX9QMKZ30kx
YwTA+CYiHu5Guz9qGiJkZbRHRsnsr0Krd4eiPKYVKxClY5QvIpkP6V6HfRvaBSoM
xj9/K2cS8luNGbvrO5Os6wLKIfBED3WSVLsSLlhb1cCZm610uRuOs16P84TfHwmJ
Dk1kPgFekFyPBYbJG8JVTAStnVuF8w+nZ5oZj4FA67W1JjjjCl4vgDX+49wKdVJ6
dOzVLHj8rPoihKA1yUgUzzy1Plclr5Cotxzzx9eO94CYeRD+l68wvXzXAVQIzrhe
aI/iOn9WGFkvBdTQU9CcheGjXd447v6hgBnXymShmxfcECbeoVGD2xR6d4VrUO7E
SSoDyIi6pznADwRBBR2eu4miQMoZFaVItfAV/6BM2UgtBbjM/PPT1joDKukNmygl
jgVL9kjDFpXtvxt3/Qk8OyircFAhI5tB5R/UaHFFsyldSiXdZX5InkdiL2vuwrTc
vEVOrKXvn5DDA5aJMy52ekz/FwTqkgEni4IN88XPfUOKZOnk7s1XAxEaDd0uQTdi
NlGZ6Q9j4pRmxjtV2EIhetAJuJs7VnE6OHflUNI6IqKJwxImeHI4ExIq1q0N9Av/
5upu6WgER9DMUCchL1kP9FuQoqvfhx5MaAbMrhZGUnD1GUJ088BpEZCLl+vtJoOo
WLTaL0CWU14W9RHT12zCYSenjoXs8oYyJxH8d6uKmDE92PYHve2/lmJAys8U1aI5
ZK8f5o9qCYFOWH0PtMNU9AyOYEEG4P1+PZYmneF6DFmEpImAU8pEb189F5M9jV9F
RDrOh5cQXpam2HmSDuWu3hQ+rXkayJQNTLrCqedYdCGOvsMvpP0Xy8lquhgOiVhH
OLrLVc/0FFJDmAOAtZICOXV08Dzs0h3G8C4fwXqpfDwkSK+JJ+BSfO/Gvypfs9lL
6sr0BKKbB1sB8F5gRUETH/RyXVQMoJblMdSyO821nRW6pFTOe1EVEyioNe88rTbc
OZLNvYMD90cZwpgBMnE2uKhzpj6o0dxsyVA21UeZF6quZQL9kuySYguWZ+aYzlMZ
M2lmRfqfNnUcuJzpl8JZmmmzJGXN23gHqq/MwK9Xaun4Hojeh8Szs3Mzp/5kh+BD
8miK9iq69VXUx2nGy001MHP19IYCzJFmoxdBpc5meEbEHOXIaDTs5SqGF1MavK4N
mTTe/mi3ADwdV6fym1z6Q0pZw7aGiZBdNae/msKIWEPR6VVQaZE3EfEv+eKPKcgv
o1e8EBbSM7wlfHxNPYHkaTo4kQzme5naqV8Xj3gp9dm6E7hjcGVYuQr+dj8oE6Hk
FmxpuWiC8VImpJurWHTISNLALFmMNdidFpm+Lr5COUQKa80qZyCaMrhYGGHnL4/J
mgNdmr1nrn5QV+ESPRLCjD1o2BTvzB+AoH7PUkSS7ITyelVFKUw/3aX2FppixbIB
DqfnUnF/uBMA9t1e1D9hpQDJYejQG5p61TRqu6dQsVMj4Xt0T8C9njbY6iA8pPLf
6gl3IAf83S33dpuQ++mnZm+hm8jlA6X70NnWYyEYDeyXsL91zMTSmFEZ7ZD7HxnN
kuP7RzhB38e6fWCClgXd1MslgHd3DXzz3K5GIXpNsOGeRMOh0BjUE9mv+IKLC4I4
2QY2Czy3MyI8d9ZCBovBpOQNLR/T1z+YoBf5ycMhPPNBOkBg6IL0j97yejLC0W6G
OMxEUPr9CQ7yYdTa7ovUfV9KPTVhECAO/cRjv7hU7BiBcr/ITSFDUBDmcjsqqp/Y
2zPTjZGr6P6j5D47P+UpmdAnTSd3ci3HatOdgyFB72DKiyhx4XZ3JWO1qvpUwOXa
GYoO0x3TD1KAsrANz5UPvtwWwVSFALrCii+K1gv+gcboCoi8HAVSYLoh+ySvoQqE
6itH+E3i241xe0UFDo1xbILmy2LPXzIMbyHNEjgCOPBWTaV4VEs/xCTwxdjVUy3N
6D7XeuEYZPqaqz3X7xsHZs/CgkrEqjRdCvLv2LnnAxBFDB9QnRJrVpwt+ZXAn2oM
GjONfm13c/xc1yLdyZ6Irg68+xQ17JE0l78n+gQNg5jb30JRZVGlhUrr/VZMFojU
haZHbPxiTSEDsXM8mitZhcumAqPubPMlKZ2iJpEzmQSsAMQSPCa5LB9mmT1vPJXp
8eeQ4AHcOsFRHu2mwbwcMMFLIVK/LFwKJvUMqF5xzo9uE5zRJ9woOw5qMj+wG/me
DEYLPsZ1v/sXNyPMg9mIM91AMgyvs9N1bp2Q7IMFuZ8a85Bg7aJNmrUE51c6vJaQ
3YQFmPj6YG+iA9+HuwEkckpKYMj/VTD13EWKveGTMtLwlKpR0+HwbGWQ46FDP/wl
PyionhCjlv0WOe0PYO6cUmA4pe4ap7PlUWzj9brdxkj+Tt1bxeYMN3x77R2H/qRD
0HC0KZPoLkQNvCEXC93M31j4pNacRCSAVia/x88JLTnAaNL1KhbEGZonxmD/4FQq
L6sb+FcwEWhx0ZSKCAq4g6h50YAKsWPYfAKfcMU/49KjKFYZCZzIwAopvGsjkbkI
ojUEWUfHW2Pp4NtB9S7XrTO30bNlSP+5+ju3/Jr/rqGRm/apJNP+J6FyhxCs0PPJ
NJyM0a2Lh4VpZXFcO09VrmUtRKnxth9nf7dO9MDsU7FJ/0VV/4bbHxDmq6cqD7OV
cQmAhhuVxLg7VD8j2/z68GfV2NJUwYQ+tRDxgYwVK3dSN67nzsELQES2zg6zyB+8
wlvkv6kdRKj2DgEg3D0Vn+jhW8/JhFQ5JNJiZCMCIbA7MQpm0ZLHnzXhPNwgvcAj
wRH/Ah5g+JLRiVbodajtN09EiMpHV8/+JfVIkibK8oR/pABLvheFp5YIiuJpWq43
+SiavGOHdhxSQdZS45h5lP09cvuglX6r5HiwHiEAnPJeVKH4hU3yoCSKIZkKvefQ
yLFEAruiHBU/dXGxD/IMj08DE8d7/nJczm5bjT+VLqZfst3l1q6m1odkbYwamEpw
jr8fUK6d5trhV1DsreqxOZ5mQP8jKtS9GbW+fJ+QChNwnxNU/iPFv//yFxxUGGoC
axCvH5X6dxLq/QTMonKSzkA6PmpkD7dUJZTS63dyO/I3KS5HP9xUySVckxbgfRNL
2poM1MKkZyOkMwdMZnAqvN14+t6cfBudt1KeJntCTQJXQLUJEcvQjMq9EqMG+MwO
c1xoLA7zO/jh6k0DfzzdFFzu3M6Ba5APRuk949CFmLWaSdlqqU8R9fm/qc6EgIAb
+4LvLEHM4g2ViMeW9ptyiG4xJZRPdh6BSMnPZW6TLZ2824nzj+WxYcsRuTPAhxqA
f5XcGKCJ9KuJ7UagKrqDNC8SayD9tJORcM3qrTcPYFHlSPffdRkgWqszkD/BFrrP
NaYb5MyI3S6LR8bmT8MD928cQLKC+N0t/yM5IjxN1N4vw+AQVAYpiNAVSszxpIoX
lif+ruyNWs9glNfegkji6gEno5TrJ6yU3oM7+yM8gRRzRhYL7r/SMHAL8ks6YtNp
ZRhkrcQl5SB5aHxKWMwmz98nstyKrDUif2w8iPgUxpM+7fVbxy3C4f9ryOFrM69g
TvLlzC8WJE8JYt0OVppJgMwzqASURteyvhx0a/UXZXTFPsUpCzJvELS6ZCBQJW+7
fE4KpywwSQdGfjp8dACh8TMcsK0SAp3PXurhaQL+1h+3LMTUHUxkRQdNFp65CynQ
Bd/XvVbhjn5w56Tr2E0b0dfAYuO1/ZPwEK9qHWFNhVmZE4PeQiM+2rm83SRjlRD3
cMLIZRlmrGWp/8nCPh65bn4Rn/SdQGg5xozLkmaISlbkjPiI1O3la+HN74Hp0Xm3
i451gvge9YgnXcqMbmlvZ17h4lgiqSHTPDh7ylQ5GM4QVxde//Qv7/jzYBBOGEnl
oJ5cVir2DiLKhiG6Q/dIR67ABoi9gbKKkoN/lxFzgeFlh5jitPItW1r2e7WqG78P
ip9czyB820ynneJftpdWnGnV6k9R7RTRVrEgs2J8Ttk23ig2NF0Tsh42m2MnKPqb
81VZmsND0HEP8DrJ/ot8oFYsqHUoFwTk3ov0i3qNn62IhEotqtYbfCmncxiJ198s
u1bL5hZD1J6KVUE7MDYzyf0AD3Vw4YWM6dSpdC/sdBUuyQSa8lNBxddTqO0B/7xN
K7nJ8VGpYjmHoERvFlj/51+1jIvsjIRgZNZewRf0eYCfbNtjs/RwL1mkOxDQq3AE
NFR8iStM4rlWI/3G1L6st9ndNu+C6EoBDcwA435PtqltoOIuoNPtdqqwcOkfQcKK
thFzA+OImYaWS3Q3sBStxJOna5tP2dSD5lcJzqz8eP7Bmu0IftpLKNPwdrpkxOJD
+aGkv9eCp5m8UwObbbd6e4vt6iqwPhklTGUR7aU4Bf1zK7hX4YnPqc8dXGSCxtIN
GAdjMuAWu9BC9i43T3QdqZD6z0rk2eENzG9GJUdn/sY1rmmi6b0IOViR/0PJPKEz
ZSfsspvtNvDmQCeXvbX9aM2GiombGnKYwoUsGCW5RIT6Xmm0T6/59Tkll7y0gMxz
No6zq0HGlMgtVqcPV2HCW1SBOTO25yswj2P5VJkKAaT02QZSQFCnDXsBMCvioiol
76FfTVbhFv0Fi42Qw/J3o/BndVkLRHp+1lyhxmpcXiaSyNj6OlDK7ijigfxCgBXB
iZVh0oHDpQfbUcpURIsDWfk0JWrd1ObO6HJ1JEpwZTN1hlrKODQ+v8bfnQbEe7dO
/vZbpvKJK9wh6n/S/Vpac2FjlmG9huD883SmryTzwzNA/7TfBsM+c7+p8ylqBPCF
VZt5B0lmaVHakgr0o/exNfiCiATUucjNWkpJqj25l9BNvP/kKNpEKDJN3s3F5hH1
ZCoHsvBCVXAhrFyMX788k+BjSTdcbRIUZs7F4JfzRZDKcuCxE6Iv47RsI3RfJDiL
iC40xz2DpRam52jMhOUq6HkHRQnk6BQ5FphWNnhUs+U/+5Tjym5I0k0BRJ5VF3w5
7NhJYG+saYjq3gzL0w6TqCqyLx8zQwUpli6EJHNkNWTjrirT0cX3rOh0V/PJVLK4
2JddrrX5JurNCwoWD+XogHePH3IsxNRDgL/v9WprlQBvUe0K7+h5cT/sk7IwrZTZ
Mw1SoEWRvQ0tU9baR9Za4calb5kwI348OdsJVtUOl9T1fFEL21pXn69ssiyRBNA3
wAXlANBGAjiRP9KDJ8PDteh9iAtiDHd4tC598CxIJM2DFExSh7rdHpsY53DfCoCu
AyubDe5ElPlmkxmYyLb62rrtq8PTbkSsvVFg92Y10QYi98z0pC1qNzDam1tlLgbA
pdn2sdIgdjzdVjai7BxoW/9SHazEwFo+R3QOzr2kBImDUXVXrc0Ov5FwNvHvJ9t1
0ORpeW0kS8USgmywtc6Iipi+gHrzNWAniWOu5V2Tpc8CB4dlMspWPjfiTTQPmKtR
9pHmSBqdkPpOrKKKugEj6yMRRd0aTQLfQ9g/9OpXiB+7OO7orkaJ3UEqoRcKVuXD
bqqgO/ZiCG4mXXcXHrWJEemeDiR6dYq6497vMB/71s4uxAEJw8rlwVtMnRuhncyh
g/blHo8Ggh+OUdbm7qnRDVzyx7GSIgDyB6z3KkMvboRLLabR1o55TgwmW+OANp/n
lIswWG1QzA0z8z4MR+jgiH2xpcB/UUVYxoZPRuHWU2xsuBuCpfeQY8OFtHSsLFpz
Z85xOr1acXMO3rjigLsfeLJRUp6SW3ry0I3PIIwaypJ+d7CYhMDCzMBdpGekwe+2
KFBSo/F+AskCGNxo1JwSPbl7IjJsygKOrj440mVsU0t1L9JqQayTjvNgjw37QOjw
EAOaPa9sph8JAgDuTxmSRlVkdN5Ym8UIA3SNn9YQI3WbOw/8C/MTZDdfwxHoGM+n
Yb1Z9KdApOGXtVtU7aaUlcrzo2F6zeg2fChvTlGoymeHfV2tl5DCRTuRATE6GDMS
SrYk4hIsHy5ZEvXEVVa64XRkMihXQ+yiH9/M1YS6T8xma5QIoU5safIcEj9caX0D
BW10ZcNaTiBkfexiOe7TqwCKD9GTrupCUBgBE5s87BnJLCshlLSK0tbaIw2GTWPt
S/+t6Bqu+vodcZf8NYMy07lXBa3WR/dKMtsUL6oEwvnfpJ2amH2PsK4iICR7b+aY
trvKHDeFm4H8RagWYN3dieks0LJ7KCie7mRXcgR5ScQz4s9qf+ZswzJpd89TsRr+
V0t5v5vM7ZX0So2RmeOfwk2xUVYhHuSPTSbCGpmf9UrMKbBIEBnbn5B5WLb75UXJ
h2wJK7hhzlohO9oBPtoatep/dIffkn8LRNwmnMPkNXbagF+Jzc1Y1dBzFf3RNA5T
dhWNFA8xOVKF7C0SN3EYV2vGal7fiJGM3y88QFqXe+2kBDkIpr/a3yfui30ReI22
OqRM13Yrk5Jvr2S801C+th5U+L8wjlGBYK/w5M0a6SWKxxQy+rFXkIfs/lmY7nmc
ZxlhkENOsHjQfKJptAHgYYCneTgmHgcmmisxLSnuzd5ApLlmUII28iQJaeS4QbGb
gq21KM5ZBpkMcceJGOY+P0xXlirrZ3MIZ3j1KIqQlwbp1DM0/9Hzl9qqnGfYSvpo
LwabxMU8XgjIgti8/wLf5dJCV212ykLaDoWSiqlzEXFDeX6F+EWqlFimU7xOcpKH
XmM/tvwMxWN4CN87axbv4WL3o4Pg3kEeHHEdCmCpDMC5unQLeDl/OtLBDIGXyvTK
20KuEvoXDqWR42yapsNgTgZ5q1rPCSZ4MU9I8WWn8kKgZABrCVH/sQJpAX5uOgqZ
xD2ihq05sKywP2/36PLNTL+1YxAXaSEdpab0KxHCRtPFiGfpdy1fZyQfZJAxjLgb
35FuecJvBRKzwErzeYDMmrARulG840faIoLfSWwbfwB8SxCo14D9ZCIBzLyp4DJ/
uYxbGv4fpT19kj0QI903pXrCjMYWpr1z3QNRVZ2S7L/95+My/t4QmRQm9L8fFS7w
yM5XRSB08tAdGSenTrUjg2g8XxYR7ScL+rZZcvXiXQgGlXi+59hRWxKUH7nbTOch
aOFtweU7wOiGb2kF1ddm+6wwRVvSg0Jf+A1wi344MnXRC0fMzK5xnpBV+RXZoOOL
epAyB5VD1pj/PKN1OFrqz7X5COBs5lpW7ots56KilZ6bTJdOjWg6tw4SVRffsp45
tCVmBTr+05ula3zK7LuaJYMLY4safpsn1G/opCY/e6zVYJ3E/hmtKshhH5wWo89q
zE5kskCuSmaDklqjWadqcuj+US2utmihZ02jI0/8MOBMAChbdzLkKHOy/S8RvyX1
twCAVyZpgj66Yv/B70BzMJf4N0nGb5Xd4LKK+3vMXS1ou5Sli8+1ESNVSelMufJ7
dWnyFDKH8HyupcV921pnZSyc0w1+J2MpcB8W5YAZQxBkxfm9TX5MBcjjpW3SOtMQ
xmgKcIRR507zF7haCAtWcYsOkfu/ny8unWDalyunlbK5uQPuvCsxssr/wdMEJSqh
ND6j8bSO8HVi0GlyaKFzz/d4V1BJFdb+51zS9QuXjjHJ8SvBkYfRlTu1Hyd7dPg6
Tri7cfn6oNMcxhCnc9+i+iPUuGW035Ta2XA3Y2KakFrXcmqYT13xhPHlC4IaFX4s
2Vsz2pcnRGH99WkP0dDJ40vlU+4glWLR3hF8jbSvwdcmuzFuv7x5EnwgYmbDLIK9
uzgcBuuG6WA4ql7q8WyHHRT1qSknaVWGCX2D5etVE1Q+/2CIpaKUBMSJ/RMOaLjJ
KemiUFqKc+yYYHy+2x2s6mYvMXecVNPzSLdv15T5URyI6uL7RiyI6/GbnqsUWPqt
ahkOyS0OsEB5RbLdiWqFgavusApkBJI3ke7qqUmGTDZadhyX3koxoR5twHkLWtHn
hrQ7fiH+iTKL/D2Iy6dXp5FQ9R5ZLIoItf7svGTtAeVwFg0thOawDWQS4NGAw5WU
1vFGpWZXHmB8mEfJbR7Dmm694HTnZQl3mknf/VYJNwugOJ50czJKJwwm8d81OebY
CtqSAjopSlmvWfng+CK26xYlowC/sjzx4WikQioAqC7Dve1kwbGHR5F1ABeC2x1T
m+FTxxYOLC751HSTkiWyKhnyh7lRtOFiI4EKawg42nCieb/+ZeeNdg1DoVkQglQb
DCtdjSwBGm41bA1HSbmiPEvEZDSSFxu/9hCKxwuo1JH5w5iqT8ibkqDgkqK29HVg
ayHsH7yvt0vN7xkl/TbqyR4gt37mfk0v9C7g2p5XmOutmcH8Li+qMelez/qJaH4a
rG8It8kZKHlAISZPxraINSBPALQKvNdVEq7ye+Qen17n86bUYprIn0ULOqr359P2
ohZWswFipaokM9+DXfLaKkpRtgpu+rwDKKDGyk3/q1fzrocLF+ttvO+TS/Mt1qca
UNim5IJEbQ4s60jESpThphbJM3rV2hRceiTmV+TE9URNkk9rHVxtekypIFnaI3jc
e2nP442dqhNmRU3b5PPAccX/EmjadZdmO/eO4fMoehhGc3nYV8Fz+h7jwVnFMYaI
hjKEOtzxzs1/L+pwLiSPmyXPxgF38Qd9VdOoWK3+glxKNUWqtOftb1o+Dy1Iz2NM
wwwNS2pN0l4/nsnELmtbE8vieaXLPAwc9A3Riz5CFlv/Y/fmBstHfzZL1xqtYgYF
2Zfo7EcxRzLRTXt/tHszK3nOe1ggAPRWfoeENvdoMrlRz+9zfstUFPVPGOhUzPDf
0OuFonPzn9Iv2HQ+YtAZ0bP+mDY1Iz9b3w6+JbezpovevPlaq/dvuUaVqhYIvJuv
MIj74umrwJ9mik9wUd3oVIL6ZAzBF6N2qSAi02xe9g3EcSbnppanvP+msGGNspti
X9nnd6jAkHCqkHsLeXsjvBO/oIb4Gb4go6OXkBBac1LgnrcNyI48tPpYb5/vRrdf
t4cvPEe1qu/R2iSaW33Bf7HZQx25BSzuYZmSrvfh9TjeGRnU2ZGrFoxRou3TTaq7
azzWWYxvJN526eVGUH1hVjgHQr4WpkDVkfIQc6VUT7W9/SJKgYUm5SMkpHvR/H+q
X1Gd73VH2Dy0iNUrAAeBPAk1LiohBOXifOCXK6b+q+eGmW1ov1FwO698ltCQi7cQ
hD8tBjnttlws0FbwPFH0MDgnRsdhbH2A13ppFYRELz8osfGz+aHuyq73qdE3wJmK
CLy8Le9jA7slk3mh+IVYX0HNOO2/pL+oEAPKUgswgNHNf4l8KiKwajCyYJ4I6WPt
Z8vBDnpJVqkBfCsMJFJelaC9OwnSHT2Z8uJXLr/h5m83RiyYldPuvlMvWMfO6NKl
C0MxewADKq6Z99QEw6kUHPS64gQsdD5dQS5ET+rQH7mrOjNWwjj0rFur7uHIr9OJ
S0CzSaDRmkVrraW8f1/lwLSspOgtfH0Mp6GP73SoyuhAEZ0PfP92S789O1thH9ap
x3OI3Yza1hOrJgDKm2PuyZB+m1jAlq/iEMsMsNtUOGnN6B2zYryiWFnPbSaP/UFj
dk3rqJTbrRcE7cU5cKSElqlmhkMtJ67IT5HHOcslqLtkASTGYrWgf8pKsc7YPNwY
fnvWg1Q+vn/Il9kcVMAsPPHddA848z+iOzyU1xyTvKDa2xZp0iLGLovpL/fJXaoZ
6Jp9gfwdaTAB2ef6kJRrIdcd0piZO3/8PWIaB0mhVUlnDK5Knj8qkQZN0bwVbCTZ
WZj440ZxzUpdemVggcUApt+jC3GawhdBrtcSS2DCfUWwqDvIKc78b1wKzWExZGCi
d2pjqaUv4gJIPg5kiiKxl/7poa64ZAc9rvGuK2iQ3xDw1ExGjVvlm/Oi8bi2hl2S
OIebZtNduBhtVSZu8eSyzcoTCrk0tzoJmsrdApG20ewH+JqvKuk0vheizuQ2mILL
ud6fXIjNUM1h5B8EhPyGsgN+IAOQgCby599AK2bYZkL2Adp/o0f3FVWod3ukzf9A
3+3UdlYmgt5PWMlWWoJWPidrEDGa1PPCaWEtY2DeeuYWB18DJoiA0BhEEtwLT0Hk
0QwXpc8uC141SRqTWfdpWzJj3Odl4NQ2w0l7gJ+rmCdr5cD78uAdq1GNBVuh3STo
yJ3D9ERrNnuL4AHP7Pv0YnpVUQIJ6MIit5uIXc1DdLPaMlAa2Tzr1uQbsWnTMcV9
GuAVacLlNc9jDsl9WPhWhqssJodlR5qj7DkJev24fP8DYx2ivaDcBpZ6IuATigtt
wBLv81e7lEgiIoebdHWgPfJKgYyqS627FtKPoqxgP2WM/P5M/fFsY/aVndHi75oo
lLRs9K72L5ub3KdnjErFC+QidBS0jtlVpuKcFWVMf2ABPqdSPWY+z0wLRkY1W4TZ
t25ho5pXaYLK3W0NntTPzGqLsNkjwJRhW8pM58CpgRTyS0o8rBIwTnmSYQXBq8XZ
6+CNjjbZQzpB3ta5CbtNBsAQDxcDGtZiXDQh+LQa0YSnMhJkPK7tT/jgMsrW+JSc
WavSj+Wpy/cwUgreS5nU3PEWp0z4QSucaTU6XGpFJTxt04/vZBJsOT6XThOcxr2N
umfDllHBGTr8T+/SWsOHf6SSq2ZNONISQMgPsQSKP4H1WuLIJPbA5avRk7SeDDTI
z/qESW4trTG1PRBe+hmmjjmN0UDTKk6+qOkPA9lMyFEy1vWO36Q24Znj4SY7Etay
kIDQGFl1TWWETCJdlKLn8RCFR+UkgY4ka/s3X5AUn8O2cHpWZe1Qihw1JvEsM1F8
6Bwb/Qo1J/lNfHUOhlPuP74fyFsdis8VUjcWU9gQkyRsyVecui7eLRRuLzG0lfuk
UFrEJ/T/e2QR/eG1qd9iAkWg0Tl8FIE1SHb6whFQ1QRcg0iFTitvazEVHWL9FBwt
MaKttRjhz5+Oyz41kglcN4/R8koqy3ID0EhwwxsZNh5qOYi3JgynYT9UaGPawluh
PCzWtp1f8Kc2ZP1p7LSbM7orgyUlfrzvbpHi4FI2Mq3CVhC5Rj/8zW3zLxzlbv1n
qEl+wa4XZph81PjugXyPsKxcSzQBSA98oyOVhsOjYAnPLSLqh/Imf/d/EqFAEh0s
HJOjVzk3iFSXlT3LywBGelZbMsOca4aAZ3vekxFHOZGk7AHQHK9D+OD1PmWeBeYW
KPWRbD78wRcbVzTSm461PuvVwDeABux4OGQIQsy5pu4VdMeytzb8qMalUXWmTbzp
zm5Y1WW57tYfo0CaSoi8e/xVDOSdrYsPgGI2HdagnjrF2vdLnVJZiZ9sMro+Eih1
OjZCXmO20fVIVM3Sw/0U2gdCCIEEltNZFOAHEdoldbxRA2QchfccDg2yJibA03Fn
K7LT/2op9/YP43hooZo/W9KN8JBIvoC2bXnxTKfXlxlTFXM9RSGCVGlPA6tcngCF
3iGy4s6TsQO6SDCz++XiD/mOwuuyRSVzp0bi+9fcEB9g0PM/cA7yY1UsaQpnQ4o2
vceW2s94LyPO59NVq/DjJv8Iqlgml+svZ0j4+AwPVWXClMH5CrPngeLeKznfy4OR
BY7BZV/w0SZKhQEfZD83DOWozVipThVYjk2SJR31EiqcQWF0KQ4hscfrCJkaJiRF
kZXe0HMN2O52WbvPTLAkHHQzKut3IYtJ952MkY0D+6NFcyXWdVBgULu4BlHB+Za2
WDxeCKGfCiJlWYyKGzR6MMrxJZmXY+PGHQeNXXauuYfzfLG0VWdBJuWY3oNww5yZ
pXnQcj8Jh7tKPYDZv5E3WWFNX9EfdMLHTetLhTW3WlWHzaiY9Zf5NyFniO1oncSs
lsZW9iKDOS1QBY3TVqft1eOCq1LtH5i1J0B5WhuGd6rIgolbc1J4mt6//HpkrOq9
DSsW+UyWIG/AS/vykOQ1hsb5g7GNzPGcQc9P7NqB7DwQRBJIsBrcql/We7XI4Ein
0g7+ICUzpb0oumdaFlvBYKm2oxxlB4Gc5Y+WRBdzqknQKryEYiQYNjuHntYjoFIw
Cd+GpGgULeTpJhrG191teL0oP/gs4IwN41PF6DWdObpvVnseZLaaOb+iBp0gdNK9
oWLKg2WlOtejF0CGaGSCBFFoFxWzpwZpQXFKxZk/fjXjbIsCv46BAVjFdTRPj3iZ
95f7CMmOX/mDN+RFJQqnA4ksPs3mwGgIt3mZRgj/GEoUllv7zwuOGjg00zO0/zIo
JJlUiLKaPvuxMSwQxO8PdJ6Xv8x12KQRvL1QMIMYHI67W3EmhY+r1+KVTJkJ30e8
d7CbVXNKYSlCiFiR1MuA9ikN0wzGez7c28Z1TJwIfElHLqsSXorOQ10CEy26HkHn
Rrdl+X9XBYAsm4qQ+vax2iRzbQexSoWVBHA9eWFPboPaiOpSi1+45UFsUewpFs5v
lLzVDs01EaWbWHXtog3EuJPXDV1LWh98nrwBi4ALRY44Upm3Xjrh+0bQ14tY/HYF
Bu0jI6ozhIgpfswUxpSuTXCS1isaWe3f6f96I9sN1ASPLQqWNL+1gU8wbMpRbPVY
bHlQmCx04c4cpRw0UsL9YxUZ8ck2bELaZcFUMXKgv/kG1j8/XWApEKYnzuj1EkoD
WFmhK+9lUVZfqhjGWomB9SFD5B2QDk3y3eBIcZ7BBgZcAT2lkzEAgMTUXciLvqoo
ajhRSbYt3oWRHK6yeftgXfrzx+FIfDVZQJ7Q25dnEf5Zxa3TbrFAoRHzOopakVCq
RQtYsUKDUMKlmjFbsMyOi6kNAJZr908YJWcYZ27sfM98MPpU5BaDsZRGJ6ysj/ha
qEXETgDoHc1xA3mrvzA256aBi7XCk8Q+dL8brosSDXxnBrED8roy5lVSIrKvDvOo
VAnrrQmni5Q5r6guDoYVL4AXiIAlmXAyusJp3RPG811cVbIpDpSfC+e9nsKMEWVx
CP3XXC71SmxzZ0vn2fq2/SLStjMa2laBZrmqGhx3dt3/KcarDjZS1BW2dzSR8hwE
VVP745WYhaAF0N1N8zy8rDWQ+hZHJ63nkK1p85o4ImS5+niPoRjD47aqYErot12H
G2Jn4OdVpWwECVN/ufeubzWWJ0pQo2mkevBOBTje92g9MImyBbfVo5IXVvJUQvsF
PceSLYGN3V00RN0RJFfzAWg+pPh/ZcUyhpbp4EtxqIovh+NN5PYksZU0GEyW35XD
r5tmo1WUO6vnxrHqst2EkiQsg21sn8/kSBguzrM4WtzExVJp8FnC+a6iw/UW8rSg
HXTNzQ3bPJFkgHaf4sdmczE5/ny+XYkZlYyaAJo/QVhp7ZIGK134iPkLNmaX96zv
B68eXrfkyi8/1I6cdhCv+YupU/s8hWvQoIZfiRgoe3hErFRqcGCcwMC0mrW05QHJ
mSI3mwgUeSwoEIZRNsoF2Ktxp2Czz6z4+rDgq8vFONkSJc1TYgG71pM+VkeglPw3
N/4YZBk87vdTbFRulqJWTbrUu/Sj1LcqSUHWx8uuIDBko0Lh+DpF3x7ksl6/EYRI
Oi6T6l+MNENMBfFMhLEo+nAx34+zXTLYerK3iChuEbygdKz5nb5b6dB6wdCfVBbr
wENCFhKkAZCDy5mfBhCArCt0sFih2nPxPVxWrA+qcgUDnrXNEkpafAvblR4MC+vh
dXqJVmGHvXBFWMXX+3oWZGEiNlvM6OKaObvlmdOE4v4Zx5b/KrqE7mCHltZywFcP
B3m97OM5vE/9TzbO+XLzgGe7gf12zvKdZ4sKWBaAyde31n0t2YvzEc5tc/0rUO5r
YlusthW5xzYkGpM+6/kCBFdbfZtCHIQMo9M8i4DtWpWM8lKc5nxydXzQcrslM7rs
mY04Mba+v3hHrEavGAmsR/qHOhKlvdHDONuFUDyIGwT9hg1HvorxJ54yF76cUpPf
ezRPWUfLI/UlQn6tk4PCbOUyFVa9oE7qoDM8h6QHLhV19oSrQwmsxjePbeBTYn0l
MQM0pdxdTkpq6Q0twJ1XuuEwg2CygTGKGPfEvUnkoZA1k41ptxENGTA+w19tZ/MM
HZG1GS9iJ6i/KcperAhqOqnTsaS7zdRwZdab9ihK/dmKznFT2f/6biV1Lo6yZW0e
vAxCJL9pDU3FCm3b79+CRkByd8TARLPFRMeefAH0D2Uaj+z5LcGWSMLcOYal8l+O
mzHd71B2yjkXBgUKHh1PDJq/x2aEjdN7jFus4+JkRtKlcmSpUygHiGJ9mbPffqi8
zpyd0n/Ue7wCBueFwrIbFhln8w/yu7/bjLx4jV3S/Mr7PUjAVuHAi9Y7sJzSat5f
W1aUG2B+/iFViaRUohqb92qMW0odX0s8jHaIGrO33oHCY/XfxslXVMiQUn7bnsVI
tEi2gz29/riYJh/U7HHtCrK3BkM23yGMlKB2GT2PqoBvhCOkd2aoIPbL+1LqTxOw
U9nvyOsh5I/9OO1XMB0jaExcRRgyYNgSYYRTB0lkNSXM0ogeVS7D136HHu+eOObA
+BJvmSfA+slTEeOeDPPm8fyUWNHoYVwDvNaDNzOxhIPttAiK4DKcmGWTdJNDlJXJ
1F8zngRKsT4vzPizs0MjNUHaFmG/zf8U4mjKukAimcul8dWJMa5bHHbxlPr94jUh
6okPfcwiG6u9H6uf6R8I/De6RgPt/UMflTOP9gE6pEcqiJNOltibF/H/i2ryO3Lg
nF3N7vtNrXKiWsPcJGrseiFo3229JXAi0fDj2FAen5e1847l1cU4fixKFTLdyjUA
Q3XNSxjewN3Z380kJnjkYNujb84SbnF2AZa4D8HFJbAUZzK4IJlagi07qoQKBK20
AssmVeRNtTbY15elK+mvvr3mN2juw2zLiPK42zQ/U3baCmyUwSNyEkLXPYD3AMMG
fex9rkN87Xwp+OdgIhHYGD37D1S4RsmdTtsCqD85Xj1gMd+nCCOcbapZj0RHhP/9
Dt+TagcME4vzXbgsw9Pw24d/Vj+QbqRJfJGKadgzPZOeeTWGQ6IabZ4VevikTGRK
v3HH1xSBfJSxNkTOB+oMD3vEwRYZJQdM7h0W9GgXy62oPM/z/8+EINwPE1U0LvK0
ILLb6ygFUcl/tDRj3c2MvoB0J6CZSJO0k3Poyzx6FEUFtO2jIld1DJbRt/+bMDx6
CzX8411RiY1Gnys5ID8YNLU7IhhPL0R+L5V41+8M+RIY1Cg7kS3zhC+EQwI8u3Vq
6fWPdscMMaBn3cl1Ib7JOd0rddkjBwotaR8O8weQWvI8xDX0UtGl4M4nB3VF2TZL
Dd2NTebsaV0C6gSnjgtxAUngsmS8feflrSl590Bwq/QM9vVnUBAgcFxcf2m2jkM7
IbHjh42zdBGv4pwHFjZL3ajx0/T+/cq+qi+zU6dzdZOV29BeB3ROes82sFY8Rldw
edh2VZ9VLdhmTwi3y5TWcWYJpTk4DWhAFvCVz8wJ3/4dYG445ieQDm9QvxAYI8ld
HIMMlj7PHHjJo5/tHQp7ImneGyQn1+2GmNm3vmqR6neWJttbYXt5SvgbOzDfl8OR
2GEImH2UOUYF+DSi/CiKbQnbXggVdEdimIV4eu3aJv2n0GvmMmXP8eGCAOCX3DW0
LuYsR79TfMMKZI2PmWwmETC6yzLf99/hc0fIAiyMUpNcafM9hSIziVK6SSHEPj8t
XZErpgFnEVL+4lNN122j9BkfroqSZfIClZfxydtnhE9uzNjyy5cZ0c4QMpY59V4i
GC0NfsMLrEhhkI3N9Oh0/3h2mF/lCUtkTww1dy1Eqq7K2MSbqxzvYsMSKEmjmgso
+qXxqUa1m+EVePOIhUXZDJWxP5YF1s92qZbn7DXrwRcwYaxo3434lQ50smzQmeyB
IdJULaljgKM6C6dKbfJZVYHambH1ziC2g/sbLEcrKfA6o8RSj9Cub0GDLNuGfhPu
NY0HdtBp6fz83EePka4gHFZgtc/rLFBAFjhIV68uSd4BLY2wI5D3v7o3hLv6EvKS
gPxBKWA37Jt4gtLPfvp+wQ+anIxvApNwHaO5JI7AqNqEUwE/O2ktNNhMuw1xwzEU
0beHA7c61H1/DZCkex3p72NXcIhtRh2UY1inGEPPdT1psyKbBFk08MKb0kRb3cgY
+lcN46sOYA/5f7/6QhCApK3cByx57vz4mDlQ/71jff95GdD2929vSJZSPrdflyos
H6w5ETHUD0OL1lY4lQsZiezybtK+l3BEFJjAs4F7S6zXElni7J69WLCJsgAHr10C
fZ2UK+BH/4uL4n6hF/SShgA6IGPbwIunnDaSCAZ+mrWEQqFT9ZCN68NS96ZDQCaB
oZRNLwqKrhZ3Bfu9SCj5+8MxOQ6LPHYiB9lc10yHqc3LpIvy66H1WTemY9PUByIs
tMlElkv2bKvaKCri4HWElfU7bWnsqw2UxGTpi4Lx/YjnumwTIyT8efuAjFMsFzi2
o8AQqN/B2qq6uznn51XQ2DWX30v9Dhb00zpyg5m05EcO/VqSwUwfiWZRV7CJON4H
7aKs9Udlh8SikFHbXjV0pCjYwnJ57/LhJWHAoW0IU7+ynmKhDtuDp4VMgMNPLXLT
iqiTtmHAHnSFGD3coaKxx1l4kAOVW3wdZSAv+lI6tlGJXMleBuS4Yhajtyh98MPU
kOnL4bl/1bgWsME4BySW86332WTbnjHltykOJ0Cn8glP/VBUAGaff/Y65CbOrKCe
rynu0hQlbZuorCVgIuHrOugGSPJB5owh2rhhlY6kSd5VsrVCAhco25WzWXB5ZkHS
OqomlZDmRHN46Vvdexc0KyxlNUyQW/E9voyaIo0MgmZe2dRm/NDK93jHXKbgCYmK
UgxRFg4n+uvI/B844EdDxDrXakGL/MHFZPUmAsCjP8C44a60Njo7OOqWqzkjdilC
ZDM8IflpQv2XaNUcX8KR1KTt0jClva11eMhPCT6mFs3Llfzvuz3SUJPjtuYIqcQF
uhqzANfsUnEgBrzyCHZ8uUhluP5xyAqj+Z6CLJ9oEmSnbvvMbpRJIFz2g/CJspoL
aVq8lCAFIyHx/FGRRewODpRpf/o6CEeHLb+vp9rVVnAPIKBV3y6L6Hk52dREIbbM
tm0E550XVnHF/HwlSKHmVHXehBlFAFrGanMrpc40sbhZgOM2ZvDntSiXEeM+NN54
3UuXbgJoYD+C3LckAsslsrZTgy0yYKps0drHccRBg5ZjXHGvpYHkAIkXJQ7VAZ+y
UmtLZAd8eHvnUwp4TA93G1oeOnLBKitFF+vIAdMdpE69U0V/HRExBhxcndDRexr+
mlyyO6oLL3FTw/v+FSw1KY8NcA5keocMkW1OwehZQnS0kywRFCOJXb2nEy6GAMuq
Rq7SHvWnxGisBhBwhX6zpx35FgaN/zPScRlHL9ZPMG3pV1g8AeBeeZbfhx5UFT9v
ryuSwC4Ajm+kWjq+CMB2JL5FsiK4g/+pnRo2mTLT5HK/dTgVHlfAhdqDaENKA4r8
b3OUHflBbPtZ6nqffw8SvkpFcWJueU++OYCin0VWx9Iid5YVYGos1IsM1odR7pIG
bGUDW7a45zl28jXayUKwl7LaL2ElJwBbc9scn8XVosDyzuHBsoVAKYKwo0wVF+9k
7LdYpGUvBCLVaUkcWmf9MGtjMLHzvMZNnc1UWGePgcxiGUU5GaRXJNXXKIx+4OlJ
GdYHPrBpIhbMybQs3ScsmGaofOZDnatm9ptam5RWKVV4Rl+5OWEgANSn0xiYVm7A
bczjG1iFtJuv3oPTB30OlASo2weYs5j6mo3Xgs4tI4B1Ja+FR+xqgVBZk0s3eLWq
9lwxTFMFkJbdJtPIpES6fGSDSc9hJq6B0JIdq/g3AQHU1eMCEnvpYGQsScJDo3CH
ONDnu6dKOxoOEDxI03HUtZq+udExKHcw7RafYhRBV72uRzu3LqyEn/g0oMeIsnEG
Jtx0F2lPvvjT1QhwNPLKe5B+K6A1iySfZcC6LLhtD/5PhQCqLEorJ8WgoHzfb/kD
G6Bl6pEOb4cxKXt8osMQ6Z3T7dMLwm+xytfXoNJNMtgpDNgYiodvFlla4gkmiNX+
S0dphguUeXIWvL3x1LU3law0KtNZas5ztF9DgwgWREl30iTXsBQZ9nBKbmoJR4fy
81/LbeVeDWYQfMz8O1TN/3OUc3IhQYi5/4oO/J2BC0rjKi15q9Lniu091tuQkzBV
cNAgSY7knFXoyHiNCvYu0Cajh9NDEIEaXSmVxL8n1QkxOAC2XtG51CccC0Su4VhM
h3GxNTxRtt9H6pa3uKBqGjNlkU/8tlBTVNfjkh+5aiT2X0SQ/AdMqqGIuBxw5XCF
9yGwBwVhCS1tpv6Vkr5udEaJCkjBjec5W82hW4ca1XtrY6pSNyDCbLuuNsaVaP7F
7G4Qy2bxbhahBjKYDxdowrMWu4JO7nb022jWWKf1nzWGGYaqTV696fWf3xLDPHqh
HT+ypKT0+jlRRAM8xZvqrCbHJl89GN1m6uEpoU07gEbM3EyiFeKSCEE6fvIhsnmh
oSDHzHwJc0MpkoAyvhiT4u9iEcI7oIhjVckVGsqpk44mckKDLQ3mhx3z7Fm5OPvN
E8Hp8ZcbEj0HdYqtE5rYTzFFzRMNb2qgVSICy0aWbejE5X5nu4xyGJEWrL5y8aAt
PZR23CeP3bIpO+qRO7S7prCJnIXzOUqvQ1STq5uQ2+CBa8CnIptgzvyLr7mlTH+N
71NdCm9rg5tvkmwPu6GEQ9ZqBOlF0sfKicStN9PRdjw4/dNDlKCV1ajAP0b1EPDv
bcNOPYU8upwCz8YQUiuN9YwRl1rhuZeFtqsh3+iKhkPPRnG8D3XJzmsoHFnnnZhn
HBNdnQJF0gc9LlXwiU8L/xkCgpxkYSt0EPY2/2S1y6JN8MHLZHxAbd98zKhoP1/6
69kQhangBwPI/qpBR3xMxovnjrYwkR61g+KQGo9tQkkpsZmNap4ioJFHIAyOvyhi
YbnQ5SqJjGXTheVWV8f1h+3WChVOt3tIUxLmk9ls21MOoXl03eQudnXY3thxcwiO
d6fSQybS7/CzKGlSPQxrzwIAZtc7yMkLmbS5u9ZrE4s7xV8jTxssNjxHiavFlbRP
G3AyTnAUVynu4HkeYZxgW5O5t3FKu3bjeyirLDDlYb1Otqj/C9g8qL78vxqRlSCZ
ZM233l9b1BADfptnXomLlo0ahp/7/RJHVgIqunTWdbBKCOF2mJGJU0E1bE0lLxW+
FgWO0MLU9YfZxECXF40Q5crrL46xurFsfWeDpcixtXPnUaQutVhvrvBzCG18d4kK
j0RZI8cr1nnF3n8sH2TimPsrg6nx22xFEI4Mvgjdym3iyd4BtFsHIS4N43ASkL2U
stqV1ttuiUiL2FdWdY+TRybUOO5nRh532SDoZgBfSnHdm33nNhLKvlub3Xd0HJWd
BNGhFekTbCuJLmGqVFnHeRKDkTnMji/do6mJC4RtpGQarfN7VOfbY9OxpGHjf3A1
gjaMmAQhvq7rs+Efq1/RYEwukGCKoAQF8RzQc0kNlTOz0fsVyr3m46yYP90Jjt22
RzWtmHpyuDwxFjJjgE6dLh1Ou+aFFHAgS3gi6ujOcnM8nm+yMhWGZX2G8j+RXvX7
Xpy97ZO/TrCB+Aw2NYIBRVJwYlwx0vb6mf7DyZBgeTjFnUXn5rR7YBYzZcDQ0+Um
FuOBwUwl2gLy+grTcc3u30OuAT1TpYPwjQTD3ITlgmdoq79Lawc/OrCWLhzFRcx0
NZF9scWYs879vijwwOlvzJnlz57Vcf/McgkWQtIEzv7pkIwp0aSw1FCemOMDWIKo
C2XkQBCJmcr4KbSNXsatd7O+p7jI03cEPaE5hlfHbLroh4yg7IKn57jXX7sSKgJO
QerhOFa91WeL7AsUvnxoBXZKsVj6DBJ4qjigHHDFQPWjsdrt4aD7RiIDIuAl7Txn
BUsqM4hI4bXwBpecqlNR8KAeJpn3fUBtDif0Q5N+2uym5w83bUvBkyrNdSLO1aUE
uS5agNeCqwudMHEYkOdcsIHu57How6+8TcmkXEX/8f0bs4obKANGmifjktRamc/G
T6tvh7nKr3aM4mhxvJ0MgpsHMyfnosDERcgtgZhyXAP2A5BBa1CTEX3nGdvP0H0l
VcVfnqomTyZDakK31DEkMd1Ek91Wep8+PH08CIw2XA6MA5lGiRC0xClbqoNcCx3R
eWFhdlFz9SgO4CEdGKxM4NdoYc9QmKTehFkmG79k6JYesVMgG9/09sYU7GezexUL
vClfKtUufmQNE1S1vL9MAaKljnSYuzYAYGffbh1HhXmiwzYtpcN9pb26DgyOsZuM
IUc4o/atk8yjfJDvZKRPwYuUV7GlZRE/VOETcvLX8vT9mBYcmkxrYvunD5JYUh5E
kOInbfGjLcV+ulEhKe+V1cRckk1g2/O597Fi0vhFrUKEPZq2VKGa+ioR4SNc514r
3v5flzhGNY2EXirNm6G8oCfdW12iaoXiG0b9QTBKScrCJnIhjNoZkd5Aq/NM5ER0
Rcx/FM51TQGeZHv5OKvwHCfTlqbvYy2cd6UhjOm4cbFJLQzNWFhxCIr7GRK81PFg
bqvOdOyAg+dGqSR+ASEoKinOIrvldXd2DmLBJPUcIh5FQvVsj5ulDJjpALkvsFC0
pSZ2aHm9A1bA4ag3DzgCygieBE1e6cFVrjjRKiUYZh7vm5PTdB7y61NUhOGukUml
yBiW7I510l5lsm7uWBuk82YXv9pzOqcdMvAXTLQBakPCh+87CZ71/OCtGM2M8w1k
yeWNFlra7Hu07cTYU172e6Dadh1ncfXU8CXxWjFtskkbwQvOZTHPei5kQ+e4vrha
SHtQHiJP6BzgHyBVt4nYXSl7U883oYJxyBFwp4XUXCldFyFPCs5THls0anJoy3EX
dmPMWFsA3ZK6cc3ERDfLgGktvRJMo0JtcreK5GVqL32IG3fgAjhvcPjkBJVqq7hb
dtHsx/e63rwYDVP1rCRplDxnNdcj84MAgBq2HfJwpc/lCieSabxMqBDUGS8gra/i
337Ty9qTiISoWg+s53Zkbot9Dd+Y+Roh+u+z00stdd40USJYH0o+a7TnsjcAIBf0
SuJWtgiyYQ8FOoYn6PIY/rkHlK41hK5xyrmYmciiaHyMOBjq5L5aS1bYH7Owv/7S
ihlPZWyhbDOL3TqVoj10AOFmGktuzAq8Tpi2cH4P8IdGVbfdxgOLgCSEQbHxjJSx
iIKeqX5SwQnLmR6ZncfdCm6v/eGbJwfHpDS9jZmHWx/n2gIMJZKZIlpvqr4ujU1A
016q9zywR3RdfPAwVp6api4maf1i/zfe5Q+Zb+I7p0eSttj++1ertpYRDaN4RhrM
c2Vg3va5MbG3lzV/exhT2cRI/37V+yv0FfRewJgJxzZHAQJ8/M5QFYA7FORxmdQ7
IZCLtwMSsdRx0YkcUjQ6+BKqf9FfZIv9XoyeLYZud0vdbMLCWLszQpv31qS1AKqb
fFww2tLZxQUG1geznI1rQXFsjIdv4PHumiTgCWPhaYl1RHMslKxo7ZcSC5FNIKJp
Qokt2WQz0MghuxVFhO/AkaqOcmjvFfZdoKeO8ergfvLRVvXPbmZz5IMwJAZUEWJ0
c84ceYcgIIQOTaDUCD1WCjl98u9o7Z+rliEps9WzyZH3gpCYn4y6l80iWcNBMn77
RTV8jWRjLixZUpNZ0cP5q7GsvHsj8645f+gMqGqYKcPqJEbpj4H8/yeafVmpgDnn
EquUc9fiJkFmaW7JuiU1m1j2rI6xNABltjCjp+bnb0DB3kBmPbl/nyjiTyIogVrg
9gmglKHClqncKHihv2ehqUMHora9X/tSXj+luC5mbD53C9CmZOoeu98yNHI0vG0G
Qh4n9YM1WidaXBFK+KKgUcjUj95qCp+UmtHRwDX9mfxAmX/UfEPunlHKAeYUEOXk
LNm+9olvZFvIwaStXl/KukZvLbauuo+ZcMKn5QKisamBkOTAQ6ivXN9nIatP8o2c
fwXjpQKF2Rhuwr8nOrf1LXD/EoY0hGvEP4/1zie5plkpha+jkERRnBzWcyRROusF
PXLYbzCoTPrJuwLseGSCskattWubHeJVmrS3k9lj4q5vcYjuQEevJ7qiT6wwvtQm
kURCWoXLx6Wm/cDCH4jOXjbol7mgnUl1CLj/we30g4G8bB2n4BujKtiwFafI99Bc
kOqCJ7V8R/lQCHUHy1tA2SEKzJ6VFZiZ+QzpISZdIsTveN/lQibEL7benJY4hu69
hIkqPhvEbxuRz4HTjAPCgPWDKtjr79lceyNKbEhGMXT2HE5nHybQRNNQL1ENjAXC
qs3QSer+cd0WTiFoIPYjt2EKkvsr4cajI/eEX/Tp/LW0acR7o3l1YtR4vRcEM+Vi
iSjYOKvsfrSDcu7a4wMoCESUlYJ8TicTm8FmhmLFd4+uc6LwQ47O4hUvco3SG7dM
1HTmiklNDr2/vjLi6vLLtoXjc6fE9bnWSZgFG/QpHpcc7gkKt7wst+kTS5yfHUnp
F7yrNhOju3XzamyTKOht2ViQXjNNWvmHy4B6w/ahwG5F9qCLmoHLCy/wC3o/oxWX
hUZjtNfv6MJuotdFzTxmNvujbfgH5XSRNaJkDcrtAa2367KVjArageU/ocPaWGwp
0fzdB472thebP+yYFDIxc1ApEKTCI2hBU+rru1Mf5aV1+bx12+y7Ek7k80oCh+ti
1QUu3ugCsogOzJOLbFS36HQWCJKhZHQhOFpZ/bElJ8d9OO69BFezs5btdJUDcE6Z
p4Koz0NahD+1tTuo/UxCHf9V6PQlaDGXI+wuOgwrRkFiAFcv8seY3ODTOd2FT2Ys
u52jEp6b5V2IzPCn8Tdz6cHZYJPjJ4eYhHCp4oBPotRMPTIrxSUYj/bzXU41RWCH
JmxqZJNCjgXuznI6qK4eC4pkNUADiubu3vcZzVok31CjOUr2HyHiGk2vM+kvavhG
6IL1yZHqAjhDA5qfWYIiqjfsZ3bsPa2jDfC/dxSY8fnAXAUjXptEwI2Fv9iz2D+T
PuXQcmuIgeKRljOI2SnIiUAdkleQrDdgBqcy72CPbsdwo9C8391uc91GKJ5MqAKS
PgHvcem6WRwUa5rgfFwwaNwZWp+3tC0XH3YhWo/XA+t39cs7nisU5cVoH0DTqfGb
cP+av1+Gp5Bfjf1fQMn4cMjTRhq9KSiRZQu7qfFAao0yllJvlGQZUEQdrA4uv0/F
NsVJtd6rtQup15WRx8K/1JYa+GCqIhPuB18p+FMfY5/1gfgAiAfcHYvQbwQXn+Mq
cX2cuUvygk2QZgAY7U5IBMr8QdjJl9rVDPpfOsdKKceNpFzx6jQIRwQYe1Z4nwtC
7Im8d5WeiupKsv8YqaS8VdyNindtJlPwOeyKOv0BCWKA5NlZDqV3u0EIRPPbKzqY
7FGy6cBICVsRo/+aoAFIQbTk4pQRGg/jl1oYEFD2wBde3vHEEKce/a7r/NhnSXcJ
55vsDmyjEWT4wsPghhu9Tp03HHdVUdT60fMchIcfXc5yZFTeQpURaYji2oBsitX5
zqQ5BucACUJ0+D4o0XYcbNkOU69JIzkfAG92exek1q7xvWbYlctMci9Lb6OAv8W7
lqdtuZPIBHu5T1mtjtoKhJV6YgiBrZWEJfeUW7idyzb5oWDAAKTZfnxi0/8jXqv6
1VgEchi0/5V/5MIL+tVzlyVzs3LtP9UkSRgPIfc8NRqEjdm9zwT4hMAnhxKF8LQu
Yq5jg63RZs+AUhFxwh8vX8cKJ3f8N2KaaY8bA5TEMhMMUAje76Op54N9HYPWXb/T
F2n6bxLDA09MA8V2l2zdAdpLvxRFb/GBmgw5++5Q0YU1iMe4GIGqn89h5krDmRxl
ZohbRPhDDM5c1UNauU8jQ2ZQWKr+YQCPv+yLWhMQUDo0sBLmZd5nyn8OoWjmwsqb
ACF+fMjSIeONadUsgh1PGPIwgyLVUFcIN5SGiklOfKKpPYv300taEaJrYuutNgh+
0jwr8kJnrrg3NNKzM+5+HKFnPwPDKj1oSnZgIRRaPDgxvQLwgKyYEa8fmA180GiG
5wUovOqyEevlA/CFjrkipbtBxvfdS/BBCOsX+qNyygNsGaCjjqjfZDHjeWL9HIWQ
QGCY6odELb6RJfs0VJ86EhJY1Ci//RjSDvAbdE1E86kkps3aZDXlq5dRSVA/SwN2
4yslxM5lO7A790NNZCGjGBCN5hqMTDs/VzR6fh9+jHGe3IvDgI9bE9xweQftu6u2
e3Ce+cG1y1BeVa+93l91ZVTUIKyVpiX/oNRKdwlFL8tfGTTFrCmquHxCT0PqgVp1
oEwy21KsvIr85d6kq0ybBHO8BzBQs7xTrJRvIfrm6Qr15an3joPZ6iEVOKXq8b7H
l8fXNOLGyN2zNRj0hQjVvQh9sXH3OQ0ZtGHQN35vEfYtYJ2mlwN9gdnzDYfhNH9f
STnXDjXcBVTvMuAY+VJ38HDFPVKWjmPi+/PzyLqyM8s7/7h+PZkyJJW4QWVF2rj7
8so1BTh//j4vSGt8qEU0RyUuHrw6yr54f7Zgw2piAJD7GOvdcHiRifrt8tl9naUn
P7/JAJT//cgqRJf0DLvMz0Va3zFBgz3YxZrjyXd3/tYaQuvzzVylZqn+WFH2XHxb
NaLSQIKfSIVUv5oS6fkdMOleNr2JLwGI4gBJQjFcIU5ljUCXNz6sN2c91AHtjlYs
1Lr4SHZOFFqRse+QU/wVAQazlWAgK/l3TR3w3e+0o/bzKyiKQBUQ6F1EAxNIwjFK
Mvkf+u4I58tzJqbrtJeVhYT4FjjK5P94HeOLIqET0MLjemJK7jmW7zSspeCZpFME
dubO8znwrxYew9zRWZ97278Br52KQFQuhO5y2zlDtJZyVlkbnHvuPJr4zW8vM1Dy
9V8COd4emuV2lCFlpWwBfg9Qt0uNechVjBwCkWA48DppkDTJY+f1LrIMN91rQ39l
dlqtLf0+ilAHNLU8sB0i2P9jKJGlV4RTjatd7iIZ5lHTWC9NjpfE86kYCOJSfbC1
XUsRKfcERD9PVaq5MoKQ86DWz+4pZPP1LqH9g067LaJ+KUVlRXaYG7ECENhYQMBp
I/pv0n6E7gUxq+cIhJ5mUW6rp0MI5VU2ew/Ps1pIeIP01ykcScyW47bpDOUBmdHH
NcyLePIeB7ZX7KTJpkuPlwNTrqAKTJ+MQrs/8+ndOWp40VlgFFEygNADmb54Ubdv
brHYHTj3kmkikqTYrlfPTnxqB7FqPiCV1mjElR80JQh2b/0n3uc929FehgF1AWav
SRpehQ2omo3X0Z0oUoZjshDxzDhOXlzUPVkmTC/Hos0O+P2gh1esztnBUA3A/5c0
nN1kE4P1b5IWxCxY69Nu/PYAk4CvOXE0y+V592o2Ldtt3XKIf4OyvoKHFMBg6Zch
QVwofGAg4WZs3ValzGe+tjkoeXBIPn4q/wORZx1wOHUzPwZabcxAkuFbbA/yF/eF
nj+Jlz7W6tfsJzOtICTb+yZ50aChtJ/hVzYn/tcB7/Ce573tjbcQ5acrq3wFK+H1
Wl9LE7Ruqk8xbFeUn0t6f3nEqiZIBNxhXUH7zlzkikQSPcKsr5j2mP63UVQQoUsI
yLLrGBg8Zdcbcisxf+9yaaF96zjqWsLx2sN4gKBRXa65SqxWKMfvG7EZhm3iMVLX
bDS76m3eBJO8TGTxrGiZJukQlhuI2BtH/PDTDUageq/tCsA2HEa2HWzqZZ4iGDAU
PPcHOrdOosjWT083ucVWvrLKq/no/DKDTNt2p8qBh6UEtAFPiLqVvcuJ8VSIw4Su
C11rQc4WbE5cmNxI2KQXZLwfcvOMACwX3zK0FnQYJjVeQb7e8D3NCT48FZyCGFLt
ctCNAu9i5ISswrV5FsQFRHy9kRghngR6JyQKSZNmnAFDrLThAxsG6kf1PGW4Rlbl
239vRUgFgV/+WoKjxe3M0sqb52gAiX1bqM1puUAqVnNGvG8brKb8HuCh1cJtUNZl
QOXlsrDuX+P1SCiG4vzRWdtEwn8dt+z606crgZgtyQZkRDLKzJbWSZhJQDjgm2xy
xA5FnB/E6nV2P5J8E4KJN1fCaY4UAAr+L9MVygTqLWIbBaxVGjm5zGRpRCxpaKJo
gfJqQQbXwwMKgY4y6KQQqDo+ykGzCyjRpblR6vPxTqNM0T3h4vQ/NkYBSzObwtEP
GSPpF5wt4akp2Bd3AYl2ZmGKgtXXZ5j4DbHKDmL8DOEVQSL0jaVuMgFKwJaa/J3d
QXRDzVim317pxJ047PtZdTWYxnuzbRsbwxksOK9rEZMVoMihGpQZZXmoOiPl3Y4l
8+dSIjRo4YBbl5XgT0h4ek31FLHohcgnPm76HWXmkSwGCCn8ROrf/L/1OYTDnevR
t4mx/Q8aR2k+jgd5z5LOrP7D7RXrSYktOQ2c54CwD3FwQMFrd364nRAprrMGOJsP
flGlsB7T1ttrz6LcLaSrXKr3q23AVWNPC8bQQRsIszNj6CI6g4eANrqjKEc3Moej
unj0Hr6aNnZvw0A6zTGKoLpesIzF0JwoCqVhYpS2JAdWrDzD1d7TxI71UWNAFz8b
53ljbvR66v2E1TwunkYWudWiyfXmgyUDIn710mJ3H2Ty/j88uQNI+ZW+tR/n/Bhy
v3Jqx/PjHDCbBdDPmf3n78ZSFiwtuS4yD7S/PhK3L0tv6RUJqmCWTJVrKIFXydEI
8MtMicIZIPRJM1YBmqpaXxRC5qlPk4cd/V0RbjHkkcsEj0LYi9IXSC2T8eKaiKUT
bmEgnzuQm138LvIWIJv/cIEuOnqKM15LKIybr+9MOo8VdfPW/vgRWyK7is1/xwe2
2KEjAftd2Q2z8uk+0FsJ+Bwl3kWFuym4dbjCegPfdFkaI6oYA8P6yHL64z4EGiVo
ltZ7xdyMacGZQHcwaiMpgySCmv4oEGlGeBkKH3WRaIh6+GV3QzewrC9S3eKZ1SZb
p4NtzTkOsgEJ0pa6W3T/nsaN7q0iCubOIk6SxaDCgfvgD/LbXEWAYSLpFOaaO7OM
H1/v/xO65/0XYjc7pO5ITouhUCtJ/LE9GhV3siAYRMK03GR9SRBBVnCfPSdqcdiu
y6uP8EnrRVWo8dt7cSXRsOItEYgTjoDa+oFaIPRqroBu6Y6MDDgVL1qVi11VPvXO
DUIp8NzM7itYK7cLc0f5EI1GO06rjp6pznSi6YF6AzKlCS8NViAkKTmm/dxDgn60
BnTBiUp06hCNZQ5l50FQRX2d908Rr/o8r/aXciLPoeHWTPYfSKV2UOq3KEvjQnz/
SI4N6vRLTLWdPBqFu5p6ljNdamEvcJdGgn3rgr4LC0EEx2eMiPslT6LMWp0pJHQ6
D3zoDOuuDdUmpO+fDKG6MpDaknq31eavkaoY/g5hU0SiX3wfdlLrm6XNEJtcmXZb
C1O6VkLYgszEVd7mA5qXucciJepqr5HhNfE8PIrA961pAJlRjtP5waXN2uxwVNYW
boTl/evBA4vEQD2Uv9LWzdhcuRS4gorCegT+72vcpZ2Qgqt4nbBxZQ5JeWH7AZkI
2vWh/wkCvdlonwjYmPA5UksgNPmOMpxveRaqSzJD9+cffXsetU4oq2yspoowmxuT
Cmfj/hN2qkJ87/KcozoDlQ2slk3UHii7nl4eX8/ujWLZ1eUF6skP0iiMH1Mz4PlK
EOnUA2EzHnqs/VOK0lRmjwC4SeFWO3Zfuh7EbgJLTjTqkMoVxZbQ2XIQT6CFIjDj
+R62dEnPOBuZBFiwnZS75uM01l8WLtdQJXBhH1xizS1dOjZY7lQTiypZkn/TybE3
6mPQxLOst6ZYIBJF7RI68oYRnppHSHKgba5FQynwD6JxzoiLIK+uXMr1DW49M6FW
Lyti0Z2ZfDy6ozdf1Ngk8ujLa1v0k4PAtsQ47M43y1IM9x05DgdtUjFsOe4lJOgn
2u9eneU1Io1AsKQTLJfJEMHBKJAPofH41qT/z9xBXrqCT+1t14Ptm3azE37U310h
DKcQ4dI/C7Wh5MmZoNW/zucIJ9tx4wes1dp2WLgPGFbhThxNBQZVYLQhSHigX65D
lBIGkC0z2jVsWcs+8q3YF1JrNQSYwVjI+bZpGWTG7iFbOB202Rmp4SiHPoKdtF1W
z32Jf/cFWL2RXfdPMuqky2NTe+H6fBNOHtQMxBNnBOziz0FWTcf+FrWhGTJMae7A
Sa9k5DnDYylpTGiQuxkqXQwK057WbCeXOTKMvTwhwCnwONjRNuy/1zzuyfNk5LuD
BATAn1mCiMZMHvzPdDPc5y1GHAXLVgb4E2446jzYsr5FnvBWg1RE4x1dE90vntba
sLGIbGGGU3yqHaSuJkUqw3ZgLBDry/V9LaruAjc0auCdmWn0qUzRIXHaIJLGej1b
GidabeISgOolLRiFQ7OMz7K566u5+ijn570MoNHNiIqhBHg/2UelVW45/VXmRv/U
MYWdDCmrtO8TFa6W8Y7bTbmWsZiPY4Sh9+KmbGLyqjRwHTknAuZzv0PXM2IoiDXW
9KVq/8vRpGfof1HB7mA+VtFmSKas9up1dljyWQm5BqByaykmiu1PaqRZu2bLDdlj
TD6msyH/AeEeFiKp20Nr9CtVDBLVoCIKFV1ApOcPr2dWvlS8vl2m+rV/7SeDqAlt
gugxM77PGj3Ex+uCW+zdTX2LIdMQadr1cVI9KryhQG9iYtAvkkGfGNUlKxxcoW/E
CybWw9r77WMtUBMpsU8FcNNf0HnC8KK9iq2plZFG7vX73FX3zB8n7mx46bof1f0q
osCKOvH3lKCWszNSQlXHC3Iq19Jn2dSNkRBb6GOcakL3xfFP9IAEmOGZxNYVEtOX
OSJb1Heigi8JbEyB3SR7uG9jAU4fAXky/RAJKQovNIMWqBSWqWX3yu3bo0yKeC5j
96xQ+OaByU4encRCoV1Wev1mU5b8lIID7Orhz69erLmnN3UGIeGIS5EPDiSy/3/3
A+5poE0lHiLaDIwNNqV5BNLOy2K+U6HGcUfmAjidTPFF89xA1UjIFZnsIe57fEcC
nRXZvY7EMBqY8gkL05xPuOVPkOL1+66vJ4MHmQYV0Xi6OONr0n5aF0kmI1OBNKfh
54Qv7IYHpEUkxbgBBlZkdvus7jd0OTZaP13swsnwNAhLeN6qA9I9Rx3Os6+wa7uo
tijU9XKaZNpLxDRuDQSMflFSel3cj/tn/6WW4petRSxEnTtg6l0+mg3cm0FvSb84
unuBWsWsx+hrZuBcBi60i8MTbZXYlD2nmS2q97inYZ8JCs+3u8qw3EsNeTu2afVt
JOo0dCSo7ytcMw5GSuOaE00pP4lCAe0diOJT6GTiBHAtUI5nnu8D63STod4P9muo
nZEi2m8ySwjzOdQhN1M7cmMHn7ACETy0jJCF0+i5K5mr/nLfgZQWMa+zuFiPSk8I
IVoyit3VphY9WKF9ZDHRM92MzKbLgWCZMSizi+41oVurp9Y6Jhr5QIfE43BvD9Iv
uqd0VbTyINWcVN+L7qkuM6+Xf009vR6/bUMCu7ZfVPEPSqSagRkmQBOaKm1Fzocq
iMddXOKnC6AweZHbexHDyhmpzeBKaUED91vzy73NrHsLlojNLiH9hxdWk/dbbEZI
5HPei699xzDkX83VGz9yGXNZp2a0kW8uE60Kg6fzFSXjnUvvxwNXUGjlNhRGa99i
Zwmuk81KynSPRYQM632xQbxZFLdK8SIYVDecwFKw+3fRWqkCo7dOFQyuyDHEMQ3x
LEHoBfbWQryXXz39q0mwryBOrmBxGC4uFe2pw411BSPrM6+w6UFTOd8hfZtgmiEW
67hJ49FAkFXOVz1Qvfv4cF8Rf9Xh7kw7QQZmtGxsh7TBUFgahlnDKXqY/bXubnpt
W12USzcYrrNNQfZW3noUbPvO8Pm4B7di3dHY8ubnU7+vzHsnFUhKrYqFxgsriM8C
HbQZdui8xpIYM3rFGfmlveQw3Z36PCJlXz77dJQr/re2h2HvrAx+4R1iAtsYSxQc
7nXauKSA90mcqDy7WX4KEYBQtLv60IhdQ+8gAIBQTRZu7PWKm2Y4GsPD38dukE3w
5BuGszLuVcoHT9slPwhZwQvzL5TMLugzYyezWRV7ru/BAGG0sXHEsDGzTFv09+UZ
Q/7wZATQxR0QSSlv49FlRg9xCvUGyuv9Op1qJ81SLR+P/FBhMD1eSuCPDPP6F9YK
2kfy/KOFq5HYetzthNL4sRbLo9pDMibJMqP8vVdL34uIIIGImpwsW2OYql0f/VHK
mZtVJSR3C/n3yBgUQBrFAvzK/E9SGWBdPBuJbcg7ZvdIwzy3zS7/dR+N2Y0ccOjM
q6WWwwt9c/Oz64UlNCC8z+l/eS6+Ryni3Cj+h2SHvSpHaMtzDJDJbB1VMPBsMhJy
ro061LS7XgIdIhutDOM6oasdHEsJ34aPr9mpq15Jju47zVHNQzC5wOKmHek/sRUE
qhIqsT9uoITjivXEm0Ey+v8y9MIiwSZ/a2biZlt2o8BChCHOc8q1zH8EPyWIa8LL
ICv2fiKDwcDdhyb3e2oPgKNqxmDlidbg9sge/kAo/ARZ2DYQBPJypwb9MhbZ81t4
xL6sI8Z/mbr/BQ/LhjeA76pkfNzREJz1QAJvmN5A0GrEDz6pPPtdVxwe+r343/r6
+v6cMtoRTWOTzj7HjCX5thMxyS3FMepMdWdKFuFjATW4QRXg9PImrOOEIUnA+VQO
tQMp7mRJH0AsXMLMuBX2555cRynUgzLgv2l5fAWlrygwfUvqhO049mb9FX7eYhOW
0URno44BNZNEz1allyD42g9X1CmMBEFtAdsef+kTEn+HljElSa9GXjOx+PKHcRkQ
uBCbEFf+cBIdyiIwcHhRmF29flR5ecZ2BiL0kjP0/RstHz9Yg9jGQB7Os1OKlIOh
Nhsez7E+Wgnoqp7oalynhdkKiH4nPnwIdeK18W8ddB+4Ehmhl/dHtOWUj6R/VU1a
MvLfqVwRuFc8ucitqqoz5Doa9g/Rs9Hs8ACVkwQKt2wxU1sd/8DTFJ+58ga77bGO
70US9nz5ImeDj75lBfHekTvZofsF8aG0XBJ31Iyd39Red6nPK8jaK5zXgZulNFUq
srM9TFVinGxs9QH4BZXx1F4xK7mdnZxnx+Fy8lkhVsH3X0yxI97xDG45vqrgVSOx
RIHNq4Zu3fVgBcn3PaHa7R2E5o3h+SlCXcYEniBaAINNp6XN9iQU/2mlKk2h0/Kn
clOCsEgdDjkzBlT8xC2ZV2Gh2AbZYiEaUy6ikWYo2Esg64+SVktRU/rKPwPrXLPe
vqubHf3Nz3xlHOvOyupmq7eJtnPCSvJ0+MDU7cJn6qB7euYyzNytoMUR49ppPy3A
GBP3ODbb0Mdrmet4/9k6x0sU8fVbELUcwb8+/pyMGiO7w0RJkoVG5FEk9NQM0HMV
VOPu+JkhEKTzWn8Q3vxqKxqKp0jH4x98InzMc7D5ONHfr7biI4A4D31DRoBhao/V
+aFUJpNb8AdspXVNStNt5tGDbDl7sDpgNWD3ERkf8wcX9QuON7tQMzdXR09LmhLW
sK8WePjqpxq0adG1EiOOaT25PQlmJNOF+Z9pxSTaZAfyf25eFNtxv/TWvGS7jDlj
ZsudzL4VsLnuxKrz0ot2DMru7gWJ+f80uD3YDX35Y2sNMID5PNsf1NwWIcpeWmlr
kLQ99+I5h8HhE0P5zU/+W90IaXHxnbFE1M1J7lGL9O8l9rXFPwkaJEFNU7JcLI1u
9gpVkKSdbnWqL7+hiTr+xqbcpzAdF+/myh4Yq9LP5T0WzxnmR2zfDdyhiwr12//P
ZRCXuA8l8E4Fkptlw5DPbwErwDpXWKJMfA24GbC9+jgTRDAueREPx/lqPpQJXUhP
1kinc9sFjTHJOndKiBc7muqWq6gag9S6ESeZQCV6q3OPhNLaieqB1B1SuLw4Y4Wa
UucKR6ADVWqii2fvY0uvL22Tg2qhQsbq3Rtc3tE4QATGt8rkWSOwe9H2DMZLatMA
Ar6TYMHzXqGWZnhhtlMDoSSmroLWvm3jFFAXDjbAKYpeCj6kwC+if1vOeY7jNxCa
sJy1z4nHVrB1Q1jRX/Qs+g66uspt+ZR2yFisOQseIVKfTfDvLV/flunG8R1d3gIS
bXAZKV3hhSch3d0dGPN4FAn/h4JOUZar3fC9yUiQ2apnnHh4H/m+prmkFbXGvpx1
qd8g/Abdc6+wtI7Kj6BU27Z0uiKG5Nv6SGZLmT+pdgnL+XnSxk5wk67cyJwYmhJG
YOLTTUYUyWNJDET2yVJqRNACWfIcLI5MevQzB/M3uOtZquwCpjhmvEeZBtj0/pyr
0iVUKyrbTktxFhPBDyR0irCon47D1T/06XWrmHJWIrqSkaX/xZ327XJOoOFZUKgC
zsJFMSTaIS79jVjnEWMFBrfB0u5pXYSwYoEy+mTv2Da3FdYYSHDhFv8XeptCTuRB
bw8ONDyBaJAfdRwpjCcQzddO7MQWtkC9sMN08HDSQpcvPwoEMM0bZcgq8FPaYLGF
BP5AQqxa5ge37Aal8w6wZ66lezV+/0EvglV1ibpCWOndFe6BRgdEpfFYXF8NaqXz
c+87cbq+qwPWHfKQvpmwDI3l2oJb4OMgSnYtnx8gRXp7EaLQHeaXKUXFELhLJrJA
+t18My1V9+x8u/MJ3uGqkgE3V3jkx1fgtvBHwQNA8R+NwDUxh3wSCax4fIwQxwYQ
aMLYnIZ+177ZaGAyHoQ8ORpd0tuLrGABq2Jt07xbAGtkZb0Wt1cbDTMnAUFzwHmx
9GMDHAygE4ib1HtxKLd/BgiZYn8O7Qmx5BQ9hX9IBf1K4f+lDuqBZ8Vlys9XhOyc
vf0XHkWp+dCa9KNnS3KEuX3rxtdmg8jHEcYw7hKXxNBukmVGaHvIUXbynZiZpNxX
0UNxRJ03/+iYzsMxm79kURJ+Irc7TYOQlJ5PNRv72gbdQco6m83NytbNGIITQnBZ
UKQ/mI1JdrbuTYNtmWLGeCgut5yVnB0EDF0DmKO/nE8eTyPsrm4Q6+bsnTSL95hJ
vVQerd5WSU8oh2/PDhMOXy8EKItJANJIaQ9MLIQTWImMGy+lu8IjmrsXaEI5jpT5
7zx1cq8YfDi0u66IP53jx3p+Wd7R5zZHs9tL0EtBGIUvZuvife8MJOrQlF43ZoS0
ptLfIQyopCEV7f2/JXJYj09Fq7sw0h5J8R52FHTOLEBmQ4TIsk9d38uaNCzuLbWD
lgV8A+Sw9ilHvI90VnEZbqK10jKF2AkaJUxpiPfs+NzNaJnH6kMEmaV62IU6TpEz
nrn31xpaOuMGe5FjQhPY86OOxfdW6RPJqdZwESNbXOW7viuqIkS57RhFVaOOjcv4
wQ9wVntbR5pXQ8FJrRA6LUL42/J16fpVHjNggyUvWrraAUja7tIp5szjOKM3yOA9
aEp4yfsej80fXC1eXK9vEv7BfVcuSVIMToAYuZ5Z9dmhPclirSVXyzW6rnLwJloF
ylvQmUunZR4JJlAo6iZCH6XjtNLqy9mc3YplW5abvAlK+NfrZyEdkfa7IEcE8iIJ
ye+HvSddyKDScuik1Ml7xI9ENx1mI/Ipx9mw3zgBiIgdRQIeXJhsppEEnS0EHMph
OqdRpiGQL2Y2W9A3421/qp8u4LQaGWP8dH3s5Oox8KNyna6h/42kjHiiaiR5u65V
qSzaHqvYnj+pLqOXNyOojZGK2wwTjhcfCnW7npC3InW6x60v2UQ/Xdz5PqcyLiVK
uB+EEAYFbLMMgU8JsZEWRLq9r1cm1M/m9PhbKhXzt+e9XOuINeSzDjs7tvBgrtP/
xwNHde1V3B05Gv+dQcrsUB/NW+y0cajqdWqoq6gZEXCLZgGExAA9x+JPTuPySdFF
sBzuuhaM628GsZk0A3g/obnSQmPB3kz2HtALBeVn133mwHVFxYrAjqTfRWsTHIIn
MLG+k/ZtZKzLL0dtzccKKWTjaRHCQxCmjLTkq37o+3ufEBmNeq0EiHVvQ4/3wxo4
IUdgKyaCaW2e7ip7JYnMIDgvtbc8oArPtPuytXeQpTZZTYSARyzVxm0zcaJ0GBDe
66nObAPIjZmW8W2Mu1hDuepwWzYkS8gea2p9pRsCSx7EwDn3dYcjaQ804p4otcJP
tcOdAhS0QEXLOSQpr3OhNwg4xzm9wj7cSRq7zcKIk4aTyU5ldYTZo3TQjWxtjin0
zAuioZorZu4VNlDGCEaWl9d8r0U2eZHRen4Oqyl971RWQRCZsNiEoOKgkVk6gYKE
H2JAKRi0kRDU/8QnmeL90i82fMggD5sDCBAy/cMQ7cIimfeAeqhCUFgjLIlZTi6J
pCHmi9m1xCNq/nFNq1kwbNCFQs4aP1Y2hr+bGMSRnGdChuZrDJ369/XAIW57ONbD
kBXmglQ7Om4cTw/ndBvFjZuPlumu7COszwAN1Ib4u9x6U1rPbQiB6okQUnnHtRsg
RKYWrWtmQZH9Y+Lq3KHGZaBGgfW3Hygu1mpkyOHoSlM8Ri20elSOtE2Z/bUrcmNs
0b0cF23B1L1AKDkk2Xg4L4wPA1WXh10P7gpk486SW9HpDvPpjnJwf87D5jEdCX9v
wDNCRLtiEWC92vNnVq2ls+3baONxlUKNrc+/D3Ju0Z2t1JhwvfmhP3GT02Mcac/w
CqmkI4RTlMo+i2CgAbzEFSKZG/GPYNcy6DqzcBkUb8tzbZpmn9BhDHc9vwIT9d+B
39r3pdAw9t/I540HCx0waRJCnwt34VEmCTaU+id5eQ7DM21mcW5/DaWUdF0Y6B+x
26secp161MViIOss7KV2g7ZKgMmTU7JLo6+KJ92TbU2IsY/Zvwvh7VkJ/pKQgDyC
veFprIMspPwRDI5ipqRqdX/9k2LF58fkOB7ojUD6hK7DNvmgyc3tslntaTM7cYXg
dmWxCwAvUcIJ4gXU8iCZWFFQiWZB3JQ/m2YPVu9hCGTq6IMM/yj/rrUxu8at5i6W
2Ju1OLwyE/rrU9koJ0OcEIxj/Rd0oiDHeqoM1r3qT1snRet904ZxRNkJoVCuXbwA
1430vMlS3VzKLAlcC1hwHK3nVdc1B3d/A6pUM8vYio35wKhI5DmQId3+vUcd3xq6
l4wH9gZC6oVQ/nUfR12PHqWL8sjpACgokZbKKfFXsRDCZEBXswmapEHsmVyZunLp
ut3GGVtfT39/eP4ea6kQosUMdi7p7PIGPw28Dg1xiGzJXRjOCk/kOKSEPfSFyvXY
YX8AV8djymM6gB/csCQFJKihB3zaOQi4Ik2wsdvrwUM2xLUcCptIQ7Zk0yqExCw+
9t9b6hIKjSQ/E68Zbs/WtQMcb6A6IemYGsJy2JOnXRhiTX7zfPYn++Vy7jPbtsbM
T8hRXtrW0C5r65Hxpg9XWudmcZxOCLF3NDmQM6z9gaIoYv/gNMAJA097sd28QtNP
QllDKi6IbIHsEuAOCJ9axwNzySHGJ9tx2ENCIC8wzCT+V+3dMDqL4SXR17t+5+Ih
2bMN3lIdOzutHVWq2qp63MWGOMwDshCpWLuphM1zYULSzyigMUDkMIWPvNXcL68b
iop9UYu4vAXJuQz+8Cf3dSGVhHfdw6hljyq4Q7YsGKa/fSpurceq+hvahVn4xZaW
UQizN9/LO4SnZqXj88dmRzRw6y/Bw6R1qehXjKWaJc3/0n9jHe1aCEpFqyFuInyK
jFBz/xrvEvsY4jXyySqrW/DKsShKrk1n+zUuIN3xrSlwN+YwP4yZyvRvZo7J5kdn
sN/4lHfrTy3GVFHu6Hc9qQlpI7X0HQf61/8tcoLN+jbXeXxba+OaChQjz01hso5+
V2FIwlOLn+xHSjAHbpWDo4V6F/esjaO/QoHl8Ou6QJsx9DcPFNfubdthLUtdJP2m
41b3QJphdQHGsQHg3y2xdEZR1rHgWJgYoXTUURMT/Ahv4ojr2LGLcNCvoLfBdQ8a
OKD7VrlAk3IehBSZWsNq+oRy0NYZJ6E4+/cMKk1kUK7YbLk9k+f+X4d9YK4SS9Bu
G4T7diHdZmPGOnh6xkWCnEK84z14KKMFEC1ahCoYSfIflidpZkSRqIeGNjat7rZd
S0FSLF0l5tiu0Tte8F8Yhe/ANmKNlzVVhFHWyhJN5DJ/WZBROxLf5PhgcL4GPwUn
TnPTNxCFVV1cFjzcMkzKUfgNj/2fOyg05Gfm02yhw8Sr7egbx/dniAYkOQyKusPC
KqI/C7U213EfRsnalgwP/npXMqKaqIEhkx7OyLXhF6aFzD7dORIyuMZrm0Y7iktr
YHWOGSHRHx3YbITkMt+BRgBfHYaFYTv9nKvJkdEpGFFh7zPYoYmRRDbO8cgQHIUR
G3bEiLEI+aSmb8ciyYHQf2PyHwMMKLe+bFsPFOet+TzO0FLEPzI6TZA7iQL5kGro
8xVxox3VhGsFa0FGlvepzl0lvYjg1STk1aF8wTnqJjssjnZf0Q451tntWGzSpSYf
LYGokHcRfBM9j8Wa7+OC+vIL/hT8KnFXpkojVshqRM9Uaa9EM/uvlLuRl5el+k4M
fYu8DPpgzlQIkXZbtnukzHrddlsm0PJYaxL9NWPOOZawwGgtUgRpqGX48hDdUozF
b2HUDRFnwVnaFq9mqFbIbeuUf0TFU2HOa705l94M5yFhnNjIfYidsdAwZFhe+phf
6Pil7jR235HR1ctqryC9vTubwj/FJqIaEC3Ty5XeRLjMDQnuaPmtuFpHoDR7JyaA
78qnZeO9YmyMNht6EFaJ/OMvByevoPqwT1t25d99t18Nr/iKsh2nTetxiTNwrKTr
KEKrZLAt9ROKLtbtdmQVaikSqgmCLHYLO4rGYi0JwofHJYUDhsGSmGiT6rt1pAsH
wn/4zuk4gcRAi1nax61LXuJlcUi1/PDRtChv+qtUGjoHZMw+OSH12FbRodV6NazJ
vwc89HLQQ3nNN1jbWDdVE6YQxrNHK+ogTJP0IwyVM1AyIILKD98v7LGYwxTWP6eD
/jQCQdr080Ivgiw/5wx+DbbqBSy8Ry+f6tFZ2vfNDdIF7QP25c4XXL1lvTQ2FjHW
7Vq9o0yFdOolmlzoiV5r+UNrL2DPJy13Zrg6XE0vAl1sDpUksBXkozhS0hsr3izu
JdkpS7bj6jXHxV9xb/WvvQ7qe+j4/nb6PF2Id7vPihzNbkvOfBU1SOYUww1Jyl6C
Uir3XirTwPfDsVExGAB5TGuevH3ZhXy3Aa3CuJG6TsQoptpcfaZRb7+XmjxBjaZv
vPwyNUCUMnUApl61po83fwN1LUbM3osBvW6ag2P3IcTXuJU5hETajvafV67bXsMs
kt1UAZ+op/Yeuq4alUx+3pfLavXaB4Cl+i5e0fHvy/hZ7tP1HbP1jWKN/ZJK+fW+
qFkWMc5GpkuRl8Wtw8JOWcb+Pvzh5dwGtX7BLS3SYDqypRDEhg8Y9rCSfE0oGGhg
4S/Z+R/ybWBd8HYZROeqbPRRjJDWAiw3UWUBony2f46nHZAeV2qjASwW/zD4smnR
Ddek/0/B0StYlfIKYg+DwUOo67WqBBLCdJfRrYIRALb5RolkTHBdeGEj+EfuUGro
TuEyK9npfxw/9XbLBNTfDJRTzZ8/9GTZ29ChQCaQbk5S3ERYLQUfmzUH23qGXmtB
+iWFozg43spGJ8Uf3ML3ZncRPDgQbPzG13ZdRGu/92Sh+r5R2MjCkWjYd4NMTxcj
wstckb0BYpi4qKGvlCs27wtLLV12tB5Q8KIreEr8aXphXI5PNeKrcSGvVTThadVz
4PUry+SpRcM7E6l0XHurdFfXHfqXdiBFPoyrqyVbpTS1sUZ186BLNzI4zJj0fvCr
9pab88luCO7sRkFMSym8QG612PZgeuW3MyjXSDDv0T1HH6iSloyxxA90t5HcFUx1
OJ7I9+Mwr7VGWERlWEt6cW64C1ZCQubsnfRxLXmPBXcKl5uQuj95JzQwwg+ZjuuC
E/z3lONWC6s19QPGyTiNU0jiq5Vcj4Dr8YefhRX9jpNdhmqLUpvZdSf8IqMRKmg+
lyMbVLnImnG065FC7Ig07/tGrj8dxYtO2Vzkw09xUCS/KTgwYhcyrtGe277qNWt0
MBJJOCCL1AHM0bDtWpDlh1jOZ8S+JaIh9dZvI22hDTKg+roqRpMzFZoxDehr6s67
3yQ4oavvP19yhH+rurFuFQB1qVjnTSYyR7NvCuIkjnHztV+j6XFobC+Mdr+yYGLe
2NOH+M+K6TMBIWkbyWp2a+srT2MXAaeRWYT4b+ngxrLtIvC+4trz2I9ANHPyrVPH
F7IDfzBkA7EZi5IFV9CurzOV9yZWhA8QgojLmsQEC1ljcyx2SmA3A4v1+uLd/FeY
km2hRJ7SnNMmCBPy6rUbVtiye5d9D4Osz0tx6vGo5OjwnXZ8ARQj6Y/15i86HIZI
hwie1w8Bg1VzakprSRJQRIxxvp8HuO4frEte7ONCYKWu2HbAxUJ7L97ZeU6lEOQG
MfDgONcADdkB6IJBWJkHXQkYUBst2pJip07IkCzDXCtK9zM5xA+qiMYfJWjPC3aV
4U6niCLcVvmOi/1O7KG1JD5jB0BmJzZF3Z0YCjxCzzTAWZO+JPKMABk+8yjj1YTl
NUTuBHubgQ5oZhnIU7rMHbYmI+6X98w+dV8smQQhe/2jIyVq/7e+D/+TJ9ybphUo
LGHDXlPlwnr54FcT0EFVYpF0HB8W6SSW4UZRGab9MGMXLyELW+35tlmPZi8QnqYr
5nvERMeyekypsPv2hz7+WpgkTb2MGUhdF3GSopTOL1jyFG8UJA5qRceNzi23Uq4z
0z/mMkjJxxtUOeUjfapD4rh27E3630D6VXD+mDVc/ni1kUNs15Exc7/Pj+n+O2KZ
nif7oeSNV50Sf8XX61gkc1jFZsS0HJ8pXXrnsFFCoCNOXEONZWJE3WMBAtLRk6TP
57yUlfzLQ1vwvuKyJJO0QXIjR0ozW/Joy6WsmsOoS6chwQvUEBxLOicjTEKHS84r
V1e6R7Xl2/WAqM/6+t6nhne6v92MSV6xS3lz5hO7hC+xYWIyeVirax/QDGXJnVL0
LIM8RzkuYjJbK9p0/ZaW4RbiNKIp53TavIL66Ojwmi3WNP8Ik0fLrZVDrz2L0Rvg
kceKfJfgeNJzASkyCsmhrLe1c56Q870OihordYs6HZhbPewh+A+nSVP/tITSLZ2i
eFTSq1sjTZOh3zQuoNHAcnOfL3oxc0cGlrxn7/9UHYa10Q4XNBlXb33APevXoN1h
Cm6KWsHawHW/a5oGNuJhKOwdH5gQDHOoheXp3ychnHUTT/WYPeA21q6h9GIYiUP0
lk9CaB4Rnr7DxJpRw8/hOPoVRLrVfjOmiKvL0bMWlgiJanTOZtr7LMqqolUFncDS
J3hhS64zMzI381jrC4R6GmnQ2LDxCL3GFIG195HYOAblY2I7ZKlA1v4e452+SeAc
BeeDhdp49Eb4zAHmHQ+NGKXBobYNDNigc58+wKMQ8cn7ZTDzoo/TuJ3Hba1M91Lu
GkOaUpq4g7gBibb2GrWiMO0mg/u7YaofTDAmz1/rLgOKezuL6t2o0dNJcTYdJkiC
2mrn7nj+GF8yQCqNCVN3zFR19nI1sBgvjHL3w18xoJUksYZFt4Yz8R8E0pvb9PKV
EtcG4lgqZQjiPrSjaIyRYdB2/RV4WN96ynkv12fs9NMPdWVbclNDDIy5vDs3cItF
CxxL8nRjMlg/WrzrgOL+utpOdXPRKso4padmIRY3/hO1fvOtKt/+4r99jZU3okP6
MUeRPwNq3nrzzDEphl4C0g8gMdQ7SzrcfRcLjoO71CRoqCjIZXX58CeBifMfcErl
ZjKBMtO7RPPk8FMuUHrxjyYUbICfi43ZBzSo9hAlxvKp5271eLeB/BTdT1qcPWjF
+Hk0pstMDG/jVUKkiNluEyBh7WWAdI4l4XVse7qhmw8sDaiJ+ULu+wjWz1jVVRb8
7nLPaROWCtw/V17GuNxuZ0sPuXpPRcmASGPkDzmrHYGYtDSMSF+hq8na5+EroPqw
TJpGeJZ7govjLfMeaLvInAGhhQtvLB2povHHko7m3ROww9aUkh7+n8C+ouJqFebH
U8joRd6Ng/5CWF3gX35u/nefy18OEjxCEpgVpcvPbAFzlfatPMElW3puRHHlZ+SR
NtRcZSnsTRfal44BKa5Oxxw/0n23Y9VXtgfWbFYV3/oXAIc6FL5wzDarmZQCAlZ0
W8F1g/Vn6idQpV7TvaYoDYQwO3AIN9QUQbqkZoSVMtCkOGBf/2tsva36AH5FzOIX
JA6zgR9dT6ICLP9n45eTlSE2Gu6EFDLRsbju/r7PD4qdKoOXwMbePZws2jNsBcDF
mqxY+bXz6Q9jB/RvrmxLnVcrDV2F4d4jDZzDIk5w8ZieWGMX6pZUE1OhGDrd7R00
eBA60tgueHzHN4W1oibVysw6z6Fo2NHiuamxAvtKLKH4U7Y4HM41Rk2KgtA0fMU8
lmp3A5iv9SLaIgyGDSausvjr8cPDYEVcOQWBUUp9yURWLM7noJ7BtBgx5mXi4LmD
bqW7hoooSzvo/DmuCoEgD6bCSTBC7GgYy2kZUtq+9gBS0jPTloe3YSo/6S5iWne2
GqjMGH+llwvmBk20z60Ap/ocM9AOdMwcG9SCn5u+BLQsWIEDW7dCubwYdwaOthDH
ckOtWiXC2YrskP1YbD5uzLLqmmmDX+lXUQ7PlZqfwEQNrm+gVvwRfoCs2KSTjoQA
GUslIg/q0lMiQvLlDKk3ryWWYo9VI3ZZuMp8s0ajd9eCn/6mS4MqT+czPfCnV31s
mmsX0jyMDBsgAZ2JnPuCLfFw/XwpYDgxyMWisTNUZGfRv1prEuLxiLSiGGN5DUlX
59Q2OaXUD8L474ZoWcK6GfBbsDNeFFQrCuQsWe/hrtrJ8odJldceiQ5qGBmcLWrF
PjAhnomckoYMNT6eAJPFABLBiJLm9yL6/0s991iOP7s7JYdOO5aojxVCty7JMsAo
hBkUuO6Ep2ubwfJ0kWw7SJxH/pQQ9rT0OAbt89L5uCafzrlg6Nqs5JQWKrK1Kti3
JdjhVgTmD9gSTehIdQDg8CeFUPzkqNMCg+LRRD1EME3li++fwrXwiCNA1lFVMXDr
6pTgNiv+nZtsK1gUl4fG8zCeFa3KtHlJDL4PDcwHaL0Xxxf/7YY1yol9dwfkfXR3
i7lmf25pPSCyWMi71VS0Sqeux0xrP5uTqMj7DbbZ+Cd+uZ2Ngajg81MCl8mj42F8
HXUmmdAbWl4XXzpVoYQQMqJV/sLujR1fAoTeXByFzt/dpQ/r/W2P3Xp4cjSn+h/i
jHeJ5PhZLHyCCvebMj9ogBDbEHbo1UNGLD3hJk4iMt43hPRZt3wN5gEe4o9/wfqd
aV3EZrOh75RyWZ5R1AWUbfzkJnLQbx9p66ralVrEJRb0w8zHxDWFQpQ12VVwbH7Q
NHkTWonoTYk8stz6TMoy67i9r34JlXPG8g1t52d6d14hLkjyf8UOOP1vrP561f4y
tfWFj01adeIsqwjQ+Y70kxIfHJEozyUyqMEOOj14H2h6/lTO89Ym36XiE1bo35gf
VOGy823IZMTHXizCjEyvNOOBtTYBjBAcd6gBz+orW9CoYNcteITvCKn2vo8gwD2M
RDSy6+XQTlUzzFz7o2hSxPX0Tlj46Yx4CPZQjJ0a/vgCY2Z+vOBte+7CpSu1oFrC
KR/Lfo5QBDRfksRPy89k1U+uFncu0XCEpNdo/t+dJrAbeZq9ozK+nGDpj8Uec8lm
9c/2ab5BB7yJgWVyLGyHU5zX9v0kB7dYsF9ztkAtdjlHKvcZYpzNC9ULDuBPKrPo
wgbrMumy6laPLXxyZ4kenLXkybBR0xBpAn1sbvgaNgCNbuYvrPBrYW/nphRqhdlv
VUnBTz0Xm3VcZs+w4xX+hdHO25hRV8n2SwN4fmaxMShgpwK11/vdS9un/I0uY9gA
hDAhl+yyl4jSmTBmrf29vIUPIAZgan6MEWOnr/QT8OnX9olQ8OrOc6J95YRgZYh8
YPi2E11K44tSJVzmvHLWZUOKZscVyajuVuXTGWZUbxdMIadqYjeeEYidET0hswHR
S2Evx0jLPROatqOpafK5icFpypbu8do18TEAP/2aELhpURAdg826sTPU+MaL8b1t
RPh/MFuQIZjr945kCWwJPV6rL0tjrw4G4r4HSL62w7S54E9oPOOWsThBCvEDnoqX
dYqbyRAiEEzUrroUxqON1SVVn/HhSSgqKnk9iJP5TFKRdq4r+xDn4EoDL6CsH60X
mh5M5jD0rg8jcyzCykK5W23aB+TENakUUIMIWvO9qELoLOmxLFiEqgpd/Z1Q6Tjt
b7e+iCFiPrJGdJae/7rkwq5NdQFnI53OlMg8NHXUQiYolkMzGH91ov0B5RELeIRJ
Yq8VXDrMlCYxmvurgXdzf2e+IiMhAH3Wx/NTqlwDUMWqRqQNKpHiuPR7lshmtFDa
87CNLoXXteo+d4KEK0YJ1jr7KhM6lrvMAbxAsA950WM/mfmYkUMPGFDPGdci4AhM
Jh4qmR9KA3byFYS8u7GSey9tPLV4EVNBaQYrC3GifEFk31T5lRIPerf3wf3Z5xYi
8MmiXGQny+uZa7gfXZ7Rhx4VyVs+emEg0vzMhKhj9uFZ98l+PyqKMiiEU0KxlBMu
UZ2hkPEgkzbp7WaT0rkShJO3MiQLUB57HXSCE4PyV3uancO3+7avI1b8Bk+Wbsbc
HXVXIWsrXoTufQ7u8RD7npdYjTS/DmpTWH07602GzH4rYgYtdkC34+Oy4OT48mMr
tDoB2dgd5LA1uMlB3Ekm3g8c0CGWuPdH+NJFt/jtFQtsJyCL87HXrcPcDm2y70Qj
LS9F+KA72Ei7Zbu9U+qpaSXzir1Y2MGedI5gvhCinq30G7pnwBM0s0YLX4jGW7mD
i+itMct84tFpIEfBDEbkadYEhOafvPsB04AlhU5jaQPEowW1WfsqFpWfdMSUDvb6
iIQwMY3PHCd8cvEPXEA1urx5m07PcGgxDPZCRrm0KfXSYzkmamBTEqhkHhMdbGvk
P23knvl5wGh7Joqh61ClDgiRmTJPb7BuEBv6IqvMKIPaovSG/QIEPd0n/fPDgCls
dPI4zpBWdnR8Dc4wQNt3gJqCmXFSoKOuJblcA/tNs9nJ33jXyP3GN+n2y9Cm5xFO
E8cAhmrpyx4YrBqLE40ApRS5OnhBLBgspDhbtysiiDMOAJEezwm/FMhm0rfzClTn
Cb0ruifAEIh6qEiltKD3NeTwYKaa7/AwBHu4nIHZjQAsm1vp48gQhAoSuMBXJGwN
jVHsPTmd/AXCfMrVUgS9nOGk3IaC3vv/fuymtCd9ahhz/h2zCnZ144jCXzIn9YVd
cdgveWhOiIIyW89/UsLL632XgM21RtixKO79Y0jNE+fpBLdVlV6RIDmbJfbUqmE/
pw1tV/qm2Qqnq1EJLHKarppGd2pUrA3rIwpp84y3uM23vLokyG6vKT11Htn/nnmo
hMWlYn5jsc8LPEhayI6S5TR9p7HN6H2gndQ0sJsPSV0pYItbB0ehWdW4IE6WMds6
8OF3ysDK+db0+xBy4GIOtlbMZrpWOQR2UyaywnfR4HPBmjg4HbGxd5fON+hFpd2Y
iPnWFbXi0jrHYr3ovimkGJDLK8Uzfh+ZYwcCv2HmvrBmYHxHq50HAJMspOzLjIzI
fiswrAf3D6BYrg6THT0ImIujkRy1G4Wo5H+HFhKs0eW01LkhcfNJT9X4d7LdFsY4
MykolMxGSRcC/b5T50OV3wm3GqrLbrUuooleR2Bc8pdBNdpZjZ6NxA7ujb96pQCL
O3jT2yksmk3iv3X6QQfuGFSVdisgWIS4h8rYcV1Q3rvXivm97eXWvLKkA6enN9lq
T8QAKpfB8Fxj5YvD//qSO7N3AZOUHLFSIYIB/1TOTxtP1OXuh6z9jUgkSrO04Z0D
I5cXQKxOlRlbWZOs1WGUi+D4InKd5jxY9SQW89aPD86f1qv8cKBFm5Occf3RN39C
r9zkXyt4P4u1V0eqfU4lYTpBCcltooMvFydWyZKbIeLBE2v1BZBGHRQXKyiDdW9+
ZvGSRURpoV6hyMHiULQlnx3X2IdOgMFnll6IwrOEueJt09Tmvp6qla1s5ju3oer0
iA93avw/4gIdjG3b/Vvx3tOGJ/PxSHBZM4DigNPJFwBdn5KTfR75VxX8NL4gCdGs
1unnFpqA3Cs1CTh8cCw3mSF+Jenlw7x1aAQUzeOYNcaByG3rH9Ug/bQeqTymo88v
/dKn0x5PJkitqmAylVIoBqG3bCIcVfADnj4Sy/xvQoXocObeaR8tpYUJqhvZJ3QF
eu8qRSI5A0kmcR/SyfcTobskoeZ/PtdRlAPPjTyBz0gmD3cAwU3HxUqif7JJXbaK
V5ycMrDZ6V1IpVKjH5oDovR1mjl9HHwInB2WYQfg3J69py1EdfAE3F6SqDfzq7kX
mP5NIIP8vjf3bOFaM6PGLKh4HP22+nnvw497BlPheW5s281LWt9aX4hMuXkmKaN6
zaHgCxEpl13DaF8duLbW8C1IJF+uALtaHnc5x8fuRTjR/lfB9ZAlWPG/XAnqUXPN
ZTfFhsKoW4nNfbI5gBFepQtxE5iNGeWEA7HV2w5OhMG/U6gJ8HI5oPm21qYXuVlw
wLfwGTwECW1H6B6maGCgcaBL2zOYHBz+/jVpHbcrGzZcYfTRtI3K/0CCULoOb0n+
cqFRuQlyaS/3AHa7CZ+OmAHKKDU2ghiPhXrrfsTJ9EhKT0NzlZDVlNTBJF4iuJTh
n7AmVgrIdRrSmQNdOoxsM9oBmINApBy9VllvgxH4oi7zjEO5NfnE0rpTzPIIYKX8
XsMfn9iLt2WdhKEEsgpAB/hvh9U86H2vh2znXPaetrWjC6Jl0puDWuJeTStSBuX6
1bLKyGjp7Lveawqx38hiVKYi+smUh3TMtuxwrIuO0mKNLEjp4hIfi96U0g/YwQiW
1TxzgLjUZghgFhHPBtbQm2h3FN3U5gAPEjHGQJhyGZeOF8Mj20Z4gOVk8qLAq6eo
qnrcivXgLhHD4FmVEqmmzk9+63OJZV9PYOmo+FTOSfD1PWK7GV1NtS6Q4DMHyej8
v89NvDh89k/VVomYThiY9QNs+hhZ0rlDu4QVAGQSVq/aeCsMYtonB5KYdhJUktfR
tUudJ1j/rfi4U+8naXbBtOZuj1cYC1zqauwmukwKfjm7Uafap+VDdz3tA3spdAJ9
ByulfEllfutNbixb3xBJ7suuoSU9/4/KxcaE7iusBWtJiNSJDZtT9X04acvcWebM
/2JVBoeZxF/w6I3e7z+A//yJDMuaMfeK/QshN0MVcJupiXAYVDMF0l7nz4+0E6I9
ivwJexrenMOBqSCpfId/slI6IILa3czYUmMIB6DL/zXIucLTHPvEDkktgLNwTz4O
jkX1tGHSzejb8FDDSKntqpYSw3z7SZYr6CS91tNHyvKQGUUqJxlP/8snxcpesq3p
+uo2dToiD7qR3HMdvPDFZY6n0st74jEb0OsWtb8ojErQirTFikh0Iw8Fp/4SblGR
0MikzE/QxnaBTwjoeu6pjBq/Kzmm2AHwi0We6QCo/8v0AoQLsBPc8vPz3VD4MAjU
Lb+jQsSPlGXUqsqTGc3neSsJkahNE/RJvGOhZBH2H2rRXqR0bUgv1RopxMBAKoYJ
wOEXv0Edyw6GMv0kc7QmRRGynvx/d6MBVPyy2Jzn1zPnxX8vI18/FO2lfsEDXLlC
SGlieakICWGWQTJFhb0KuBAZsVC9HLk7Ly9rKDRNt6YcXcqfrgbaXYFg9WDvzYth
t7SMnDabUyV1czZZBXsmFHWGRdPrGRoSZHx1ZfHkARdYjRnJyqjWrxsugSZrnhtY
2syn0amaIshGJhQZckiYsqpZnike37qrLvRivUKbwLEflAYuYYuBwz1axhPlkHuN
POJUab3qk5o/kGkH54oUpROJajXAsRbd+6g9VQaQWERDrnIj5mdyvPC8LOdQdXaw
TqwXCucCQW1JRaKeJsESMrNURHBppC+FwOOqcdamcwWv5qo6LONO+HW+4G0C8RM3
xtWIJ+t4paIeCyNbCtmiXsMVb2lwFHqlf7+nHXgNxlfbjVdIRDeVbgKa5a19jWHK
U+tFVAGpQCUZF9OYNNJXbzFP+q+VmwkeHas1LtvnmOzzVP8pS+lSPRwhRrYMQ2qo
uvi9HCNZ5iTkCvtg+M89y25FBNgfxd8AHXoM1zw54/fh1DS2ld5OOFHVKyaSXf1/
2VAS6bjmnrx43EKJqcue9NJ63AS5r6mQIHuXK9cgUHstlL5xWBZg7DH62FAnDgkf
G4lUOqMEmUmTaW+/oNOIHzPSpJhEV6AkbxWX4rnRditpxxpfJXw5erT+DRVvUtVl
A+VN/lCaJWvkho3//kTHJ+pUKsQNgZJ1XuQ1oD1jgf8oJ0D0ZKPXFYEMQKgSFk8W
3MKKjsidMZCTG6o3PHUq/Ck44S3eZR0bShT3otAdPrcbRzb4iY9YLIudrsVeoDwc
ri99o8T/pxHua41yl9cLjObshWTHPq0tmUl8ih2AFcrRWVjg1TRFuTKL59Y4adEk
gowSKhqZjIvAFCNPKo7hKTn8VGTeEpChhsrfa5U+d2cN3VVBLk0Kx5H9yMDDD3BN
z6N+3nweifteS/OeOL+VNJDJiGWh7DLHzXzgJGJf6905fzyGFtu2ozjY55GQySNL
TSz9mHOr8G5dpiUjk3tj7Pv5qWraOUbFvjwBgwr5R3d/wNjUXriK7BgWnyez6rzF
yIIrMaxtauoe1dVLV4UhstNasUfggzj1voIXrc0SYvrxtoKLk4i3OnJdFJjJB6Op
Tr4KQd4ZSnAltfOtFh2aabmNgREWmB2kuoe8LYNDHV9TFUUdub7Isix33qYzHYck
2aF5VP29jVPHHXe7MEq8b37lhK58Tgh9vEf7zJLvRTsxn9oyqvLUWBGXiB7aJmaJ
J6/DJ2KYLnSj1aOKt+9c05jXZol35db6ZmFgCrGK47XEVvNFlfJeQ3vByR6dFzwa
yThigQUAjQjJC/NrWiO6Q0DPhdd00Ypqe8UO+zCjyC0LASx6oKiO9Z94miIEPNWY
haSHS98Jwc6z8l5qsvXbMIteLBGhGpJG3cMjFko3qT2pL0URV/2ZPKEnP1ez1tHr
poaw9//cynRmo+59jaD1qIngO8ga+oLxr/2nwCD6rSZlCC1r3DX7ZuIuRZD0GJJI
VZZQErU59yGscSjSnm98nuh0srwM1SdG8WSadsV946xYQ6kv/Fr/L9Ch6cQoZSvQ
sJdvosTC4dIcZubULKyujICtL7g5VfTUyJKRTj8/9mPs/0ZhdjkyqtZFOQoZ6oNO
tewF0iNDGqSYKeYDe13LOVsCsCPO6nnhFO7QIci0MjXhOpM2iYMxsxEk5Ume5XDp
9PXDz+KLvn+uTGVS8l4BRpXTwyuSwSNb0flmJdEv05qEpXzE4uWEe6R/f7njF+Ng
mB4Ud5Q8BHxwOfpg2v9cbaWNzeGK+rY0myAj78Ku26Rs1b+5cj1Fbvi2wDqaZIv2
B81WiJd49kxUP9Kya4o1mIus1B6u6SxUebUKzjx3ynSUeJ7zIUdcrr1i3vpAbI7f
CSWFvPqJnzpEiU3eiUpqDm5Tw2m2ITjWviF2qYPYL4tMyBofpk5yRMGkzZGr/t2N
LbeS+aAEvuvLRPuZBhV3NALUYAstSkTPerbROwY9zJ2eHNx+LU6BGyUI7A6LcAtO
UddZ5MMaphn5whorKL2p2JoepJyLcfZzP6mfa1ND3R6WswQLLfFKbglfFQBNbN+t
Xq0IhZPVvs/S88z+jhMOT3Y5ro3fOpt4kgghSNpUiwVQD+x7tjNnJILv8okEC5fE
FDbdJuTPAYPVILm9vCk1xEMN75PnZxl0QdNsF/Tq2GXwokRC9/3u67Pd6COM+qry
/+wno6OHL5RNsw6JekG6jQBQW7PgbHLP+uPutDYi0vfuzMYBdmmljGXYx6WDc3/D
isY+dL3QrYIvuZDmmGPd0dYzNJY2VWs5616CXyrvkcpx3zNzrJ/7PkOm3ra7D1gT
OLxHkcVL48nY36oFGKCF5RJqGREwUOGpaXWohakL3Bxs4/zP2tE3ipv5ema80AIo
2PYyQ6GmCwulymRBnN7kZXk4Sm3XXTtqxXG0FPbjdad3ydf6dmf2veYJzAKi3oMc
E+CNVyJB+nevZnr8k9yPakiSvZEu75iYFilkrFgkKQzl3CmXlAe74N4c5KzfGmhP
shlXdcNXIsD2bmvG7pxvFOjXHUK24iIHDlRcwP4jYBXYERL7s7HEginqXzN+VQRN
WX+1WmzAcVHLA7dlqdUrcFtHekyMZAqI0RGmZFYb48egAWpw2yfpuLoa5Z4dZHr2
y06AGDaVwDlNNJioVx3RhHIMRGBmH//pIIo/LGaC6DliDsHqO+j5xHx5OhpPGcT9
0eLC9D7+8ObJhH8mQO790Vudc9EBZCC9Z281CmbOeFlGvLOKjFiwyII/hFg04e5u
jMoEnJwrjAg3erlAojuWiigYt3RkM0Agc0kJ9RINH5RCxD5Y/BPrPCTRyyR5NhrN
TbKuELSpTQFF3Lx445FHTgKUxAeM9uTp8p7QDXImsjSQuYySfwl80mCUAOoo4HPO
xNIkWdIDSdlQVmBsvTsIYrBLoZDAHW0r1WlZyR51T2zg7SM4mbScH7WaAI4A1iYZ
WNT0jz7eMmuwlNVVLjjabirg6W3m+9LhE7YPdzhSckdcpVIqCdJUzdC6/9aB4Q+K
jSLnWO77ZcIuhaYwUzLKvrVtp9TmgIMIAMmCtUvQGeDpM9ycpUl+RF+8qjOECOHf
BEGOeRaEFdRKTWB4IMlGKL7oNG52Jrwbiug/irnjKY+dkcsqrCmdUkYoIgiHbRPQ
GNQCrlkKbu72Ej97riEoL+ofcqILERwzal3P7T12vrD8wHPfFBR5pUD/UULkYtgq
dl6+tHqLzuxvWBXiRoabjdXYlw3Q/J0oGVnqy9a+W2ZOPjDrR0vfpSkO3z+mTLXw
QhLq+s1PfweXmRfnpQD4fOnNle+bu94fEQK7Gg0+rDpqyfEpBIEVncLkI6ULf9kh
d3p6n32/SZ/lX6ysrwPcHRILftMguw8lwWgH71ApvdBbGl0zOxtE66kEicogCQ7h
7upKO0iwEnGEQ3B4ZNfHGV6hJiVGezocON1eJJaqobADmrCHPXn8otnGiKV1INDu
mbRVJbt3I4tnR16gcLZfP/vWULvJgcZcmn6asHoQkVvPcuUm5a7RWkvR7fsGHFw8
1eydttfCASiEa795/5i3ik7SehJ9ckFscqc7EBzfnp1ds73PGOs2QpYAJ86UdMZD
2O3Yp8fedZGE37ll2/iXPIZYQ6ubVdM05CpXfOV6D+ToBcfZfF9MuSMmrSEEMPZV
C3vS4PxGq2LuWpVCS+/LBRJw4kO3IbY/jk4GSQ7BJW45gpxV4n8M6E8RIAL3z17g
F3yxP+/p0YKy9S1QXv4K8Xm1slQskF59fZHhTS7GiBOn7uIAHVFEH4gnlLfipDNH
m8ZH0zboZzIdJ2BGAktaa7DEKCFg+LNKmjmCwtOazVLQWnmDJM4zUGQwBN7FCV1J
sLcBs52+xjZClb3uhtHVrCnhSl7B6zemFAJrwS9bkmHWg+OJwpGjbO6/q5NQQaei
/euP7e071W0C6EHmQOCKuZuJmlz16YFJPQWQcphiG1poLOxPj7SfKIEyvsd/ACXD
2d4uJHIqIDSmuw9qn0gq9QFeN2R1hN/ilYWGE7iGQVts2rWLrnKJh1PPhOce+aOz
Q8grWz7YdMJwg/yD8GUnQriNnz7AUUYHIXtA1TyurqPxajOUO1KZrrBeqqAQMr4F
mcXwtdCVAyLo69SN8GzlPgtY4eayh91YQN51fkEG14TsRkbA3UQYod1WKhVaVIWu
is4F+gUpP26kHdbRUxkB8sB3w7u7WmzewIGXw8FEDrHDEzz7k9hXztPNYjYIFoAL
pNqoTTa1usTOQrH+QwOOKbqOKPJUD5GsF8oO7IdLIgih705o3wN2tIuDcUZmDNJQ
yRfOHuW47aVFsF3rfoKFmZhJ7hRjUFwi1edXyDB3WOjqEhTwe2jUCT21CkrGRwSN
rqy1GEKLkeppaJUyXmesO5l5Be1nHdmJYBcP5LpEjVdAiLt4N+V1/5UXH5omAMqv
uOAcC0DkU6YnSTgQzyYbsKu/jHB82AxFUxjuVe9gh/VoYLbtR48fecS341rGs0Gg
bmjzdCKR6g90RdtbpNJVJppn1TV+tNpdVJksriDo7ef+D2zOTxKbOzgGm7XUFvUb
vn//Q8SaHy5zqStSb3Qkl9HMU4vigMDHYZYy8C7CdXkJeNehKSyYyHDs55MuA6ee
j2HPttEvh+p0kARvtJOx6MqYs1b+tK9dr+49ELrenYZYJlCLmb59knknWOBGZBNU
yLaOCI0muwz9/J9Tnin+cfj+RxHTsO6vHp740vOcHrBtUy6u0eoV7quJQuSuLhGU
N7X8F3KVGckFusXzYOBZsLI8icpSoaPqyAA1B5gNov+DqreiHFYpl27n/V0MSgnM
SlzD8PjZHSTB84ypITG3uUW7zYQVR36nr9Q6Pcstye2nS20Eon1iVj7a0clM27lH
+E+vcKbJparTBC4g1lWejfbIHy4H3hDRpihnoVQvE0Ln6gDkl6zp+gAQ3r+HSCS9
2ihT5bR6ejQHgVLGi3hr3HdcXt41htkCaPtLsQva8JgoFLoBmKTpTe6buCi0wRgG
75tSdpGf35WUDD/s5NT23gWAtYTJHAKDhLWLIDDZ6NbE53WtI0sfH4DSv7zblKYf
XpjivymN5GI7PDL+JQ0LtiHKglqUSpYh0cTwovnxM21TFaQcJ5nmTa9qBZXqOQan
3OfyEJWmDWWS7NU2EyBsrLy9obf32WdDP5rXTtz0PA3H/X69h6hryWhXucU5Pwuz
28qIopagh28hRFFJDJNepL6K7va8d9nuKLngPMT+6WJ7kXkN+rM0OBRBAynyh/3R
ex6Udnf8gjk/LxEl9yCVcRLmvjK9b2nqOl63RgnfyXd6IHpc4IXuj3WKGPHWP4Fy
g5NOfuohpXQoclCdFF05hWnQWYesn35c7ir1xTaTHV2CVlIeozQx+AtmtsJEaWeT
fJuCmPKeuAnMkOcPyxsluWyni42R/vUr4RymEyeWGhvvOm0SUYTBkjUKL4jZQRkm
vTlVPwLissWiBp8yWRcYZOvXfC46dPEa8GmO++N0z2GC51nlmONUX25JM3xvtvQV
RFZpvLYREJhwaRlncm0a2KUGyJJjzPvntOxk+vB3r8mkXLjrANaEu0TiEi/NHvg6
8hmek3AjnmbHMeUnlDaeaW2f4uzGp3qUJWb0YUrkdz8CP1AYrLwKtuJxzIfhW9ti
SpxhrXHIfVHWuuuqHGodOutROl8la3oWc5zoKlYKD8qEW+WFzDcUdcwZyQAcvqKI
0KxIHXTh2OrQ4wwjc1/HlvMy9zyCEkYvpnns9O6WfhSK/oHBsPlQP+PokuI/T7rf
d/66MYt83E2+shfYLlLZopugqcZruvLKyoeh4eNQGn/mm1Q5iPJgJTAojzXx/CIU
/z87jGhsjlFJVAvDMYM/mjT3kfXDBkfZ7PQNieXVrXB6S72l9m590Ib6G5AGkWks
lL+c1HgVDNSHPWEWAY/6PelRVkEQgzSXZPfnbukmzGgzsJi/jO9nBhSTyqye5E7U
ECXdWFYrjKtnRnBUrvFHkQp/j4czoqcmsXIMNtwOOt2atKcV/jEa+JGLMB14hjAU
vE9KcnStpjh6DQWmxaApAdyRc9W7ma0i1KSdoltxRfxo9s7fnQ3BWhcuGwYlrF7h
NKLH7Ozbys/3c5NE3RvLCMnG3XJ4OF7E1EgHva3XST1dVyrBIf003QzVcRsEuPIt
DJ3kmGwLb33KA2HnwfhE6ZpZLfU7yffhkmV10tE0psimT2JQ30W74AkDc3oAOIG2
Fnsal7/zBaEjXr/Gy84VzbfNasPLqU+ELk6hwiVUzTnqVRyfAZtAiuc5sQOiAEMY
57ekQCa8k9dVJ9Rt1IXGIUuZwCfc7s3PGyXzgotz6NPG46GjGWGo55j0PjhfPE+i
CG7SrCOM07PYO2ktfCCagFnBUPgVwpBa38Cy8lS3E7DoE7C8dBJPV3N6yQydHi8m
SNsJiuY2xI6J3/0CgjbMJs2+RnTuIGH2r3CcOba3NMkKFeluta3oLv2WcBORxPye
oiQ8kHQft3Gck47p5EyORVVnUqZLOO0SPeEneTexK54KMFnNxYxpll6HCADUmmGm
1/lxDkA5nLQtCEWrevoTWBcAcdk3ARNGamSHCO3gV4QurAQzo5uc4aDVlr7vAfv+
QHyNuQTYcRiPdGGm5293iRghk4MLxuqr7p0QrxLKurZMH2pyvy4YIeq/Sgs922HQ
m7533rT9q8MGfZbGk0BFh/YSmbIFHAAYxph4h/wMrN9HWaJZLeDxzuR+0/pcLD6y
nyE7Ek0iWnkX/xEvVNbeCGI6MX4W1+badsrn1q3L4LM4BFOykUkT3zDjJaFN7wAc
Q6b8XkGgyBqJI2qpTNxIDyvUqYC1EPV+3HwFHb6sgVxsWgmzgcP0QW1lTauEqpeJ
vTdNMcCpPIS2bTxP+gPUpXXs7iyHSicTag3RR+NTtFqZEMPOySWhl0mhigsxrC9a
epEbMUtmws0JIcqtWxccD30bkZwp5rVD+aLCJQr4PNWp4MCW/D+PnuM6ahelvs+R
PoafyL+Vfqn6sDHiV+MSl1jxo8Mq/zFRisRJpbqvKS+PzYUWx2bfqlW08fvs10zN
1GLGIAT7KhDQy7IHkC7YQS7BkZmZMCGZgRr+tLSNz5VneHmXzuQga8BsNKtv8Re2
RdszmUYcwcf+r3PR8hLin7XXk5F3PZeXiXiyrkxtDCDaY8fnk1lv5MdaEnqzHmn6
W8EzIntqS0JFxksVbPD/H0xjWLZDaMcXJAINC6pcU5jzjc5os40u38P2GRZv/zHM
xB3zNUdkCsT7eAJo/FqtIwXMvjkCKdv4lk89bHSpyMzODAy1voNQ/RGAvjqQZgyC
6MuvUTadCMkXYmPaz4Ws/77QeDkG/CL3zrJY99dRLNTMdbGgBYp0c/P1ZQ6f2uhm
ODiYjg8WqSf59dYdzcWJlwQ2up+Z39Xz3g5/uxSW5wFaiuSlw2lkbi2wf0OyFrgY
+s4xndBcuqW6fpmOCtWtrRc2jyZulFHpBtujSnvik2bUFaA8IqamP+2he3CxpMWH
xFWPMyE2jnXUIgU8hKMwkpMtxOxVzJCmgwHAXi/GgMBEgetUEnpwJkSG+gaELSKo
JJywbYNMIEO+rP3fJx9AJTeLn4rSLMJXfgdbxC5vnJyTXHKnlo3AnHw60t1bHbNM
uidbdMK9j9yBrag+JARHclTfUHuzvyhL4b6LsonW6vEGc5VYBOQbM43XDUfKOT/4
PdnnQ4T33tVAyrIQIhyydrnlwvIlLTHGtKxGsmH3seuLetfFtqgxQ1+hSHJMmO7W
4qLmf+DYamsjiH5+8NtO8QfMqg76FOk3dovLt9uKeySoKSbfSrumZazkjBA85Yjk
7L794r0GQ4wrL+iNxCB9dYaR4fKjLCQZsc1NulnjyuaOBQ1uHu7HpiYbk1vNbkwb
6zOJPOQ2UvzvyZq/a97b7iyyCqfKPk6e/MJodqGqHNNfbbvNMa5BtSuUgopAxhdQ
q44dOg8IZLMx7VxRd38HxLB3jp8zvvw7H0HCpvblDOw8jGSpVWQG/LxRTrZn6SYo
Q3wZzZZai4Kb/9s6XzJdDIoxRq95u46ESHdu0aWel0RyDy+q1r1sDWNkWOeFR4VU
NUtXxQA4eDU5PQ1G7+cI+u9Kb8AS2A92Kj79w58D2GpPRoedOqOkwsxzqNGdd3na
Rl5/ymUSXi3CaF8JPOy0+xOh5QH+3bpldgqpvoJsgk++2K5u+30uu7LaV5e7LdG5
inJOuZldX7X+FyCR5p/5jrJzPYqu5QCTw+b+TfuG3xnq49cPfcCuNMHeLWBAFpNt
beWGmfB7EIip5KEorD3Aqug1JnmT2ywpVSyy+jSQ+ZOg5DjTHZ4d13Om/ij4zjWi
bUQtbqgxIZ3bSKGcQ3KciR8ngZbAQ+GBAerERZ9BvVP4XqmlpXFdA3G4LFGItcHa
Pl5Sasd+EmwgueXo5T8BZNp0c6gbRAjyyUWgLaNgVJSpbaS0Y0xPYu4cxzJUsgQ3
KcNh2cRug0FHHK3aNhz9bCUim4usahkxbeGlRn2KnQtxbd4eSxtdDsfolfmysTS4
1TJV0zTYng3fjKj/VUWiIJgvmYr+AYVDo2NiQP8bD/bcHoKOpSlo/bEXOZHnrjOL
24I83tPgAkeo3NjC0D1uBqA0lSQi6Jr89u9KG4Ki4pmZ5bb270ELpUORNTY3te9h
dW9jbgnZtI/kP992CTFp0kArkoJTX7KXh1aDNfE/FTRsV8sfUCe4b7A2YhVoBqxp
S5vYg2rO5liapVcuCXl30VR3FnevI7bJ7LdOkkTmOEy41BuqMbRUPXDj+LJZPzOu
RReAup4ph3w5VVoyLmfxoXwFcVXrKTOLb7OGmsB5ekznKoz125O8VoWkr9iomVnW
rub+rgeG5GbGo7hgOVMvAs/essU4JpVmxXzp0T3MMHM/sIqmw6ehOcA6AvM5h8LO
wLSiD5QOgeqvzhAg1601DuD+FucoViX5oxkBJ1sa8UPYZ9UPFi1tOQgfSuob5oVq
CjxelrzONxpvc56HxXqC+22Q1hfqbHDtE9TXoRGvDIlDRunjtt7DanAa9x5qLILH
LlDo73GuW0/gl2lGXX1lsgRanqCT0Mxo1u/dv66A0IqnoDtFqIboOnZZoWWRhEIF
SwH5IrN+38OeDmQxxaMFaXscRYy0g8WDIP9SH+q4363laR9V23zMlVXVpDn+qqYH
Dad9x0sT/GOzk4W+Vs/YlsfX9yZM5VaCESL/Doxhq2iqhYlDiAhKbb18PE8opwCN
jmGcjH5uaDTwVVZ3w8OqTsycqu8ctjsruwo4xPFiYtQyvS+6d0lO1+TjGBc5B8Hr
IP8yHZza+oz62k+1ZgAYCg+xr6KuVo55TkcHTiq4/IN/aAOnBCO2SMuPGmqT9agz
WoNnR7V5o7Y35L2jsn3jQiU9+RavoKfmr9MrwnVaEGA1YpuAuD4BlEosuijGR1PM
0pq58t2MMrMussiJ8pCaVZqjCUifk/yVFJ9AaT1Gq6jCO1pV1JgiKsvNXjF23476
Jt+q6e8vV5H0Ki2GgT7Waunr8b6LLqdUMSIm7noYDBMf16rvK0PFwAenEHS64s7y
EdThY3n2n+t9e6JsAKNsmUyQth/WfYVhjy9r05Cof1t8Oyn+o0GJtrGHkGfYa4M6
Y4/yEiFIzKZjZcZwBNhkV5p+emz6UC9OQQL0f5B0fGZ3hcBy/Jhw69EvpYA9yyEH
/otUQW3GNX3Wdul+zUnLXoQ2SIcxbjt45l8bY9ogrcK0jynEn7M3t3mTT2k2fU/R
Z6k/CmirFKZgt38eLZaEOAmCgdFD0EH6Z4n4nm/mfHuPRQdLuhAuxJPyWg0rjroA
xagNHW1Wtn9deIGpp9L/RbH1rwy/Lz5BrJ529c9oLuyXFocxfSrh4J4XRgMTP5t7
eCPLTfnOfhBgqlPRPTzjdyceDvkJM6GoZ2BwX5HgDvljgLv7vJR5vD05r80bscFV
+J8dNqF1Yaq/7nEBqpueYeLGTHcppg+mzSeN4GkGCkSdaWgbrMxhZoADmXmXzWeE
AXjIvPeBvg0GVZGzjzDuJfmJ1ybH1917Q/C7dS5AP5pOw3S+GzIjp0s5KFW5UNCu
uYu7EKcsh0BJNgJSj7TDOjPqrl/x+/3KfwekQEgX3+Gp6uOKQmw8bZTjw7b46Xsl
DA8YbyIYnyLZwzX0aALWt4WObMf0Nt1JMDbQnVCRNt0ExLl7fkwPEUM9ET66c8s3
Lugr9LBdXwYD0CzldQ6x3LyrqgfloFip5G1p1kaVlo8fx3vWOBomsis/2cAXBA3w
1BgmKPCtylLS4a4R4ZsXrl1IgveCCEWlA9q5oLhyMuUFwFYkVyTRdQjdxuWWv3rr
NVbWwzPwpurKb4L161KNENe6g0jNRpDTSqEjD1IspH/mTbWs5gDOBlu9/521lwp4
vwaKibIw+Fdhs98lBtz91P5JwVzwrwxL6YnBWy+7rOdbTb5BDtoyR163EThNXsTB
Z2yGlT9Fx7ymB8q1Rxz0KhVaWsq70vcA+3kUE2ntO7T8N5Lmhb/+/JFsNdMPtMHp
Fkpne5BFDWjhrF55rOiR7BzlITQuXqE5f2J13+AhTvkJKcGn4ucLdgxzoXccqXYC
Ykym/DRy8TpHNIIRvlxEdZ4e4c95Tnsp09RviJpcHuJAeOUh+KZW9QZQV1EtQg57
eCfqygLsSh7G3duia5LAnTHJFp44sspWy+pMW7KUtgLGhNrfD18TJ+avewKQ6OSG
n0EP7mMHU8cSFy+fNji5mB2B4a9lHX2a48BZF9BDOziDwVEP3k8I67FoooVFN/RM
qpyOYgygTiV1jByCx7yjuj22LybpVpscpdDKyTnVRwynpCmTFIewTw1Hb+WOocRY
BepBaCALmW4QSnnpecIWs4RYN7RxIKffimEckmgbHHuocfJYKZJrM/sfVGPAU8/d
5fEJjydWhbX+0MU+i4UtSjgILYGGsjleJR48oFI1Ff25uV2Es+2oMq1D/IfQunlO
es6cYuWsUY156AIGBWY1X0EOc16ZFZSnax24Rf9uxpf8PL8OqZxod+Ua2dxZWHFR
loPN+VOacMrjri48w8/qWLqmR0ocWWKZ8zdR+nHQSZC786xAOL7yNrUn0nsMztXZ
FWSIbCTxq4Sq+sKx78QU8+MiIvjTkSHi5HUpPQxwux8WvoOkTiDHq1gFzHYBhMdC
c+h/Dx8QV7aWA23GHq02F70hL4eGNTSQ6YRvnprk6U0l2vk/OGFkTlNroRTUQdK/
lyVrT8c/aTB7JcIVhL/wOj1P5jyEsZD5MWMMb8zV8EV8MmJ/iRmLrhjQ01LdYCdY
znBNvSL31fqKrpln5B8fv1eZ0xCTA7WfUMlW7DQfgjHCQwzlf+A5vfmnwmFxWa6C
H7+4iewoVNlJ1GfLc4UnQf+7IOMgrL52JLAafyBYejRUFvPLw8mSdVFx1CMat5lO
2NBvj6tb2PbUvlWw69Hh2wR9vluTs8gHvdMrmCLr3JFnHdLMpI6Y9xVXWPegMXoU
DcuaEAmFat/1y28ZCsTcT0yT55o5IS3+tg4yfAqVcwfMp8mwaxsMiCoUbNdH5t3k
LZokYXeIIP3M6gOk1tnAWmHVyWoV2DnexifzXxLXAhZY1lQNdOYKT5baoJVNLMSn
GInDUtoCuceNuvJJkghYJm8OfhgEwCh0j6XtVV+Kz/RrFqN/6kuYRaO9LVuBRMhb
Xk1qbX88uek2fzrIDhOVfBjeDdnh3ZvU8QpGksXheYEvT+xrm/c90TrE2J0WwMIV
PrGZAsvNMyiLf6kjOcoxLlORcbBRvdBCHDpEcf9c+rn4ZljjL6btpAEy9s2txXfC
diCslBzEuNN0H0SjTyI90SHYuhQYx0kTF6NPPRSTjU0wbhXAMnaD2v0H3m19wzA/
xIxwVkE/1DH86f2ghOZdNQ4uDXQQ50tXdN8G++03t4XgjWJBiCUlEO6uZfdQZdDL
emFZgTHvEtbtMly0Zsdp7XO/cAlJ4wE4DmREynnenS0Tm8rzNs4tpT8byEF2RfbZ
MKs1Uik7hXcVGHBPwZJRQRwtXiW2f/cuWoOgn9JnUavS19ELBqJi6CDutx5UlBps
SpRN1CAQi7d5UoqmkD32W0qClzcDpttgFIyJxkZqNvjD1YgYrOdtvJNuA08QL/O0
xCkBH0Vj3uV3gvf+5156ZKi/GwU1oGUVVPMZAU49zVoux0KVRmVbW4z4N3u+wijV
SOB6LJO0WQzS/Q61hb3zw5L1vkXOacIQLRAORpLLJWAs8ZD3EgNaqHMTP/I6YE4j
HWWQnDiHa4eI6j3vJuHMuVuicQdL0EOpa2s71/aJiqOkq/dLTNpbiO1fqvRGWVgK
ygpt04i/QOE2OnnIjwMbd0EHGAmSDjs9Ul1QUtTXoCGBZfbsJvjsaM+GlZhhEQyu
tGVrSI5v3KO2dqL5ye0O+tSDV7X5YWMyKdL6myeI/cxCNC2upOpBKe5J3QtDDgF/
3iDnj+V35CRRCK+pRrai75SKBnchxM0EtrqocVhOMGl/1J/2v4NLJFo3SL8hvSEr
pdxVYvsCtYVeixCGY3DMxI9PW+PLG0mW/dkh7YLmX9GqudNIWU0EgV87FffvfRyx
5ikBdokFDUenv7okHUO9etLQHArlXGNRkYTky0HmQyQGRXqi4BVGM5HVUVfH8jbY
uSfp4u2KDAv+U6y/72SlV8/ZK5/GxNPP50y5y7AITleVoirIbB6FYYZKAJl5Mk22
LZucYPjqf1jeiFX7wIbHMnJOFGQ6crdMPG8lQbHsQ/kxidWGiknpdo70yaUPjkhv
SZyLPqThgrgVfEsoXtBAiyD36ER5nMQRh8AsN/TRrieDrE2J1cv/C8cfqU07HPOT
pnw3YkzWgv6d8qtq6mJjJxkALUJ6Vn/ubtjBoTngrCdeF8DnDbM2N5J5qP5KlOS7
pismr5gBe7u2IToYOMLIQdoZtkyZRdGqHYENClGZi/ryKWy8TuMfHjBZeKme8lKC
OUwNBhvE3Erk/Y8ZfoUdU6kZIjvgdFjdzDuwQJF1s+Te0+tZQiwKLuUVgnyI6Qs6
Cc/94eclO/SWdG0A0YPBUZDuAmv6blcQRgvdStaB/UrNHFIJym34BXDWTDE+xQpE
Tihcv+Kwytmv9oumxiQewM9HOzCzvBhv4Ki9Ci4siaVbW/rgftqGtoPlaWjC0jX+
tAZ2teuMVhb4MZDAji7GypOqi1M5wtHujYe6gu/aZjJ6pnRDvpWngJ2kkE/Kke8g
nteVkIz65iiCNOq1LAwXWc1WnpISqS1EhUEnGJwRF61VqopfKVSd1/HPBVRqFlSt
7b188Gyi4DLFel/PkuVpHDzksYZSqPz+krV7gNA5u/TIsPL7Y8r4yLolb/mh0XYl
4Vwg2fmvEhGis+aezikxffZXnEFR55FRUDBOU3TubcYaNYrnhPCsEMeWe0CK35Fd
ReRoX+sUqbHVx13ZEzOsmQZAqv2YUcpA8fIAce4LAFK5u47uLXlZzUX3w6+s7jsk
uUgW+A5kc9jlvoVmhAEGcrKqU5P7JKPdn9lAl6nUbBaiduHSr3jYQQ7i632GaeyN
1cCMSGbTyMkX/pMJwy/h6gQFiOFWO4G0gOaZ5fXGFoRhztQP+pw2FT6JNCQd8ayt
oHJHUDcXzS7GHuA5lFdy8nq89CNGcgfr+9YcReDsfwtZEhRoG5IEAYmyRciLe9S4
ff7yz65XmaV7jCqNwq00Tty6qdU3su3sdp1esUQGM/VXReQvGbdg3iWUN3aOGdOR
WXCxjm60fs4e5/DSH18Hi4x2ccfElkUwt8jOW5bP+90a/499vJM3up5rdEmMwtLQ
j6NKHH5kS7DowhX189O40PHvaEIOKTWT9Hhkvh8N3x9l06t73iH4tbgPHKvEbXT3
memZQPsRCdISA1Sokk6EDXS1pXdcfyWuXJh53dF975lulDkg/FUy+We7SH7blbFj
Khla4sEHimN5r6xsihqWK0/4DdVNNa3L8ss3NjYWglNRfkfXJtJoPgvpPvPoGRfC
iXy61XgHmt45wBLeezHeCCC+uesk7TNrbfQjV8SAFVkNd6QWr9tT/cIy5Ta01p6X
TRNlosP/UTtoR7AM1LdN12ywCnZmVvKi90LqZ9ZawkMHHX3Wqg306oWkgC9iCjDo
tXND/U7b2ZecFWNcLL1ytubsHtV7KIvqLHa6TsI24VEsoUHrrUWRwDlthdCYYdEc
Y9iTp40Ifj+Cz6o0kuF9vmezNBXIIZorT5FqPPf8eddMOmVm+bwFSTj4rWsnNBQZ
NvQut7TbXYJoxB35aJ9/If8rcjNMJNUwBDVRgDRGSd/f+BF5dQ+l7zzdGwhd6eVx
gv1TnL8N5g8RBS7vVuiGX2CcoCW0k+kCK7V8kAqA8M2rFGsGulZc1S0KtixzCmcw
9moz1Yn95uSfJFrrANC3IZrUHrA3v6vkyvZ3ZXvuLAXKMlJ3r8lU/BTwMvDt10S/
YuwUjQIZ8L0r5HuoMQiYdRJUJ5M2BFgZuWm1tXEKRy/PiAeBCqrUEawT4fL7yKz6
rZfenZtWffXD91HEjAg/JkDrY6U4Dkj1hzsghf8d0yrmZub2yD0CxpLqUkLUqJ6L
OUBvDVbTb3VeEJ2+d4VJBZDV8zCi+fca4yebegAbuc2C6/sasNLkXrzhFelHLgLx
w1qqLr1k3h0pdi5hDyUmULdaw6lEMEQjTmYOhctO/bz/LdtN3VinxiQ7vYX/3FQZ
tLPu3XZ6lLyC5SMxp0Q+avp+l85mmQTLrC/y6FIXQTPj+/HeF36X9lSWZ4VKpvap
bE4HWyIruGVBuG7N7WDRm0gUbg7hf1+H/zoqQ4aVsEdisLe6a9K68CKcVBoiYy59
f+VqFObih8tSiYHaV1A5hd6wYCudp/WiTNJJ2I6S9v28foefTM4srq0Q50vimPku
Y4ZFctF0MFPkoYfGHfsjp2rsBBuMQsMekduiS+l0oUnsfp07SaiONWPL6jBhTa8e
NqApZxGRiO+XIMnoIwtKyr7F7N9dhjd0I/FqDeVbJ7dqASfjB2iV8R+lbf0Az7Fm
n76kGgS9cbfANjenQdcDc59xqcC2I10DhN2Tkl91bfmAC+P2rQ7BorjioUuWSqql
9ItE4n4MEU8sTeEtal7xohmjkDIgRS/3o6+3ZpgdyJX8iO7M+x2ViiXmAPP8Sslk
LuSn4DqoLVISXUj3CjLGdfqZKjdaJ1fGIrNENNQAFKZr9kdwgSOuCw5XF3I2U0s7
afBiEE5Ab3Es/UaHSx8SfDm/QXiDU5D7tyZKJDAT3G6tgCJeV4kUONrKJxTFQNWu
HqiPfpxpR6RpSf1dU0AzOpGLdNcVsjYwZVo61U1rylp+O5lnZumCpYPcei67+IMs
ZpYAYFlkbL0HejEe9kcVuEbjWfRg0+Cj/JglGmdDUBnsqDv4SJIinXJvMVAN4ZbD
S+04sMb+o1Xr8N9dM6J5QiQXNcxUCqeo16o5pXyoPtrVGGga+boXkfY9qsI9W2pY
PD3PurgszXJSj02l0slOdrox6oK/+JRNqQnsfaqbR4g/tpi0qM4mlfz3BPoQn9Rv
MpADePl+ikTTPgeQUppPTBshXbB8fhHqgV9FUQhMaMNlXJZuvAZRr8TJYUrSUN4N
ac/qdJ1EqdB++vjtayLbALUZhl9b0a2EwoIEzrxAUJKTZhe9Os9DGBSWdwR1ZbmY
bMTiWLKh7jGgRmSCOZbzg6gqCcCwH/vqvS3q2tmy6uDsqPar2/Jvq034PlNxAfv+
Jh/EJc7n/qoDpyrW/MuKQEGNb+M7CWBOc5e4UwB/aU6uVVQcbxgPdU3Iobwe/8gA
KLd4eqIlyxnCsSRmJdLuDHm/d2v9EBRBBTF62Z3RsTv82ISjBJqGDiTTgkNO3CpB
pP968OGm3VaDtXGSzoDftGGruPQg0UMskSYG+6CkFCKR0RIFKcb8k5VFf4QWpulF
ABbOUOYfOHHualNHO1lDjlbyPQY318iZYUbqnWKrfxoNnI9qRhpDJryE/02W+CKe
/DN9Xoms+oxtukCxz5C3TBs8g5nsUbif6/urI+RRruJPQ8OCYKkyScxrePa6ndfo
XLYwVc3NoXh4AdYj38LRJ4J55ZWuZEA0HFwDBg6q4kho+aHNjAsJofFUJdlb44w5
OFuFGVQN6UqJT8r3w/6CDLs2L1oLJyUGmtk8hR9jXFWmMHiLWwB0qV/yRGzrxPck
hXHVrDmEHzp4OMb1y+zAElZmInGEd3FNXsHdp8JW7r8fX38KaUTlpXvqZXBu6zB/
FmxuW38U0II8/cPEHTtdY0sg0mtGwaQZMkEIeMIrFfc5fZW6kd2zJUeXRD76KReC
JbhntzDS54UAsl4twXvGxPsVGHrv4iYbYJEwcOLZLZre0oZnXf+p8jMeIifMZzL8
uKk5RHgyK+/6B4SAR58HjV/L9IWAhBv6WhA908I5EMhVsl8/X7rJSyNHGOH3CPzd
etvcBi01h3n8qt1qrPbtAVLgLpFMBcVmc4mw9MNVqk8XMiNXXrNmwytTMa1XQ9AT
WekWeTVWjayyVDRVlLJKwJ/vAw0TJqu5sNPWao95VmBnBl94z8iJct4IlXAcOv+2
2+ULoNWJtJVe/AwLcV0xuFus/5jo+K3wJM4f9BVB4qQCEaZPgXrxVa35yVwJ+IXQ
TXORlWMmhCCTYbtEY4WKwx813GbugKTJ82OORYlIyG5cPyX+F0pIINBB1g7wC+aC
HKez65hB1ihxSoLmLezv9qTHpBvi9Chqo6kODS9GZgilgsQulnvlegxvKPu2gjZn
jFkg9Bd4TwjTiSwzJD49yvKqPqi9iLzSApZYPBfEmDvYoQOYYAN3RLXCudum1V3i
kmanv9URVgFADI2QZ6CYLSbI5HUNigQGOF2LQH8Z3UL02baIsmZ9O/+9UleZbyga
G+WLwJr5/vHGDh0o71Q8yn19EIpISfoHh7JoR+jOP/pv8EP3u4uDjKFx1eAiEESU
Z4Smkytj5Wm2IoSGB6xHsW0ekH3wjEzaM1saXUbTb+jEFORfrqIZ+hXRwvQRIecO
M6daJ2Ok2wAS+PbZk9kTtBuV8IQfsBsVmPPchAmORd7Z8BRe3+fYvE27wx5eNoOB
7oikmbz4qoFT1rSCtZteWP/zr53szkD/KYv9Du7NKFMYqGA4I/9ZkkvMrD8soyh7
nhw7Sb5cqubswnkn8CVe1aonRD2lv3j0ckgc1VXRp49oYfRsdkRNoqGyMg4miim6
8gY/KWl9NkH2kCllDCIbKmNMkpWWsXrNRLAVd1/pcnJZHx3NPLkjvjRN95wCCLcl
f5PfB6FAX8BRcTwSSx5VcM7w9A5w1lSsKc3qlOz9QCokSuaw99ySFuQMheivu/03
mICHNOebQW9YfUivlmr4ksHz4CilTtw6Amb6NhO+iaBYpMfiMtvqoTlty9PuabM5
+H+lPD/q5qD8wpTm8vhkXFkMLiZhsc7VLvAe08NSFA35+my9xYq2KwW4r+VJrnw+
RtldgosIsLo2yzVoYF07GL5MjBTy1BzY1LSuKfNMxKxQDcXLsC3bwCLz8B4LNr7s
bajy8ClGO3AQd8+6fQrsX1c5kJWCr/ibWOo2xnh8+oAF5jQk/YZK3M7AfrF9H6Ee
mJK+6wBFipmWrTND+V8ypsm3+a18LRyeifXZqXghTyULi0jTZzQw7w23g4uh43nJ
BccsefGRByA66fRR9CW2O4xcjuzttrdZ1yjV/+uzzkY9t6l72cDfevzBLb6ESntZ
0WX+jVup17+hW8uCBrZ6UFB94PWEiPSo2OhnPaNQOdC63pVUlfTv+dpCZA62N+Um
s5m9fQEiJ2JBCwMr7mA0h4qtkY/6BicSLfgpw5tWyiTkerdUC9DC50LyH8c4FdpH
17wccMgxWWJfvabPkcrXKg2I1SWQsyM8u5lY7GeTGnfarKxk6BIq0TyLZP4sq1aU
RhO2nS95A+uFS2wYVYqzPJWUvkEZjskWQ1U021Lkf6Cdun95ubVayMYq8VuHWkXz
zRPSPkgv8X/Uv4CCZXyg8c0TNnt36jOPI3lb6hDrpGqUsuNbeHsHFw+5pCDIVlMx
1pbJ1/b2Tbd21NdyP8hXA3PSATbyGzvZAwHJb2/5+qPCNTWze5D4FlBjU6ItdMmN
rn+qMUcS6e8BS2b+74CpY55ojJQQUb5tAEmSERIwy1Wrwkim5j2FtWZsseHISHFI
u4VuvGlXpE6i+RQ8RAnX6bUiJpIk5VWAatgd4j6hvkXp2xObYyqr21Q+20/E1aqa
c9lSPDPnSrEcS3viAk66/ZO0J/teKLfhBRT6aBGSnbV5ytN7RcXPNt7ngD7TU/72
/y5ACVILnCKpHZ4Me5qIlhsvLq6vv2byMU9IGtDe1lfHzV1ToqadluYUekzQL6A5
6QQ3a3dNi5RHrHuYFY4epY2enAuPKZiAeiBhrOoOzYIfK3SqdA+qxD6bFK8xl/zp
o+XwG5i7BwQzgS9BQ5jlzTUtR84uvwmAxd45Y+pM2zhgUxW3JQWo2/pQ9bPnf2fq
pAxlx0F19yjBDVQ6CDHk5k/iUUNOG0zsJ51jncnXCvsXUIRC36yysGsjSQZNneU3
q3zX+AKOR8jcOm+3E6luZhG6d24Qg0prl2USaNrVfi4b4jhfTxN3ddZ5GWavSz3f
yw73qg4qSwD9t3UMKQja3NRSvnF5layoE8noC4Vhal0gTHaMuWfYw07WV1f6mfJF
CP0kRBwdA/HFjf4qH7sdKlWl4AxfRlVMnicF8zPzseGxoIXSdppKwfwiT2zAymI+
DFAFlkYsMPesQoshROcUXtv3hR9gUYSurJWLWGc/6AfKV9myHEnX0/yMB+TD4OvK
E93FLWG0ZcWe3iLwrL4qthUX8kY2D7eSqa4/qSvx751aV8MLX88gyZB0XUH+T4ag
xOUJ6/vP/l3m4optbwiRdDWAMPTIJsMXDAaAIaQVYL/Kmg10CjxBI/kmjIDWon2x
prTGdFfprN2TLPetZ+Lli8O8Qqaa2LZLtLS/79s5T8X/joWTPKSQkvCGyQcRtyhL
cEYm7mVSgz9ey25wm1bn8/VTw4dW5/Gr5XExxIIUS0i9PmghOPjzxwyBOuD+ripB
NqvWMP8cmFZLHD+um/XlJc26AO4gQTaFgHQDABbhKUlfbP28s572NSMfEeIn4Djh
Ve5gc0HveAJ6nCoCBnQCsjIM/Xa/Bmsk3qGshUSbRvHw6Xmx1Ft4Ue7udeSgX/vG
habqgTja2YXjxVOrX9386NVp8K6386vR4bG6DMvoiTxenjFo344sPSGhZ0l88LAx
MMQ1dSuFRlsi3v/xUIsu7D2DVnhbBc58nHJkQIxSvZIyfk98eMrZOVj8GR++Vdg+
/YMm404cHpdUQfS5Gy/66wFxHXQUmmmU0W8cEnMZmy8B6aPN5uhonB05D3SesPvQ
aOOctrpwV09yd5lKt0gMAApL+8e0weASSHIs1VUy5QvbtHq49eowkJnxXSfpr03K
5X6l3kfQZxIC58woqYxNvlLAdFuVG++lg6HnduoOJdZ7vipik/orMvU2WRJ1FW4k
AXYsIipQlK/ZPMUinuLNDC1VwBLfYHhBm9V0Z2gcb9FGFzm1bNuPMULLoV/HwIbo
OF2zz5+kzA4tw1PQk8db4c/rFapH8G4LyqP/+4n7GrbNNm/GX6zHKu/QOmHMdrZS
iX/7D+LGjoJJ3hKf3j+ayL1W89OKBlgesnvReicrNDWS1h5c/Os+Xcn0wzdeRdaH
uQ5HiImM2yVD5SeivPJvuIxE2B/5pVt7sTexmVoaVV4AGSRSRYmVFlPdNsUHgE1S
huvTCyOEuTwfWOPLcsbyHyqgsxptYvtEeTCH5TlsGLskdjhL8nGj6WYyPxjZO1KZ
36cQe2moBJ0l66rC/HgnNELaLB6fjLE1XyjzQYBKQAcN5HTRjsV9Kr0P7g5Aa775
sGDr13mihlDqw/NrmhfHz4z+4S3zfSL2xEknwgYzNPcp7znG5MQFsz0mWxCZrt+6
n1NSUEZABaaJpHhNU+j2QJGgGOHrqKdkzpTpg+Nuy6VnHHLdqGsYerFOUsT5qnUK
dDDml/r0EvQeV0tAac70N0P4cjnIbrNEe8YSSXC6UdE/n5Th9ie79ElU8qKFHoN3
3TSFHP/jORJWxuS9Zun1UcQo57WY+eY2A1nI92xD1IDqJlnQw7PVqFE5CQ/3NS/L
PZ+9M6TtgI8Kurrhf0Sx8y/I9ohcNVj6v8jULUzhiCFK3JXICGCpCoHJatcttRzz
RX7P0KCpBCfAKIK9U75INF0UmiIQZCGlp5sAzhDKWIT07MOhWOEjkUH8dfHPCGry
6fw/0HyjoCjUUgM8+pbBcNv8fib2ioLSvM/qsjFNXNit4KgEdx2ryKcegXXxDzeW
vKyb9ug2PfmI4Q/WBo994Adb3pLWXGDa14/fc7GjxCGrVbUgssvmJH5bL35u+MNa
oiMZeO7vTIBeP3kovZ04hEEqYQp7XiVsQVfYK/RfCP5zrdGg3k9IcVq/o6ZXwODK
3RW1SUMLSUDjiGCWb4DlTQfoT9w0xDtryAr9gnytXSYhNEkl+e5dcw83q8N3FmNI
OPPMIIx8ghi7Xt8DPmaA11TGejTyn+Niv4sxxFWx0FJMLZbtG+aLggYjlEOlalXm
ggkO+5o8k2gnQocN3CcNp3Je8BqkV8AEZUOSj5LzjpHBDwuX1Qhv8kUwKFLXvMWT
D0dBhE8QDHAnkhQAMqaFn6tJRevhvmlI/0fG1sBUNBYv90l5d2jqSRTyNnEyhPP9
8noOsvWC17dB4p1iBBMxe8KaKaXbrDID8lwlzvawS6xEfCJyCrKXbtIrNQ34Gitr
n3y6yCK6G4F9yoeLmU6EONOCDO61wugNqHtnz0Ov77vCixqjFFd8MJxkLPKjioK4
bkRG/Regd5VNWpfzWYshAc+8AILth27V8hhvwlGgP6PiJq4oe29rnATMmtzA7LIv
EcXGfpjqVlee1VP3hQh7kh3eCotNP9V/oQ8PijMBlZsZPcnteMxFJJomSBXJoJSL
vDLKkb3G83lBaXXxb+NWbrxfq69GO2FC5p+qN0r8f/unFfrVNbwNYgECHjO56RVa
n/B/tNvSd+Ib9rEu8LdoGc0+Flz/ulnWSRiRuWd0pEQVIeO8hBxO4wPcgzfigGzY
LREDg/IwgoGP8erXqaSSRnMhjFHSdRHlO1qipNvNoeWrmJYH1eFHjq9NSY8GiOKj
D4vwPlYwucf4+bw7BSBOxjF8UhaNq6bhpvWfB3iCbFe5UGZfnfa3TnUk8SN7JR6J
O4nVHO32SlE2/FlqpJjErSR4vU26xfHYwDIaETnnOd+Jha3o6+OY+nM211yNkdhv
+mu0Au5zPlFYnUzWw8+6Ukytx9sqZTQGBaTfjI3FtS7Ul8gYDNUucD9vrCFnTuiJ
M9jxTZ8fXFC0GjiQRR2zclmMwJiVe65n+S+Tm6I0CvwCGPJdlAvx3InJ1SJOm5y/
O4IXXNbAXPPlBgPaJ9NYYUF5emLAkpW3NcVG5qZsZVZqP1TQcYlZrQ7lln3mGw7J
p4v76r9J7z3elDYWxbFHqs75qQghUMJWaMODc7C4f8rHEJIB4Mqozvc4nn2/p8LF
FBUMFqhJeVfkTqpOesPDz23d5p0Q1GM1UWXcaGU1BhWZJICSHtT1fZko3ni+l2xE
2XW8oP5HIFYvTxnCPNeFkNGC+ebM6+WE/U44WPalCFFsPtXDfnwftdqyssaE/8UV
uTC7vn6M36gClWx5gNP5cM/Gu6wP0mrlJXyn+zaUtIaJB1FbP+kF1UCQwlbwrT1e
EzHGrbvrO/JhzIrT90tGpBe4OI2OCQloPdgXy2fMGIpkiFqLQZkVhr/8EKGNmBAI
jfRogIPCSwav59vPwP5mFPKPzXT/piMmld/XSZcaN8O3Mkf5rnijFoZT2icamj0P
80N63671zhVvLlqMCDmjK0Kn5NJHT94lmPuiVBH8UrkQabgivSa+1ytwWLqrrAoB
M4HTYdN6o4RZEFybzexLGVZ67sH8aRISnGlnNsACu8u6kTx6QMNbtdJwIeHFvRao
qDJt8nHOdYeDqx+oJQm5kOOLAaRIcVvG5auxCuowpVzoI0ok5yYhfnhKyMGrtleH
oqaOjfIJ0WgIp7cl8eQrZcqWszMKoZdXQsf9Ts5CHMe1FVpwAnG0eaNS/H2E1uE5
jOYDn+JhGKOmjjXdZm+eRwiVMJf0+UrVma+p9Dn5n3PpEFm/rZBwO1Xll4TXiZzY
OTC1Q3423vgoqSUmw7A8UG4mk39vUNHuU0QFxqZvdFZeAXZA4cjXdyTo7Xjj3cKc
nrE34Zklc0K9IdEOm255IHd+EIJ/U5SFdipdZ4+6qRMcxG+RZEVC1CiH7xn2Njl7
VZL0+yjJz4Ypr5MTOVyyFJtRMFTRfObHD/rHZFeTreIsoevRYp1UENoFJVNbBqi8
kj1L4F9vxMAHmLxVlWNHx7VC76c5vh8bWiAdqsyNeCnB4aaLE/ccFLmrrmxJAabW
uKYUj3NJeV+LaeEMo27phu16z4GNbQCqY921nmqPAIszV54UkLfuezksFt+DLxZh
6JsAMg7dP/wfcZ2csdxmY5C2a20lXOuxKDc97nI2OOuBJKaF8u9deMmZ43LEefW4
QGok16NrsPvxKDej4eXuyTs1xuwHQF8mh9JbqUtsK5lRFyM1kqlsg7R2LrAO3r6A
wI2K6EQ9cBT+QE1GHHWKeK42DaBKqFYXpQXdrklq7V+aGvvm0/w8CjddwYdP9er2
dQbVDAePLU6UTQX8bMu+3oyFLX56axesj5jtoOXbhEN8cHRFgZrlUf0Smrq1bxrg
u4AJUM8HcEDXt8CIsL2wPGud6Cb2WnJE1rGGDI1YFjgj6HoWF1DMhF2wi3xOSXd6
OcWog6FqO7Lf6t79rGtGh1SW0lIORfAk49NM6YXd2mUyybyC+407cmuyLOXX3I+t
fX6DzPP6arPkbv7hA88DgwFo7Ylez55ksKXPVVlaP7tWvv+g5y7XSmWv7CKIs361
U9u2VmUQ/2lK9m+ENTeVc+ltWWYvWJw8Iucu7qBk6kwkRMMfYGbX5aAySjgR1Yra
1tpGF+pxduml0CS3m1H7b5zbSwv0biW8vZ1G0GqJw3cCEZsvhPNRABI/NuU1j8tb
taeFTnmikhms+J8Rdnz87a04mwcTfD/Tf+ETOpfLJhvaZo26BNk+vXkbRezuhEkl
Kpmbwn3jtXwsBokIYWO6teNmPQrIzYVcTfv3FVnezq2WjTbgjw3t/21/A12keWWb
Yg1AK1UU+ic290O1cjXDuhMWtaGSyfLLghSeG8PqHgRsO+BPYhJiMY5R7ifgm0MY
+imNpJzojgsk74OUzH/ZB907sCDXz/jdw/i8nlvQdTnE1h0PJFxeFOtaInO37Se4
EQNT3E91gDyfBjbyqKvAV+kCQVMzQGLc2uGH+zchE4Ht9Wbt0pI0JX6ooh0SZoz5
wxEXTfRY5dUI+YMtwmQo/vpxSpJMriE1jHMnVMbY2ahPo/wpUtX46XZfgHWuhHGF
/DddQ4v14i8iywJimV24k1UHC091/qY6GQwI4UNvdBcDMYX5gLGBsTXqY84BSIXh
if1ew8tOTz93n8TTk4v1A6CayVvt9ncbUExYyDIQTE03RJvWUnW83WRjqkZbxHht
4A+ppGcP+k7Hd37Z8j0BSYRCWF3uoqT4pQ0RzNDJNA/W1hPljb7Tp4E4dz8zbFzu
j5cduzdbtMvdRXht4YFw+FtdCMaVdnR3iRipA5528JYauIBon0rLE6I6KoNLNp95
fBF14TWvLAng98jTVVmTr3S16QfZ/gmUK5WR4PbW6ony5EmCCkb4KwPX9N2EpLCn
U53/Mt7DNCOQBgPO6JU7yz/5UACZtcGO0fZlHappOvFjsz6O+olifAl+5HpinCqb
e1hA9zfP1P3NDcH5wzS0z5h95terjBP973VFQTIduf78cu0haYQAerocZifasJME
mBhgw99+9R34CQScd1H39u428s/ySajjPgIplj8DjCeC/Szfx25yQejyEfUqbzWw
IKLjoYPx9DCe2o1WlqqBTOMRczgzV4G3j/ppFzxs92EfgvKPVFi+Yu0mMzSOIOTG
w4VhkcnqjusVMuCz7Gn7Oc92153HFoDh6QP+MLgLmMjrpbMIHlm5ULY3cruj3Bqf
zPYM8NjHtLbXS4nygiGJ9/jT2QI1FuWvBaEBTiNd6lVDsDBp9J5xb0drzxSxGuR/
fXbViXmed6ZqyHO14LZTpMyY3pHgt9g3lDaOhF0hIf8keAHtCIXuWmPrRFmSo8Cm
jT6xwpil70v665lyLms2tXPCTgOQZ8vtV4iNnPqyWZVg/DrX6lzPiQHxDr5bpgJK
m9NKUzWUJXYlLmMcvCcaqsBO8Xgf8fSZ3JMgHxNvTDH8XwNOsZsCLAz05XAXnC+u
4yPo1ELd5BRIdizFSWdVA6HyLpkN27ago+wOetl0ZKMisWyjFPkmetI/fOIJ8rKC
HnuLhUVfnlS1aFCdznWS1ob07PD/IyKaYb3GD21BDdPSta5jrc1/Gf3cvOl85QET
DH1yH4Qo+iIt7/RAsvy27MoSNHRhKihfNUGAatY9YyNXhk5am20P36Rtc8fAAgaG
VszO87MZ1VLWfUmOfEBrSAyg9MIBVbSxrR85+Uw71LRF6Q9j9bX3f38w7ZGrEK48
vwMAV2MU1ofbXzIGlS9uKMC7APjDE0a287S+t1q4P7xbJzwwjwFX9uTcfX75XbQU
wmP1anPG6tB4Y1PYivUptNyCliKnhE3aNPwUe80ZIFuNL9JlBgsBcgg5vQ4gMgLC
rdHMtOfDSA9Ksq1vz2gXws35X0XT0Zos86cIKwhc20ctmLavimg+RfrBDRIqumzh
rO2dC39V4Pu9u0Dw2GMkEDxEFmfOm45cOqh0gRbeOfX5QoTZUTPydcbdSi4Y1R8L
Rn2zUGoeTiHFG1QXo1GPjhdGYchb0hKJAVuBEFeIePfB/z5/fRtId8V5YoW1tWe3
MRWNJtzYYgugYKFWGxqdrouSxLbW4YHVW2Npm6uCW25CvnKgDS4/abCWdqYbswY5
rutFbApxK0bHvuYrS2oLE6VENigBbZfU6goKGtgInLJdQ4j7hHvZakSy9PNGZVXc
pBtuyKfbCd5cjYM20qdPx6TMVyji70w/m/+AlNXGPPRDVmbB/O6mAxiZGJLfa1Cq
9kCAufgWr3foKTz+gg/hpfXTD1jG9KvncrA+Tgat2CGbcv9SEHDhUqYCT2A00y5Z
blZ5/7soUWdyem3LtWiBG0wt6qdzPFFKDMltgs7wWdJF129VlU7SZlTEtsqG63rp
PwG+XpKIScxFPzvf5h7t9SvSwE9RcR3ZG7Wi70faOyCfXT7wpPaWRoOo/Tfcnt5M
tGVh8eLdU08XqF526Fixpppu2nRV02/Im6kcQOmgj8JSF1Wzi2iLAIN47Kb/vtoN
6q09L7g4xScuiMK67pEpl7l1O7btHYaLFuLRs4Ps5hvRXFA+OjShHZpSIWUlV5px
foigYBSPQVicIoIDnZureELSe8pL03q6YY/oIMdn68FR9YUwC4qmSP9++/GkiIFJ
IX8Ae0lub6WkCZKUe+jkOxmDfiRgGZga69XNrSO4tT5QsL5tOW+chtCrffnwzuEM
VnaAwNQzj+6leOoYIfC05spvDcKQCifEQfl25TUa7yGVvzhjeXTtyC6azx/WMoNG
MLsx5h+LpDVsjVuvkhOV8Y39FcTreYE00e8r6woh6XGgHFRaRKfwxkNI5bdHaRP7
MAb42HcTV+HDzFHnVXJwqpIJmJoISqee2/lBKhSzzYSyW7+lpw8SXEIgKTHgcTEW
7HycypeeijjXEUGgMqMSVoacyLxCji5xFipVxQVwQExkxH/asanelJdiOc5pCNab
y/Lcos+nosGafEJEMJW7IoQLZTCLOOZUlWUwkCVP7kuooGBrMTTYjvR8LQW+lJju
T61crBU7nm8mdJBYnz8Y7DrQTFJzUDHmAD66DBs8moxkIRjBMR2gJwkVMyrKsHHK
ygaMSdICxdJLzJ+bb50HvpH85d3JWivwFOqv4/EFEtjZmapBqbeWmIIQvFlZOPzI
IdTMfstmjfFxebaSA+Js1oDfe9a8z5gi7lRcn1GwPk/sKP8hTNYHt73fZsS6zPvZ
GzVrwrWQP74znvr1NKzTrXtRt6MZTj5zBp1TnxWpJbamfEFdyXn1xL8iPgkKxxB2
IEOIlA6CMLgzKlsSPZH/Fb8Qw4brD24gMEYfdaMeE5B4rGiZRlj9X1kNeWzkflOa
dC/MN5EFIFJcd3o4wYUNJbvNo+wjXfFtFSGzE/xQFd5CYfSn2Nj8owC50s9YB8cC
VSCOgyvSn2RvJV/w14Wxmr77JJVwKbrpZ28ajSvkkncK7QV46hLvbew+TqkmHYtN
s1uCnMoo/81EPQrMTeeb0RdHEZ8leAgRLxaD7I8A6Fmrb5sbIUYnsfEEhS4wu6DJ
UNAnru/xGbqg4b9dXV3FQJXjtV+ecq6Jbp4xE7AFEnaa6aBOKpbYz6syPwnGM9Q4
3oxWjG4bzeroP52ClxqApRzkN2ILzIbqq2WWXlvAJvj2q/TEX6obB4e1mIX/bv3V
tf3GjVxmSn/v+SiU/Jo8mp/ij6gEq46lZrAJLC/7FIIKUDk/cEmQsho1dGynlcOK
5mujjmPTPYI9nBbgf5/0TVRp2cwqVIvwoyNVBS5HiGGVfMSUV6CcYi0VCS6Autsp
rhT5HM6wRVqv8kVhbHup3IypDRSm37s0nidKiPcOhNlmOKmHgVxd2yrVM4hKzfDl
RifpccsGoQ6/w2AQQp84lxSO4OhFDtlbSD/yYZ94Z+3DupfKb4uTgkzU/he1y1nq
VSZcRAMwTfCMOmMyHm2PU9J1547VNirRWECfUtD4Gb/wkW7H5AcG5UWpFtXgXyD0
JoVBD+/ul7tE44dmyohUv+xGnzmwvyBHURt8AUI4lpunWSR4bjoK6xFeJRUyFnXz
ZhqeTrQyVe9ZpXJTrZIufKHDs49ZU8pRK+uCQYzeXThu4ijSlDFDHhioyeZgUEp4
N6hVjOkcgOeX6F7qNyvFY7ZlsoZLkKz1SOSfha90oqZOUe1WgcpRuEbCj9cLuAwQ
DWtzakc4doi9VOq60MdZQA9/uruhpevJC6xj/DBqyNoLIeg2PPFSTEdXZrzOAjJE
XbJPpr1U/WDNR859HuPEjywiXFPnT7uTtkQF5wczUq+JZ3tOWRuSCssP8257J0F1
JXXca49uCaFg5Ql2D+dvmaapoeNdqXUawXkRRmJzJltqSoIOm6tCQUEiS1ZxzX2p
PN9UZsYjo28FzwzvsXiU9I+YMDFkj+Ln956FSbw2ADxluzz3rlPfDIDbGhOvwVFx
LNXcIqd0kAjs5Blx2pJgtEa+8WXEy4QZcmGHFw/i9YlUUrHmnNURIVJJQRFaSm8J
I7LoPgk2WC7OZiT3+HxXfLcrrTFxa0i88TGE3yEfMoA9a9uZYdRvoGMYAo5D9l7l
Q4iqtpOemiEolEHYuN915gFs5EHCa+5uil9n+e+z3ygkA7iGFBbXswGOBPWO6Ugx
FOHQQ/5LMy4NeHLp1phcYwdjElupEK0NLgb1Rl56wesuhQ0ZvONW0oMBa8RjxLuH
fvQBAl6Ya5CwvkuByBlgisTEtfmSO/xNNV0IJGQvgoLHEIYMRoasB1l5AbcKZxXy
cd0BTnra2Nc/7Wt3xAdKtRSDu7qRasDd383Hae0lbCfHqKGRnnxvDGsf/4KvwgUw
ryee8al7/vsrDF5Y3Pni70tk7ty/AlJh92DXsNxs2vNG9E5J8KP0rZGhDVQ2Vs4C
oO1iiF40HTcA24jJHG3om1SeF2cZLrMYAL+z2TkCSIApyav7hahLrFSXj6M8b6T8
QgjnumKbIQvbgZUV/QtnuuelSxCl0SDQRZ8a4Ihjx3dfoDmGFJP7UxBs9tICarLK
Qfz0techrAtdnO17SJLPyZy1optTgHP4yTou3VXEVx5uoi2/+0ezYCq81oEi1jJ7
SRNd2d4pu+ZHt9yib/NA5T3rpXfvfjy6D1E89TtPZld/YMkhBjY/DhIKUTOs1UxN
xsU1APvVIbjKbn4dKSewCtXJtix1i/HSP8wqDK1gd3zPMB0N1+jI8tJB9415VocR
8lTOunHAShvXXkgzVn/z2OY9bnLKbiEi7/ag3uYrMMZj06hrcRnL4v4oowu4QB7J
tdEjFMXASsuO0XjAiuncTAc/IbaGQI6RkSZCU98Av/etN+ZADWRwUvt0sL4BMuE1
pdmy+/lLvutiaE1P1hOSmbQHJaEUoBgwMlaQ0fk/TDBHN8bnCbzSgC/YpWk9CvbJ
Cth9pkLaCrPfvA9++0PEe+EpVVmD9pYIWjfRjSeW4A/QlF7RjxG+weFTlMFxPojl
C7A+R6LF8dvbp3vN9Ptb4n54b7LBpyYr6T1YOQZdSAV76aZ831EU46XnxFknmlGY
twCgV37LlAeR1igFjuRcg/5O32FkYMr8y9whbsQS7B9acodDcx+frV5FVFxV7wfY
xQu3DQrCTqrjbP2I6S5TfitqGadbnCUq3s7qqZZ3VB4HPdqyRLDFCgoK7YSf3hn/
psQ+VE3KgDysrQ/qnmULwOajNuQCdYKKIDcIrJ7yBxaIeu7nm3VTLbP1zLPL2vt5
b0DUPrd/POV4Z40oDpC8BjTlCowFYO5Uw7ssm1DW+J1UsarFR8iV1dU1w4vWbmLt
W5fn4A9njqu0y7S2zVGa0OxEYA7nZLLS2jbfadGAcSd5RXXI4tZ+19r2JFEIt7Wd
34yv7u+U7rOjY40yRffc5K3xfv0ab7I7Hi28Kyj7JKyFOX+Zxh2tVs23oKqWQYN/
UV/K7MrJy0LgXlqHMZ8A6LQzs2SmGnPueY078jtSLr/KbGvaqgku19mktoLyQqBE
HV0KWXkEqNHMERAc1A3mHdNDk7M61QeLFK5xHpM6AjUlwuWctkzeeBihzIxWCyIc
cKynyBUVDOSzri3nlkbI/R/bpBvMNz79wLrnoNS/EOe6Tp4p/nHwytErh5S8T+7k
a4rZGyPwfIMlabmPU7m3dn5SEu+F041DezoVotlmVX2agUhZL9tkSCrE0ig2d23X
XmhamlGudKnYfpHRaJ19N/T1g4zOaOryQExQa4hxCiZF2yOzc1Q8Dbcku3de5svD
n/z0iuQkKA/0SLXhHer15WhvEDFBJkvzY7TZK3azwlJiixbl4GQXOmgiz7FJSII/
Ffhm6ZwbJcfbhVdgY0fqZPb8+FyF2SnC0HhgE+C0qiGxhToOXVFwY/wJ2/SlGLo2
5db3m5SUPPX24nE6srehJQKxcPRoGZJRZyXal++BA23pzER0ZKT9JOt0LvGkIeXy
CxmvNpUsQRh9r8OWkap7T4B8p4xXuSl2P800kyaaciTknYX57SX3xV+Jcgwa8zWU
C/VZZQWFYglaqu01ds4EwrOxevw/KzeqQBwgP7bqjh1elZtE6C1uxBPFfg7HDXfO
6GxozPRvqI0Xwxw2cpdUE4I9A4Qa/UEcLeWAiaFYiYjJJsPG4D1LWqS5adAEkHCH
BB5nVgRV17RrwugwOpmlUFJ070SNDf59yoF7JRgfh2GA9wEgisThKNhXlOajAgn6
EFbpf1NJAivOBWVvIFCpWKIXcTXDvQ+Lz4drXCIXvhsdGyOWB1crxpB25K9CiCCT
PYTJVJiIC8nveP6Lb+gP3P9yoEy2Xr9g7L4UlknknSKcAm+IPUP0xvbk6Xs9PHct
Aa3fOq0IL/CCv3/QOc1TCTNuTOLQ5AVKx6I1TVzg9PIfKdHQDIJj0B+5U+AfJks2
0Mas/duY4pBzQKXzCpJ/xMv8X/igQW1P25GeEMDGd0cpmAZACy2NxFxwF2mCETqT
lrpy/CgEoQL+1cfQZI+9bo0OySX+HsU1npnut4L5H4/8WTqG5YDZHRQ6tbqFEmS/
QuMdBrSyb1hOmtcd3tncM2HnNFWIqTzPCcFGmfK6yjfu9vy/9kiEkEHOZqpiiFcJ
1jyV8gQoUoMuHiBa2aREjfGuw3XC7+yEx45tgR+4O2MzIekhU1q4MgjJGCuHK2Ze
Drp7uinIDjudJ81ATxWfwOn5tR5mlVL43p0XwsDz0rXGxewXrX2dbwMFNtMLP+bK
OaCdoGMb5pnTYhVDWFT6vnTTeFjhEhmWQp4jU59VXU+fQpk+sQ+puH0HRwy6hnYo
qSyViCnLqoAU/3Cos5ce/ZcLIjns8VjkpsHJYoJKtCUNkDTM35sBH4Sct5nXyCkL
DitypNJIFePTYexGueO+WOeGnj6RjsDVZWsFekjqKrJCH2DAJPSNB0dX3iprHiD1
tinZuTdBOnrTY4S4mCuCPjz+cPTqNQbqiTUJzkq4wE4qBimlZPIJt8ZS6onneGPS
FBtjHrd5bGQ/k9zaCCc119yc6NY+5eQPgqO42sa3WWcTtP7GpMCCugC+pQETiuoI
pohe1BCl6WZ4w1l9MI72F88Qvth784AMQgQxJepOgfvia/H1ZfKkq1FsrZqCBZBT
snTD/avuD8T8LISKT0F74y+rxSP3knxG243fYfdTrpQlsp+N84qod6tLWCaDIbp3
5VTiLox5CZ5MNv0M/TGWOQUYbk539C4xUtrXRhNubozYBb+o363JM/S8rXen2lf9
D5Cfse1X3uHMDqsiS9qZU6tNTYWGmgpTBx76qaZ8fsCX067nr74UlGr1XS5jaN95
3km2szaErb/mWsTytid39xUr1R6wqxxr+EKQu4uTRGtwZJONFXzR15j5dBP6zLS2
AoDqvUojBKpGTzPM2RR8JuVciuT9mVfPpv23J03xFiV+Fx4cfQD05sQnfs6UakMv
qhR9NY36YeAYgdKgo7td3BeeaL9qCxzJhK4Cqb9ZpJM6VyPVpCkFKW/sVqtCdlVJ
HzPxCTdrsclIFHHZY1xv8RQKUf6PbgYpMlP8HjUrdSIbH1X+HTVxzRS7EAzqz6vt
by4sS2mbrSdZpIugW6SW+CWMmoqK0ShnJi6cMBkD00hGZqwrcRRyu3cuPDlbS1zZ
ER982e27lC+eAwsRKDFgUxVRtc9ebWrgn47hvg7bgC1/lKZMt05MoGshFR91vAmK
2/5Efa0QVcKmnngc0sJJmxfeqPAVTzB9pG+OusUe5nCKU5S133x44Amsx09VF86Z
u9aQfjWlhdqGulQyCR2Pe73ysrA+bUsspYZwkdDl0nbJe1C+EcGssiMiKCDRq5vj
Cz4+UEBeFYQAS+G/7NrrDl/GmkcyCIfDD2omXfT2Qx4sWFw9PQCnbmMIyXUOW7s5
XhanBIZ4ZA/fDGcrkbDmGkBGB0zAdtp3axQLhxX81JcqwZC0zfYH3uqiuL3zj2NW
1tMkHkouLZ1YLDdhKwY+jHEQxJOL1Nm0RcugyLewDoirtI3IX/Q6OL8LB1/4OiMG
yzaqdiX3g9HY2Mxyo599GuX/P/vrHqmF5mDdYORcwS7l7UzOpyzYDfFuDSuWQCSh
OFibxfayt4z0DU871vS7phv7rpg/cSH9P2H29ckhQNgB8h5hPbUriqE950G3/GkX
2hNnlf5e/Co+1ev9fC8kao/UkYTqY4eNzjVcpsK2T19EsShJquOT30uDuWcPt/Ee
eIdSQ9o9tKw4yfFeTwBqnawJeXv666bBLWHC7ZAXp0VlASEcWXgyjPelx2JqKC/v
9QeGeNi/HsJJz2v1CVZ9/qay9lqChuajoqwEk24lnAmlyJz5Vc7vAhUUMCRgjv/E
eG/tC6uevBh5huu/p97E3ZcK4PMPCmpuwqMB1/yoMmCVAaqJvKlQQTK2P5OmlwYT
+wmijvHLJmphPuVGslQkK1HmuwF1nMlJt3Lcbwb7FMoWf+pE/wYp+atIZTi2ZLAi
Ie7Fki2T4Jp60z5ZkCuJ3ZXwu9OAXJPSpbyl/qdfibSQOnbEN8arlt00LPY7iDRk
pYOQPKz1xEXtHSX0rUp/azv5z+X1ruAJ7rpcIPhAs6uMCwLkki1SRMcKbV1LOPNs
GQ8yCl0fWGzAYtQyPCmOhythIfdueDQWlLccDxou/QM5q4AfYynqHKxbp+/lAaKo
JaUdiccIS5AcErvAzIMacz144sKUFZ1SDc1PCt6bNFfnROZhtUa0f/TG8vC7PFJy
l6FsCF6YL9RnZkqw9H6T7M0wovS8aBIyIDfgDI7HididYhOU1GSfL+c9IAIXA+Fd
736ReGK9Au8N5eduFOQ8jhSDOzJKO3Ojj8Qnv9WfjpyHf2daEXbQhKd2k7cAiozx
QfUhr9eSpu8ZDNBz//dHT0i8XPjRyEoDYcQQf9Jo5PSRIwNKU/Ws6hJ3ITHdWx6T
fQgu1hgqHlyR3hDMtv8bpH1sKrjSaBF3nzcdWga0T3926bDsImfGSvq0JTi9MzLh
Z9oKjmCMKFEbe12WYnlnOoyk2mjiFm/fJDCdEo24lQaW54/G9+3uKGWTcqoa7eqF
dOpTucu8yWYPsseQRyzf5JxTJTgkpCpSapH8LdbSzNZzEb9haax4a9qfFzERFSzF
4m38G1t4CJmBZ4Yx0Z3EnHSYRdiWLihiJ9mfgOqU8oNhb+XRU7QEsHRrmXSPfUWv
Qun2f4ah67vAy3e8oRz7YHSGTgQbuuMmoLQhFa0LA39/wHW0xa9C2SHgN78+WgCh
9hntmRWKbRnoZHmxI55SSHt0vl/P8st7pEZPid2DxMxVP3+rFrL52NjUiNwKBu5z
+aiH1NSLwPA+BIc+Y/twXnFUMbygydhHTx24fIkGgg2TnxLUKwXRIHyaasvu8a8k
Ea0Tfg9Vp0nLo4qzaC1pf/Z6fzDc+VQN/+S3tZy8OiEx3bkLfJJEDdPgycqiVPZY
MDEZpz2VbQ2QOpmX1rx86J95ge3j8PAN1Mm8Iwpp02i6Z1Qzc4OHZOhbk13vKAlZ
hwo5+oYVdtbwaxFo7GzQBu1+oEb/D1q4dJP/ZFJVyrtj96QH5PxIi16Rzmk6UxDw
2WL32ps2NqGe7Ks0MNKADUoddf2w2yIEMm5AiPbPvSa7Z6OVMQLbRCFbCyyWwROl
XfMiDHviVBI8TDXDYLHP8+hCKYa4XdNuBDP9C3v0s0txc+PU1JQYYDqffMpyYK8Z
/pBaVDujyYQFnOh6hA+d/eOy1UrsYtPZwDOAZ7aZTT8Qa4RgS6VWA2C9GEXTJKYD
kwJSwUYnavq4A07WxSCHeyoN96PoE094xr7OA7jrL8VaE4jbwUBbKB2sqztcAO4p
swu7OEJYsgnKIBHmu7upG5tQer6uscmeRezhvzB6CDEdbzwf2L5A7ziaKuzTM34Y
nJ3cOp58XjjPQZwxKVMI6oPpAozFjde4hCvevOi+73vKOA+nvEnRvWKJd4a8a9uV
m5NblXWx77/qYIl2bK1NmJrGN92rblQ54XSBp8t4jFGuP20mA4LMafmgA44qaHcD
Gr6czZ+vMzfXBEmg52hZeF6eTLEr0IvN7zLtnr4CO1eFgh5y+KzD5vAGYMggu60T
B4lRTo/7u7U/NWu9mbvyhTbimPJjVyidlxCgVQx3EtSxRCqUWrUcms7xuWXrklBv
bovavd3ZZvsvWLkm1UxAuxO8+2JOUf4mh+xs2QxOcJcmastR4O2cb3GbUblxuBpN
lzbc47nDSBIqrLM0WUEFJOCH9uFovMNJcucZQ2UX4efJW/ZEiDYSZNMygRk+grqf
NVtzbFJ4Y4ZPnQ49lyg3HhRMUjIbZaKqYJGzvmUy8lZ7q7Qnbuecb9I5Pl7rYu2K
QkGglVOt2t3WJsCZ13sSjWeQHoXN01R6TmbIG71OgDHSDgBVCoGsgTi2R/li0qkl
l37BQRT/KI82DRyMGsCwzcmx3tRf5GuH38aLazE7UxSaP4uKYAOr5re69UKWEJon
W1jHaJr7BIPaixeQoc0E0O9buodZTvrIDMxrnlOf/pFnEBPcaa5SzzFKHd4joNmE
qWJnSspIXdx4eQ89y6AElCUpd8gJuFhzz4DYFVmDS3oCPtDdv61OScTABB7s8/bK
kKc9B1lf99v9qmQr7ytekJKVtgtAXXQr9HFKtHQG8NFU0p6cld+EsmEAIvUwUH6T
DbohjsCxnOms/U/VuHK3y+9eTgNSJ4q6P8kTllTr4ggf2ox20Wy8p8EogXori5jZ
/MeObwkt3em2I98WwGoVRX1Aga6MzDIQwJbHaHzM8VmeZm0rqrwCfws2fYFheNnO
0rT472b7M7teR2JRVwyq0EhgIgDcQ8kuliVuDYjidW7peyCsrnPs9XwkoEHfymyL
evgGFSZG1RPFCxhANg8/s5/oLYHFzAdzNsWePleoYCAjoNLNPBubkHFKbLB5Cfal
oUCPZdtWbA2JrSCA40wyicFsf6GJQPwgFMs8AnvBpx2FsgFNxp8Q4rBhkljOkza6
DHzCNSzlsr2tiEsNd1Ht+ber0NFmqiTWf3ZhrAV733FKqj3+pNCaKj2ul3ZPRtPe
hTy920I1zKHfLIj/few3OevkTU7utp7507nS8ZBBFSAlJFOgCNCSdmP4rJE+iGOZ
wfMH5mfw1afkTU8pjobQY3XLm64bGayxTFlZJFg0iWcTS8Z/r+hVfPtVhtFUBXMd
qM4CZRXQ0skq+Hvm/cJm4w7hn5AaSivIGtRRfhWmQy6EYZ0i+hb71QWwrt5hGFq0
2TEDM+RvIsw+QLwTgr2D69B5HS1zGx5/nsVHuIDQg41ovlMidzJw9SK4N8GaY7Fp
9Dgx4+Unbbg+f+1KkoPvIGKaCym1hGFaXiKrZqZ/Kmfsorb8FPAPPGFlHWN0u5It
lupux4w/kg7K3B8tH5y6xnoOtaUdvPuH26Ls3bMlGMa8Qwon0jfw+yBR+4LbTbht
P3QIEhTJdaAjKuaTxpvEFRdVdoqy+dEFY5JeNxHI49xCiaQ2vuaS3Z5dog0SLxOx
Mh7vX7nrMyZvvD/7rQu3jG1wURuKuSmlQFnVZ9+FbwG7CzzlJHHbnIr/EC1zH8le
PIvsJgqDwXtsDWhMBeaUu4rrf1kvyVTT8Vlx75MvpMbBQftAMHt6YJKOphYcPBE/
LOz1lsixqnsO/id4lAr5DB3trArDyxHK077495gHncqDwp6A53FX1WtynrfWYx3R
Ogfgt1fywGRTdN40rLYwo2RZeij/AR+Ygs9fMSO7E9NHERTZA/m/CiQmDn4xRvs1
SrsLGMIv/scjT5h9IGZ9gvFUYvMjiU90hbUZwDjaa529qSoJm0TsM2+YgMBuKkCp
Uv9Ca429QLbrv/JPYIHVcErpaykR8fuwJ2rsYyQj2q3oMTYQt5AGEkf9ukwvQhZ4
erEETHEAaO4Wu6byuKjzPEM4ibLvcZsFtL5cEqdCyjF24+oCu8fRaLupdkDg+YI7
o4ni3b70wwNaPrEzj3kGCxqtxlP3o2ON7nU3Y4yIUJ6zXnrqLjKiGClRfcZjM7+k
eetU5MlwyEnSjP2+DlzhhLbwlNytYGGgsv2gO5eFvRA4aYLByQFP6NXTmhJ4rkei
hYxQHFMz+AKrCogsOUdCVPgkj9U2cV1e5RLUBJhVVzzVYPcimX8AKoUwAIhLMC7T
hlgxILxfGEe5QLd795TpN9xXjNKCp0MWSple6RWN1G/JSJMWyoDn04AmMWRssgkE
/cuLrFfpElIpaiO1hcjD5r634+XoudKyhZz+dQfikaSg+T1QF8PfzOVS4BESoy6q
z7jIONRIBYPvwYT7l2VJo0omiQZ71iK6ZKWHbuRtwMNljPV+69wAPmASq6Yem06l
R6sqCMdyN35GoAqj82EW4Qa9u15ibvUUAoIQ+bOusPkytn0f/rDC85LzV1KjCuxZ
zfGmzLxRAsmnF/rMvXH5bNxDQ0xCvbiyvCtIS5iXzmcD6bCVNiOrWb81KyE8uQzR
YfXZg6684EA+c89NEA7MvAgM1c/iROiBcOIfMPhlNtCppmMcz3Lq4xnbQnEk7+UK
3pynIOXXcthfZv6SaHxpZNjcUZGhTlznEsCAtnc3+ac5ptZukSmsyz9qrxUUIpf1
uYVwOLWTj01CsZxrxdY59CG0i3dFR3DxIWjDK33YVU8BaIP+YQdcPfl/8DK83SCM
MhtzFYVF2HLI9oyoGpT+BglNOVOsGd2TYa7tkG7b279OkGwsg+jacgVHFWEJECnh
d7oQr6JYZUHXs7srO3tlKa8L0GTU4tRx6fGcBJMqkVjhErqKQp9Vqq2Y2ysEXwX4
7w3TkgUB670e5PJx0TGJcw099E9SF3IaFp7tdEyvBDi1hz/NNaqs/21EaM+tDKLK
ysDHmu0ZeDVgr9afr+iKS3n18zwFIARBwsW0NBbX7A9sNuo3bMw94O1NDZcRtJpE
FH2ygE8YjQEPaGvAWXbCLykPEyqmB/55MgJbnf8ja6rHl6SaLdg+wqJqjGlVtNEI
tosqBCo/b+wo8S7+I8y/vPydndIXHEQH7ERPAVoj4RXevomi57ISSAUB7LovIR9j
GgSqisC7CXvDpmlBc3pREzWEW/HPpF//ME8Q5lkbjwOhQqge0Sfl2Ni1ZZk3fjeH
Lo/p6GFdYVqAEIU7gGPmuEGEzUghEgOXPMPRN3iffKRkAYwqtVnA6Ndil10hV9qw
LMGHZmZ0VASJoiMmmSTvNqAfZzXN7I88rb5WTkkp0wMvWmOy3raWuzyC8KQW/V+v
zDBQJzgcILd67f8mAAicHRI7kd97l8vlM4a8724/Zvyno7Gfrp9B9DUKTk86EZ4Z
/Mg2zajwJ/SnPMAHyj0dwZoEiLB+wzKB+tseFfs6Sx9c8mvQFz03n6rCzQPH2Hxo
bnKymgBlNVXK/GuARSpUlMLColsNdxclh2qHvRLT6S1t8ggxAWx7CAQB3JveG4jJ
OE9wM0NG3OLj9e+lQpGpDvpBkLNgPAB+XttLDkkRhK/1+QHc3KbPMiZ1AA0TGgMq
RDdu7getY0hXAZq0StiGrjybMdFpHN5tL6UNPVjORB3nlEP1KS+H/kaBc6PMjmoO
JtSh4GoWLQSTMZeiqqXiJucoFd1EK6wWrtRl016bXiXVg5/YvkI7iWBtq8n8pawU
kyrL7Q62YdIREhcewuoYVPPy14XvGLJOlKnUtU366DInRF0shNpJX0XoWrmZ3Sjs
XGTHJO+wSglslRAi0wPOd/2b/ZZ7JQgUcEzVLvEHl6BQhJBfgRPnpBaIjBZRNuY4
hsM+JXXmqodAVh5vAt53D6WCzBiqguHHD9u4aTcva32UGVb6z2DS+TYXo26NAmzX
SmYqzzPDDWKKaJ+o1p+YSFPSWzIP7U2TlD3fseWkRecWGNgIq02LxQt83aRmTEkg
UgIoNc9wpQhSExDFE0+a30qsC+Rz48qcjpLSVJEluOW57G6aMEPAs3JMQjRVICHq
kNOwCgugRObPgjRd/UOd3o6Xjg5E5BTMKdeakNi7XG71ggkygfsDcI1txOtjqlPY
vdLIzysMgedBHRPwFtjNvjxxku2JrRj0DrjMLpOZLg/G2WCUanH9DlpM4OP9Bm5G
+o4QE7b6fteskQyidC1oD7FnLy37z8d2Hz6TdpAnIbHubqV+KrTfnkqvt272xFvl
gEEykjjMM6FiSEaNpNbieG7WwVBrQSUgm6y0O3qnG1VCuN8vzSNzLRXbFFlh6CKJ
5n58qEOM3VlNgZFtSWqMj2KVaJWttQwXkcVjIGVbBclBMFE9fsHLBwbT6IQ/94k3
XfAF91GAQtEAJjAyiLPZcIJD5FUGYP6YOAEP1xUOelyiI9uNEacMJCyQibIKGCyP
PSuK7GQZEC4FeEhZdvD3BG2IegqEyOXMqw4JgQrCTwCTcL3dVKTpUNQpKztDOX7a
G7UeUEIx41ocdXNJ3gkSGm2mw0U0+jm10HjIosm/VYtK+H7/BdhkAS5Cu9HNfF/j
5MflxOvGpiPCN4kUDaXoz6EFGsfS6LnrSsmj4+gQgJrTa6zzQ+KNlUtQ87MXIbis
jq6OiXP9b3VORznX6W2BvTCJeutf2DscfxHg2MmqLstoU7s2E0dwB3B48NcvNfdl
7u/aQzeTf81EvIRCzFgWw6wLnBP8/+T5FRePw+FfWRfe6/dLrA6OkJDmM63JcUaU
9NfpQZSi7gsL94sTX8vIwYf1/xwW/oRf25FnkeaWNaMTAh6whUYDwxJVTrgpXjzF
bQYjk0w5hG0Y1tZnrOK4PNqKTlOIXhK9AKD2BrFLarDoF2Lgf3P4vBzsKusR0Wg7
qUbi/8oMJan43dQBCAImdeyQoMxxee3280wca8HHbpCgk+zf+E/wqPBupfMH74C1
RcUmBN2gunSiX2jWaDxyboOwr8OD4yhcVLtEZ/NQPlySHmSANmuOnQzTMBbYkdCE
uiEG3Sz9nyOhW1bV1jKkXLH/14xPjxdltU9V0iE2edaqkjHpjqDVAOzvNbXbLFn6
+LUpoFlKvOmT2aeLQLj7sTxzDSyueLWMx8bGu7y2WVAUhQ4uGRqjcG6U3xJYAeCg
rjrwhTWzJt6Y4YcKERqhzS5aZZbIM/E3rxMgIMRYk+3vc+ivYNWrZt/1ebrBm1YS
pvO9DpSIVHyLEb50YAduJ1q0BnG3PXyMZUgwK6tBIdMfPDhy7Xi+z3I16iNB5Mbz
absC9to+YWDEjPLJ2sP8cC2JyUd8Ua9htUv/NR/mhqOXwZYkU+24DKKe2pUIp4Bs
dSygBo6Z1oMprFZRdY2hyVXP9tVI5E9O/S6wMdywO+PiApCkaHoV2s7J9SiBM9c3
j2tjMyrWiAeg6jYNwIOSftOliqMRl7C7pjHxQtAbcQDuIzZMu8fvpQ7lnZw3ICpo
IAhID1fIYaaXARguybqUvD9dRg/VLn93ueJn13n9rTMB8xCUVX3aGT/7IRxXOrKI
p8+7IidPr+RipFY2D+8jwPBOdy28IY+NzVzeMBD28Ev7wFC3uUhOJQYuY3yWTHZi
NaQFeQEhokfcbjs7k4g3upTKHxC49oYJMRSQAbLMzq96kg6JUEcaNkwsn9yFZW45
TC0ECZrQDqqSuoHG+WIziXlJT3IKzh6//utJffMqJwf0SGK5dFRclJgSJcDSj1eL
JnI1sd33YZNh6ETJ9lt/s9soGxR3qwwvjFfi07oVgKqsuKQaF9LxMIufs0aAT8PB
xJxNoqTZeSiCVYTUoHucyrazZ23iihIFMtN2eU3473a23sbOF8cp9IKp6tOXbti4
eOmdW9q5JyzYBnwzLn93IisSxlQnSQL6nnJkrOmUL0RFjbBwISK4dQJqyTxZwXV0
IsNgV3M6RHj+YMrjYNSa89utwkhtsbJLx/UMAh7Cdaq40OUaj7YP5p+ThBXRaU9X
/fHt23opTa1A+5T7Wy5+fUIrVlazPjLmWyYMoYZKVjxnIcqYUbUdl/2A3WyZAehH
lCtTB45l6gNwbDAj5NJRhAYZF2w+8q7e7diUlqLoUVivcKYeWyfWkqhNoYv7GmRd
SFMnRnCBd6iQamqvx6xgjh2OyArSOiCFBjUWf7fvm2xdpRJ51DvSEc8xaflalpXp
r4JomU2JlIiIcwp40YxvqSIZ8YntKBRjlqa3f+dZgOFc6oV1uetSZW26gYWUfBWM
mBeWCqF28/pALAGWXWYywMP7p7Iei5CYB4I+wKP17Zue6C6QwafKkWTfiCqlpKRf
rNXxPQ15/dtQNPJd3T65WXLQORJlAbI5lNXU32i1uhrl+5VZ+EWgE3fs5BKfBCLE
rsCZ0NDcDXYc6DbYsiGYUjjdzsvRsPYmU2HYDTG+ilL+ppQsE/kgVK04TpigHosK
by7wdFZBFtcEStfchX6ji+vz1vBqbU56x2XtqV+lv9cCQayHTJ/x7DIi2qVn901E
Zl8aQnDKvX+YcnwwrWlh9XZX98QrGsU5ypiNgxxEsMmwh38z57Wc0xymvP/bm4gc
b+M5sd24keBTfPoJ42t88AmoGXVfC0WO533PMxHLmbD69FvsP3rG1DAdKCvI95pf
k+bPufN0XChfl5FgvibCxSNzBRoWA1NsweWcSfYKjIJWXIqoRHy/65IEQAYPSAIh
t6lfymJqnvaGsBzyVkTL7p2kY8BT8xG+jiUy9UQoh/SNq35qMNE7k2cRttHBBtId
5cjXc/8DvR689wPvkUPi+Q/rfllRLSoQetN8SUOWdpbviPfA4uMWgs2gQuWH9IGW
MnhKbG0qKFAm2EgGbc/2X2SBlc0e+UyPwz/16r9Fq1R9lxaqqiQmxUqXwWYjLq6z
9LSZXzhiGEDj/Cy1A6QodiavrC3Qq/Sn0dd6AgF3e6YXWx6cO5SUPY2Q7ctI8wOx
2qxSBdN5PdTYbUhpIGJF8C7i8aU1+OTDZ+LH8YZJkKB1W/hlWvSVPQ2yjiXSMyeU
Ulkln+c8Id5vni+1yyFS5HUQpEVUnLVR32W5rvCrvMARgsBvnzUo75EWyHV/GV9S
TorytbWfxvtEO3MPvTP0cEJ1RJ0r6WuM9elLb9dA9lp1m2SEB1/LX+w/llMBLPXT
rIBqspX4audYFxE9XrEYWeEz7GR4TVNcs3quBVkhaQ2TbUuLGThF47wJWF7i2nOf
ymvRntSeVNAT/58uK9dlGJAg1JbrvxxnNqMB6wtG+WDq9rg1i2ulxURg2eDQSkfR
pPytVM74wmdiomNMDv4FYxhdK3ZZrJPBjgCo7dNIPp+lX6uwctuMBZBy840Vchsh
9RQPeeN57B9+HLkkd1xBxEFjD+rDF37yY4zNe42xMnCizZZLe/oOyhFLwOGUhF2i
dNxCZDMOihu/x1DAv0oEoNgER1E9ZWc+s61HGMT+atyRv+shzoxyR348zuK5H+fM
lGRfF/mqwQuBDfUcklcxZijvFD2yW9w4l3XD/h9BnYxDf3SmR20DSWh8Y+7VDUJ/
R2FPMuRaW5lWMQCgwg3ZlrkRUtIT8gLw/XpfjcBDnawaSLRVptIKfqCoDSmja2r2
0rgtWiRvBO1R/HZLMiEdopSmkIP0g1uup1CH40d6NNpHwt5f5rdzGewRqP0WQuee
/7hatYFOnPmOMLEke+7N7egQdnNJC9oQpcaHOybQMK9xgANbwaUuJQfNnxokkXc7
fz+AOLSr5n62hYxjXBfZZLhmTnYUsts3Uf6yPwSfA7UljdoASbgIp5ijzsNsCwZj
fvi9JZGm/zFbtRxp2IG2o+4KSTD703izIBwl8p7EoT4gwm6SV5yj1ocDbi/jNdN1
zGtdxz61TcchgW/vzppK090i3Gln6rEsnEFO1WcBbTpjWCBBIaj3kjQR+YbvgWYO
Dlu7CS/+peWhenJoeMcRzBhvOrdxqoIA48qX+8CpLbDzOw3dP10PAL5FxHWphZCM
p8XFEuiHrEoKVGzsnlxoKqu4AJqjQrR6CpbBd9ck+Htwce8U74mfyEqqifztGMep
lwN8XYjIkMRT7yv65BROFvV6bygGIiMoONXnVYPzGchYNx//Lzhickk9/AI7HG/g
5Vw8DHVrnQz0/MUtLWKDEpNwSkpFbflPKwGAjddPpvTp/HbXKD/eEFSQWb3CNhAB
1dqb5L/TGOEzIbL3mUDL+Xvu5+xDwlj6ueA3n2oCjuLuZN83DLRm07e5et/FVZv0
EweM5E9Npinw0ZuYoaaNy3tbimuUD8P0K/40N+BrQ3b56wAF9quSIvtG5XZpF6og
kXd70qE//o+tfOzCNHCSJpVu53dc42kPd81xRRNGSjuABk2TqDas2jmWcnlbNz4q
Frk8ScBc0bix8QnAIv0Z8eWktmJeo3dctD7xpmkgF33586wfgyfgty+FlmUPUAa1
+3MjQDCd1GIObJkwGDvWS+NnjjHxNFUJT/34Y6pbUWrBIfRvxfndYVtKwJFaWXhI
CBzt/MKGMe/5la9o5MiodW3PXMtX5xVclF+vLLz6NoEZopeT+G82CNjeYnCrxTcD
gVWm87Cr9FUa2Z1V3y6QFhT3q9wpPHzrmCcreX0ucct1eivdLp1St07iNKzedtjV
j0oK4SQr7OpVrMc5SxP0WfNn3T8JJmUUGAkBXx1VHYo8Kx3Qc7d5V6Dlbkc99H1H
zkrwdJZM5gAFU16KnLhKgswXCBpwYo5e0aGXK6ypnhl3qxVYNFovALQuMHWJCdEq
cVnDt6/NZ77pDj7GVyboNQA6HdcCJVfRty9IwtoyFbfVr++iNV0zPj2cdM+nWgPj
KBLwPgZ7W6HAkU7ZRtle2QSwzxTCZ+OnqcjN7I74g7VFfPQw0lHg4qlbCVkT6H/n
Xdq7GhJ8BdrVWzfm0b1YSgv7CGQ3kB1EEyqbJR3AD6Pkbgc1sdyQIDLaxWYDTocM
wIszSZrXWz7FFkg0um8QZ//3uUmC7TUWjN5vUndwk3+4wqjg67u5HQbwcmfXRlg9
vWlKIScwXvpCGn6zykcnqHCX5XlEOqjb2T2aHaE7mLCV1AHAriQdw7HHWyOE8qH6
l5284H/uZ0Hex7LPpY7tuQddgSi9SfNbeljTwcTTz9JdMHIMi7LuoNZEARrv0xw0
rXsb3q3ipAuiaveaP+7ewu2dIly8Ip++tSVyTIHAcZzqQ33baZIX9EAPfK+8PnjK
qZByp0j2//Ftc/qIQHhjugxPn3iNd9zqncirUBPM5P9HMRAIxCk6Er9nOC/YqnaT
7rIoXZV37XQ/baOCs9G6pQojLmXF40Ri5F7upJV4YSSehW1iHe95SHkcTQbuJBpJ
HGVOziapv/0bxBKqSv1hSwvtF9YFzF3vIYVofUecAlHHVT0Q+kZcGn6Owe+ysNyY
9citB45srU/W09Rdjr9cNefiA2tf45YXEKtm7CPME+LEeWXcprGkwy+deaj2eJus
xJoyW5yJbIGJ59yM1kHIZxt5596/KQ8aWsoQ/cQjZfdUBT/mPTTy3a+NoNt8ziAc
aXzIiDPzoNQLpy/8CnHFOc4e86+Dqk9DVzw/GHmvqLcekxYyYgRng0kJjLS4yOcH
41dR608SqxC/3zRHPbqgTziwff7xNStcHaBrexudjEeUzWW9K5aLl2sNxTnSRaI2
20gxYduIPt9VjTcDDo6FaWt18SgknOeJmIeu7KXWIZtrE9vC1VGVsWZnvJ8ZgY/6
YNa19XnEL/ZwbyrafOCA0P/vXd6t/qTv3LlSoY6ElNWXVq9g8Z//jEN+lwg3/AFg
sbAVF8VNE1Il1fbUwcUvJ7gExLbFXTzyuNnOshfs7dFt4IT4qScXbnSNHQcTVmhe
jfDvYM6TRVHam0q9MvcWXKPDMazESC3yTb9b/trs+YzjacMXCVdzrgatSxK9rbsn
F5Duq2tNxDpVWE9S83QsZEV9N/2Iyb+mB8V37YSM75hKiIgYtk3TCFp9ouG4Dsi0
SXC/fmBHiWXxP7EiI5RmjqSUvP5mDjCElPjv37q2c4wLM44Kyy+YrwIY5XeVzi7r
H2hezapCF0dc55r3BFCUk0yLmDth+i6OvYq8B0XUArEBCaQ8yNDIQcr6c8tqFRz3
BmpnY1wOIXsO9ZrXj5sTeYTfTMSWzStAl4hlEmZAWP5HD/v9qmjzpuTCM+kz2U35
Vtv+X2RoNAP/OwNlx84mP9SuUccz1qCniozlzwnXHopz5EJsdO797K0iY9T5euHx
nR3/yH85QB5US0t8E21VUeJ3bLlgTbrfQLOYuwQEbuRaRrvvs27n2SdC329ojw1K
BMorGX+/uWpvv4zS7ia68qwlnrxlsghTrBYL8rOwgzD5D6/qqa7aiGc6OtBa5uDf
shcW6LcHU4LF8KO8H1IjFCX9qVCPMXqJ/egw18SHpmwIYDpAA2ZoLhW9dOQ5NuOZ
j4xxKxY9vhRzwnypLhTJkFfFJ6ZHXdKq6Z9PdVUCSzV3I2U1ddXR/vFo4szjOpqO
IzI8t8GHEvnMMsYd4CnBLcsQnCTKteoYQvt7sNhnnFRbV/q6eNjGXAuSzDp3Eu8r
gh5toRyBkOOJoZP2v1mXFRT2N/EKsAGifT6bMkMKKwLPjxTUwQHaIZkJ8hSuXpFC
qU/DOYcori+HtsLqULDVgTCmRu0S7BkP8jKaMGPaHSmTo7TRhIEH0i3yxCq2JBEv
zqiIp7RX1aqxOfM0Ni2B008Ks6VmE7vFyrKMd6eTm3Ft1zT27ANtIQxZ39pG0+Ax
s9zbEtdH41yNTHGLvsRmmsU8xLiN91Ps/j2f4UXiKUG7z+NbzY3Ohjt/9t1DVnQG
nRALHiDY0kIlbclEeZJQTFB/SBMfbuORDaxd0yM1XZAfW0xHSrOLCM8yO/tO2AMm
0CQAe9g/HZCW18SaLV1C81rvqUyEgjwpEhglfUx6NK3FKhhZiI+xeulp2O3IW9d3
BM1HtQWYJ1UXI5OdyvVYqlye+vybJazsYUPHWgaGxyrZt7HJvB3lXdoTxxlDnxjw
BExVMcdghXK7hMNDzUEOns0PhJnXT8J9juLI2qgJw2eDder/e+IiRGfX13bN+TyB
9HO+c3isUCRJnQltLdy7htbjNdWCddYpcoPtX4af4KLb60h6jQrub8SkxjqWj5MC
cRKWv8v1RBt+V4bqbIENvgaUXY9EpOKew6RwKGfWL/UVJIGDP8zPiljt4oXGoDjl
8lfbDZptlNT8Pm0I2tufJxIpiH+s7niJjAjqTjxqSbTcXZfoPgXWhouyLXHqmkuv
Nv/oKPZzW9XakAQywxFl1az3IOOlgOy2w8H0xdd/ZQDnhZy4guhCps1ng+59Q2Gg
1eRWGr0pSuLYn/f5Yo8eIYsl2vHA7SVPhlhGPOwZ9+JGfo8NMb3VH2X08zpkVlGG
JSqEUdYOq3kFut1ilUyvjcb8FO3/TwuNIAZ5g+daoKY2CklEIqHFaA+TDmF11rxJ
03gbnP2UP/LkMIQSQYjRDl1niNS9OCbIjHh9lQvuuZ5wmRKCaLnKXXm7IVQN8eEx
KVfo+fgGVkPVWeE4rRVaQxPSXevKrM3PedSWpgJ6EteI90p2Tswmgm/oNv342n4k
5J6SYctEZkjmqC1Pi3FNx7p2KxisgzwB9T8YNSY8B2FDLHUwBEwsYrHuEKfQCAYb
N8VDt+s4s8KXY+6lAlOsOeGa/5M1frgQ9A81vCWdDzR28ABpbLc16NH2YYXnZPnl
QWrjeAnxUjJ97faUNF3pNg8eMahDkqoqRxUKDgLHrxtj9c36cweHStRTfa2T6xS3
2//4afWiIhkhLf+TiYZnyGfOKDurYAKdZ7fgxMDEcONt/hkrgmEdoT92onNfmVKr
RA4m/RCiEM4Zo4BLYnbvb8mOEYrKtjKt91gxqKIGji3Gu39/FNZ3UQx0QhxUfgAb
aHcy0HC9Y23Fjy3jVflEOMf3oxpybWe0hNe6qdVYi01DIorDGsgqF3leeA7kIVD5
IvbsChFjeurtidM3HWgMLAywUFm6Y5x45DgabtP+aFLzzUaO9S0nxfhCpX5GcFnV
GwwxDRM+x6mczk5iIr4XSZrc97X0GbgIWx3Cy/leHtNrDcUCsTDJVaJ5uQABvX62
jwxqW4yKu5E3Kcpwy8nJmU7UICVP53s3XwDdpCL0JQ1e+Dyes1Qd6GIv7dyqExbg
rV2LJCzrnQWxz54UADcWhaHid5y5eL7nWCuBiySxORMgngE/c68+KMAICVurI0A+
fBtN8x4pbJm/qdu6xT+I0NyWm7VSjso5vFqW71H5ELEkLwoEev6PWDQh4JY7/tqQ
q+zWcBc5dwTgzy9ncOMMXMnH3gEawuzegB8zkt9A7Jz8Or8de1stjGNqVI9rBJXN
0dGF9gG+ULasgGuA3m7l4ERPt4GbGW6SniyVvXGF6CV3IDyZQsXdqGwLV48Di7CD
/cUwAnsiNEw+NO4a5+y9SFReJX1WUqWGmDl4HfQg0lJv87gvQdhtGnZP6g/0Sb4T
pmyXPn5B4MN0tExsqNNOvavn+ddslMNwDHaXyYKp1BFbEv6eGj458wuqsyYxBPX9
NaKgPxoQcb/2P+pCV8Z3l4/KFI53RQdwUvYapGhbj90noQkmsTxq4tdemHCVTeuA
PBTB7ROw6y8pXKGzKjq6LR6oVMmwYRH17e+wdj/DyjYF2AC/IW+hiOW5NoEnbBiA
DTIASNeGK3Swu65bb2ELuxWu7oPGU1epdeDOODK80IKBenb1cSsoycu43hDLXYJc
aVfAm8D5N44e26m31fs2gwYbx/xkdKmlF+rRaXlGNQYDOTOeJ/1p0WNGkvrlNQON
9ccXtkavSuGQh4N2RkHP139N99OfiUMTXrB6aEy+vb9bDEx4bpLFFksqdbUcCvL8
IKYIhuPADFjc2hDXF+gRJffkbbnhX9tfkz9j7/KrulmzGEGBl2rLUSv4XPDY367m
L2krvhK0EriQ7gcoowSsan4uH88qAW6NsJQiKXFHbMWumNurwCsmGDVLJtwVSXw+
Q76ViYEezVrfiY0Vf2jI5frFxuX/yO5nwz/IL1koRcsjoNFoB41qBC8hXgQ0OGUa
FERYj6/Cwg0UJJt96XmTzf6oM/snjz0nYgm+ScKwMSLoBtogGHrubKQCWEnVrW9q
PJxd4X0r5A9oQ5zfdbstW0eE+QaIG2CUYAfCk2mq458xzjrJbV2NUq1Ez3UmLrss
ir68YjdoN/0nrhGGXysqEyInkBKaOBF/3VguakvG+KPjZDA+lYhJPvT5fovZ40cC
dd3/vFP5ikLeXPbA+pzjNF+yKPvUnNfVj2XxvxjlE/3gLaS0vlLWLbUuMPvjzmwF
j71Yy3vHPlwWHmKzo3GfjIQiDKDyNw9zFNKoBUrf4+cTWMRpMGfMSGzHmIwQszZt
oY6geogXBoipo6NrmMHoHbV1eA1uMBfo4i7fw9Nr/APgy8uPOzg4+GccfwGspoTH
C0Qo2S5WYeyiJvTWyCb+oQcdLqXaJeR/u1L2JjTtZyzpVE5IxVVIp27TjprLmtBL
nyjLdsX2FaLlz4MZkPC0TZFjlTrUSq+Z6UK0q0uEdMUCC+SNUsn8B9eHC4cHRVDB
lDjtduMtE9HGAAIkGOQF9FcMMzZzz8DvzIIZ8GetZKsyB0TaOFips0J67MzgS7FJ
V47JFtnmlqiTVAuA0OAOAJDBkEisZF+nOMoJN9IKlb3j0anpNnxVDPBLb3nL8SwI
jRMFpkhQuCMZfIXnw4Yl+oHrAOSfKmiKR5d6saGwy0Z/CAoxLuixo2pcbQfh547m
OLtISOmuFlErlZFsLtdVpBnzRLOa+bhW40bkbgBDKc64ii0ONf3uWT4w4D3/fcs8
j78luRQCmTLvrb0D22BNtS1Ok9asddZXDcgxHadFBYII6zpaktvmE5yvFuDHlX51
DsitvLKSZSf6VXJnc+VTeP63CM6JISbXEXYOeUKbpG/qkaIMnO7dX3sXTgI5njco
7vLLw2q3T/0uVq1tHXCwFKr6Ye413wEoR17Ahw4tSiR3tZrwKlqD56+SF+rOZrqE
eQ/nWbXVxgCfUp3ajfW2uj/itVTBdiYLzUZd6YvirolqRqAdn+nfXEnX+bCH28Vz
i5w25iSHwofLLyNsi+4xRaWfRaTNvM7B9/aZb6WYr/q5AvjWcpDY2GBJeJlQayN4
Sppz4QKN3HHlRMG5/jVjyh9FTTajTtxTgInVMu3LJpG1QVTpuBufqjtGlqe7CL59
1BNJLkc7gw/uZ4ae4RNKYRiEIuOJB2tqDRG5bbVaS38qg36ax7YxqFOeuiXP2NZN
z5GBCjYKAXEQ6Jzi6wX7pzQGfKPgvF9sbDTX+et1o2ALP9yxhNNoIrqdSCG5hWzE
UdO26B9Fx+Y9cxoCTOvagXLkwEw9ADLO9OZZ+QwIBldzT8yl/wnFNZEg9nPgsJQL
V4t2+j9k2caX43MT/LRHOSXrPXkxNzl2Ddrb4vVtb3pLS/Y8guHxhh3Ss7soJDFz
7ZXRUypvBm4RxmvFkgxfwzsbEPZT9HZL+og3mCPyNVC4M/H90kAFl+QA6Bl39Cdi
VbXCggRCqRBXzQEGwxMSJ+yWJ8xEigMAqBqyh1nvGmX5pUc3kHi4cbkL4HQonHWs
Oy0umwWF98mmmRwjaqY105SVJy8ckOUsPj2Rz2i4d0woAqCbt6k/qneg2fZmwbZk
tZItH3hSKvBDhhDFp1NF8oCFIVpMM8B7G2VQunUcL2lN3g/J02ESZzVOHTcbBWdv
jtgRODnDcHipGBo7aEkgNchET6H89/TunK7XcLHjW84OzAzNG0ieESIKKlvJjCu0
nIw4qURWbmfYOI0ww/gH5MbAyuZ2LFgOnysPAsI3TyGB2IkN1GqMq10uc7nxLlHh
+Dw7bNCgGSxt3LmqhaS8/M9QFEhi+FD6KdUZ7NqIDdxQEw/v3PdNQcExJgdfJS3T
cmspKiIGEymgqRsVYWaqGxEoWRko5PZSgTk3iM7xLG4xbsVr0VXR2uYbtRY9kKb6
ScVTdq3MY0+t80+AtSXtQ1eeT75Z7RxYUS5TXvFIgb8Xcqvl5cTk51Y2MeLI7LtD
O83+HpT3jDav/5jOA2/8If0EHqjufPNM2CBqr4zkO1zk6RUxfajBGnnL8Y945TMG
4RbOp8fKC/AklWXPQyWX2sbVQ8kQ/QZWWq1+xTK0BXHIM8l3Y4vRE4Jh91ZAOEcV
qqrJiYzAtqV1Y3qGo10fvWgKmbooaqR2Ca9yw6Xc3cTyrjzpNL0xh+N+lvvvK2SW
VgWwKWGw7zOKNcQtCmgk/tfx4xM7lAYkd6rhI/aPoVjSwD9YXuSmmWTPcL2HY5hf
Hu7reh7GVb4mSR5XSoAn48+mSBvh/RUC5CVojVJUxvSsUpTtYXAaULrbLLybHp9y
eV5Cvtdm7Pr2vR2ihTmjrGO1WFHcgKGhf0SRmJJG4fnkev7hMIUEcLGtLF/Ouyq8
+xn3pgci5yHJFjnFHqOgDwqMa8VOWNWXElU8QUeFyo/jqrbpEJAuUUrhc2aoPvUj
8gww5ek5b+9QXTGcThV+lOWvcY4mvQM5Pv/cFDqF9K02Q7VsIDwk9vT7iIsGGhne
OdCTimpkhAOEBFke2KG6h2J6deSnpV+oPuh1Ks7Y9YkUw/odcjbaCoA+AZSS+Wxz
ld9gNskUxiepxhggONy+ZOQUyD0iCcxbg3EYnwftJ8OVL3Vhqw1LqOAFHkOCjrlh
kXlHs8LsVwIGQJeBOt4UUZvia6MOjxv/GLQJt0vrt/TxQEPvuLuh+NCFDyQZClw/
eflxd+79yObgjcErkdQC5YRKUa9Ke4qHrx0cBwRLnDPQXmTKMqDIPPil9rDyBxvK
MPfQVswYqkk4mZTXhwCwRQ1wIh0C1zxjYh73Lq5XHVGxIzrq96YOse/QLAeIE3gJ
sl8hMcPT6XSH0BNZtnm9ox1i0TKKw8NKtZBnb6r97ocsbOdk7VsIWrXDJeZKPFsu
bWc2I+MK7WNZWx6cMiIPEKOZGnJevZMax0rp3AEwXeuSG1mSUseiFsCupE6R8RQB
r496BvIyEwNFD+6yPkRq74MOrXHRfOQubpgUqBvAagIjsLmp5GVl1Tt54QKGMAf3
kBj2jRiBPjugN3Z7otkvhmDxjYe4cjIPk53MH6H5yVF83V6DqpZCZZ/CXLIWbs8U
Xg0SJjJrMZ2XTsyI430O2pUlObCGE33fove8MFWpwjjx/jmExOS3zzdDPFP5i+/g
m/9lgK+5eMZ2FDNmEqnC2zhf4hYsSILQ9F+nz7q9Au4IYZFxaFsDrGmAlUGGb22i
3dhRBVL+IcNkqStZcRMtDWslfPFhFNTJTRP5rtPXiaFMoWdaur8CkO8s2/yZcdvK
LC06Faf8jTpB6ZsOq+tFjocLv66yng+8tQFm6126EJsPW2e5T4fWXH4PZC5gKcBp
x22UNo8eBgl+bUkZ1d1ZfKd1Gz8CHKGl81tLjczOPhHsO2SgOvoHWEavyhb2QR5E
qXQbEfisOF/uUpq031yrL3gI4yFUthih1PqtA7EaGFmcKEjHM0JtAOdCKtMDfVz9
XdBsQwYd9zlhMmiA3jbEewDtNYcAWBMR/VB5mCAi6PTyYJK5j+imprCIYpZiPLLj
MDouVGXXx86w+WzEkHe0f758v6U73YmWdi5fDgN0QDKQKwYfW6ENEchDyWH2m+Zt
Fd/8BA0FoqGvkzJAmPui/UtlRJnMaRfWBOSrx5u3HE2Cxdy+LsrApVHB4oo/QLN6
Qglc1A5AknMJ2uJcSSETVMC4hz+pAeSnoEF/1AsOTSQq8mnFjQBk+xKPr3UBT0GV
XEToSuCxg/jnr8PoeqlZcgZwF87R9hu9oJtPVr9evoRfy5nyXwwUQKUqDhDb+UbX
VEPTzJ55PGYXPdmdkgCL9uYpmWsS0dWs/MLpX1rCyOLQWcIwLAtVzcytgJghQwHN
q/oqClmBHi2BaU/vQwS3YRDbnYA3KDCaKL/uwY2aQqyGDzDPypt97yISdlLuKe6W
KCxFT3TJ9MJeuI6A3l7GJmBsyMW0aOiKNLYOnF3d/2gqb/d5PShtJuO5tKRDKBQ6
br7rUSTAzJkkpf9OougD+cb8FUxnn/9P69L9XxQ4ZpokEha9WHXVL6d+WR7n5pyA
2t8rdzaLXzIwecR3WGSYuFRctMwx/uSMVpJwTMeb6oSOqeMFXzfqXY1qn4jnmJ+Z
cAPcWEuEhCYKDenO/LDX2ZNWbLqF73l1Lf8bU4/hU9bwC9999rjRW5wNa2u9NDXJ
4WaQVqfCAqSzA6/SKIdJfTihmHWIxSkZyAmhuB651hw8DBCCv3cSXGVmdDV25EuO
0V0GBuB1nylPluAh6obCtVKxpWzJvuueSnsd3ckcCw6fPX+NCtmz6qnrEztIv5s1
RrWiyPoN0EjwYopbOBLqt0VymQkfQQNWctRc6F7YDjBmVujiGTisXVztjSuZJKaL
LjTy7Dux9vmdntXJw/lO5HFkL54YK+JuRu4A39JqCto66FoTEJSG2TN5I0Z61Wby
uziDUJVlsD+rbZjrwijvpfe8hoe+8Qwdtq+1b0qT/2ixXzbgwQkMxa3n5gVnLaY0
Do5UIPIcxigy6aqjV5VkfcYuDUuHxcF0NP86rxNc3LVJevp6Bv38JXPKq/4R+lJI
R6y7xJjVV46BfDHLp/MWiVc06dTPeJCZlQa02YJKl/AZFrU1bbIswDlanXhP/G4x
ZkAoGylKqHDE84sAbjJR1/NELsJfJBmmTNIjxmv+V/B6SqRyHPXglsa5M2Sv94lq
c2FgZr5gwmEfHJxJJfhsdE2oJwj1vNpizKJGP3exzZEq53yeL02fYAHpZIG9rlHG
n6RLRPLuuYEeyoN7ObSCjS6xmyu8MRIUK7NrMbutyZiQbIDYvkE80deBBfN/Skfi
0XvocxRedDz9oe9CLqompAKcTKEHp5r1gwjLzCtudVWiLTl2LEszIWeYmbD3knlN
iH8/Utjaz1c/zWz6mV1p44X87hRohYdOSFY+LKeCPjYjrBn3NmameTSMyGK+rY/b
Muf0zdgKrAG7ETYJxUQSUDoRLOUYhxv651Rb/wQp9kHcMcxXrjL1ZY0NKfoTMVxn
alzyXEBTDNx4QggbNPHnkEfQ7sKPG0kwGQmozPPklLD8bjS15oGIPd+l/me5ExBY
sVFzrBECuCoxUS2kq2pti35jiaGjPeMCQeJafTVU+9Gu1PwhUun+m6ME7cHuqIr7
kdAX+V4/ity6bi5+me5VUgGE0sAdI9Ld2ThIMg2DimBeh3YRYxJfnVNARbNC89wa
uIA/fOrYH5ZZCJK6M2UGQNGGlcVJCWXQfbtXmvxjDRg0X7JRPMVh30LgoiWbzd30
9Ev7NP+0+wenhXFKxDdgPAv+ejoIddSY+AAso3gnjO9XC78ysNaPbDHfiHh24KZo
oqEAjzNIEXvPt/V4mr3+A/K22NpEtRv/ikI5G/18+znUOpuGG9uSF/v2V384SUlT
IZyrO6+dCrNg0h8OFl31d4FuKF7zNBnxFcMAh7lY47Mlw3vXQhxQ25qobOTaZKHV
OWOPdDqC85L/OS7gxTtpGKrz6IldpGIKCnMU9GZsKVUutn195yktAjsN8n1tThwK
e92QGEYWCqDAnakSXG8yyKBiXAGfy+b/rja0jn/HU4rzn6/x2C3qQ8R/O52538oL
yTqY8/TzZUr8/muS3U3CFZ9NEpvv14U4ADyCQC9v8SUgsihXfWWOsBE4rddtcYNO
RgmgW0hW3rGT6KJDgc5PZujiws0nY+kInHhyDuh8j7wSfGaj8mVl+oBoT4vLn1sB
SCe4uA5R8QJch/G89TXdNgVagYEsPNY6tRyJFtuaVrovEaNDnrZ0+2N3DTd6WWn8
qiQAWKoJSqMV44XM7FmOlBNd+k4IuDPDuY7wLpCbZPMH0L0LsOX9w2TW/kwJZ+W7
Bk6YxOGEtXXRzFsKT9R6p73liui/Ophj18XAz6GhOcipGji2nwtAYBLhpQueWxFz
GdsQKzZ8pyEuQXMzLSheRZwALbkPUNdTPK69mauJDWoay9h3F79nr32Uv/T64/IV
auqeCEh0yLu3k/Jo+HGUo+98Qnmvg9f+ZGjzMt7ICLn7CtrLd0Rp5HUj0JpkUlXV
Ti90IzAPTOg5cT+x5/jH4YnQ1kS8/qAzaP6W0nra2MhAPQmBMQZ62V/T1nj4WkCM
jzYGTtI78zMntDK37jRGkT+mBRqn+YeBQzyGwz16Ym18qkRJgUD0uuMATAsEpy6Q
xAKpr1XFc3jIt4S/8LxkNH72fzHFmtSq/uVUoQRjA/dDYq+hYzfXSahIevve4Waw
AuYsljk6T9fISPepeXS9Vsf85Cu4kSGC6HiashPCnOToBFLgLc2yYtOl1c3FU48I
MaJWhg7TdhIN3hEf2cwwyp++oItsp+AvoMwRsCJTeY3ODIOYXg2Aglz3fWyfD4Me
e5Ee8GiSRYZqb2Eksgb8LsCbQBF4yRdA2KSzloeYSfgQCThA1DG4YWuFgUam2lAI
08jTjwbjcTW2bzFNZkGVonHTvUttgBOIjNHcHIjmNBTq3+Kp37ypXJ+dP/qLt5RQ
cMiiFkGpiY/b8+V1v0ha1jVMejath/whJW/UCpQWLor7DbkKm4EBCXcQU9vDPjau
pTGIxjm1ogW7KgOmY/92NIPmMn7WYsntRonXL9wCF7EBUDEfltiEVAKIu+dzgIMT
ybZT98Qu5MrZGIQIokR41FFMsn+/ZrzQIDWWgsrtaLUwgjL2Oe66DEt5vvax/RVO
ndiBNDCZSxpX9ni8ka6jT4BorUZeMlniVjcdgwSS3tHw5jUAXc8kJfMaZ5EvijY/
OkQbw7tcnB6TKFzHe5lJlWEr8UqoTOC7ekGYgjjLe+WhymEgr8ZKtR6I186OGCFR
oG5BK80qELWwY6reHAHqhkVxPzL5+zSqncfFe0+OWxtE/STONK6O/m/5e0UWmFBk
Y7gIueFLXZTL7Ae9mQWWLyKE7cumcYuH9Sqgpnd/2dOENOFgk1bK8WkS1nfWTXug
dYLJAlShZIA4RzTSTH2pfhrd1vyRf0kOdFRl7apAel947yjXN6OSQFU4MIuM6QP5
6r09gucbJzsIl0ou1urkJmN2b7sMBwT3R7Tl3HIYPqjcloXcuMRN5IrD1ZMwLWtG
OwrnvNR94sSQ6Q337vxLIydZpdzkbWXQ4KYnsFYFSluYmg2TPmmO9gA2YGJ7wizx
kkr5i9F/u8IX40gk3gBP6iOkip1SCygBGbf4jXnLQvrn7FruEZk59ARI+lK+5wcO
oop3ybVi+0iCab1W2rX0XtVlqzEK9lUHMI+GfjIdvpy+gO1OsdiaoD6fTqrlzKuO
tzWO1akGNCSWfAv7Kew0KEr/PcvWLxOwc7kDjUim9cVJup28LHWpReMM7c9VL1Vj
vLWV4Dk2AC35yA/ZWsCvDNX6V9bqVKJD5HqjAAxtJjGma+TzQc1uCBg9Djk2sBvm
vHtzV9Edn4ef2mkiu4fTOAmytfHlm/MeGkcId6ja8vQ45Kh9V0taCsUDzsw8ZABh
JUB2lx5AYP+Tjs03nZGt1T9jyp19VOQDO91t/CUdBfvpZfd+hhWu/4QU9GHKiDC9
7WJIDDeIGcg/D3c4emtrJRdmYVqJjarvU1NqGJTjWWeJklJym/L+SOxXXzgIVz4e
MpxiE8arvRS3lxyAgPgj+UVYOW0dVNgCrHgfyW0bWzM3G8KbDk2DzieGrNvPZNOl
2UjSTmsdELGmZA8WgkrlvymeukpZEsvuDKZBpKi/kE9C1DdFQUkWsl3sg/4YV0U3
OYvRZVY7fTryNDgmpOGxzpIGD16hdkDi3PNMnXHpQdIhgd2aop6VjAVPkDUG9hof
nGRFSXBpfMyWcpYTNUHF8xGToyeZGtdJy9ucl62oQIObS1sMGQ9OktShpWdW1uzL
dPQJKbA2aWlKT8cFIK3Zvt9Eq5PPLtKoQNU5DGOXhCJ09vpugA4XhZ8004I+sbDR
D9JaxOkN5x+YxzkQwLQA+nSUx97SnaN8gmScAlkYR93qGiU1+O6LpSl17bhG2yg9
bfKmri5uyHGRpKu38s3//GCXxkKlPWieRv+jWcuyhBknRFPMz3HZR15KlsD3txDx
MAT44v3tEveS3CIyFpMIbmf22tzB1OhbLowfmKaIwF6f1SQSzSE6LCYdgloIwhMy
POduNQ50cDHaxeeLqAPJbbxC2YXcRhxwoXAkmLIUBskBw6m2AjmpuVpRjWxXpGRK
tYxF0PrGP0wO+rS49ZFarf4E8rcrbJJk1/rNqBn/7xuYTOVqCJ0EkLcZQZ5Gy12c
A3NYJrEoamXd/YUUf4bsMfxZQHCs3bSlN3Y3ik/PLXbznnckAmwDSWbxdJD0+OMw
TsbnDyBHW3XkabjN+H7nyqZRybufReXqjMMS9vjShLgDgPAQAaH35eS1s7bKKwE7
zBLb1zuGhcCE1HDkZjwJT+DNwwpZWUx3vZucYlSzMWvGhrTGFuVjTYkHt2sgFIdH
GPjI6ZX7fBN9lcRLPl/EHWkp9zTBkmyQ1l8FYBXUUeY0a6xfK3gndHmMlUfiZvW2
HWnlc9DYxwaGtaAQC4XUc9wbsNSVQbPqDobA745VhGM9ouXTqYHtHGWLdjS1u10D
l+A0gRbMpDzmLMCWBboQrRYhR+0+4mne0dYLOH2MZlyvhuJiIUA0QtPUuwsm3PTY
rPS4BUugTFYS8rc1z4JU7JgWHIT8IqUraJV5jNzeKJZ9ENjQwqHUVc7FPdjU5rau
p9W9BquXx7r19TvB0EJ6rUPIkZwucAhZ17E304jnpYRpk3KAFj0xcTihGA4yuNiZ
eCmUNwnYkWXaqW846YM4E6L25j80uLskveJxiGhqhVYMXRtyfYYBQA3xQPduNdCo
l6WlPpPYkU6rduUjxJCxeP6cRQc5kqkfggp8bmBS5wl2p4Z1CYkJPNd9aRNrheq0
o9D5ugGkhhKpTwATANpFtVYLqq8DWoH/gU3jLvn4NzeM/oLxf7qnq4bKt26tNrwR
pZA/XNe2nT8OXwbSxWRftTPknVCiFh2dWAwfwNXwfUhMYZSuir3KDEsHs6+YYSTO
1RUQHP3q8G8lSpRuoUBDWXmejQ2kh923b8pDXldHXlOmEM1LdHC68KJgq2zmFZVd
ajl7fOWKJ5lvt3z2HvQjSU50uYabigAa+0Icx1AC5U9oRe+fE/28K3FegUL3kAmH
71nhFT82Q7FDKN1mqxrZA/NrTw/ADEsI+GgmsEptoktlG4InLY+CQTjX0MmV6Umu
aXfPg0MLcg4k2u2zHUu5XxfVeKIR4H2PPZllY0RD0pMPHEzOEypwrLqHuZpAkke+
WjMV3nS14a83MVV/oefyib9h1VVcOVx5y0YP4GteDJPM5Vl8lHqCqMYo7cgSI+As
GtHJQFs4irem1mDcoMmRRDB/p7MSJHDhw6wYU5PoZcYDuix2szQoCTzXvxyl6cjy
5OhtnVF8qM1UK4JzeUWGYLdo1axm9IFUq0TQonbfWLfsyaYG9zMI/yK0nxazb0X8
Tyz+PVoDTe5R2cA3+0njCg8aJQ0o8YGHU4kIt/xE+Ps+3B921LCfi/NUo6U6kUnM
zo6rIJi6lN2YrFiarD72HAjR8mt4XdquhUQs9zyLmr+afzsY/akCUj7WWvrNttup
1xfm5ziHZ7lDjgSdEccAc1KCGBHEzrXzrGq/hs5wX3IGVMpYbiYZG9vxE7n6uhXR
9RDK4/KpYzCEi8Pld4uakmvmCXXzI5le2BcyzhZnKEGCQoGOFS4L7077BHuCglev
fwQp1U8CRjiGu53KXAoOzXNcYyC43x3V8cCvXstYbATBpLnk/F9OAJyLAvAUNtz7
TL8cSsozLWt1jZT8m/XL5oAlZeOpy2i1go0GliPHanSbvYzNB3+N7xQGUHIlRYBK
asZefStIEGCIdGK6zlYvldhE/t/vqYfCFWAyBZLMxAOAs6XOD9r1a9WvaadyKe42
eSEjtYuC1OhSZslrGlP85qcl4Ydn7U6hseabkGvvl0I8snBdjdbx8c2sM3F1ifd1
xJFOrAnDgnf1j420DT8fzSJ1upx0pEo2nTQ8RWpgaalQ/olEVu4s7TA3TIHIliV7
jPCJ7dLE715eOJ9sJQEIxxpLmgDK0Oebj80mSZdb9Abm8eDBphGH7gjcEagF/cKb
extCoUuvSpcMg/ccEzMtZV62SLXT8XpF18BjLxJ5MLs45OMHS7Jl4lBe+KljNcIe
StjxfFUp12XwEpArvLSIAcE4zkMsSMms271WIMxjdcxA8hqEE81ZDzWO9fF/s+g8
MKTi7Dol/SwfDOA/ojL13gvqf1wkZDXsaMsHI7U24zwlAlBAjJZ6FEL0uk7Wo0gg
AZ8qEkcLPlQvXWNNj4HYQD0pTj6+WEAnnkQQ36D+zPG7s1Ola2+elFALi69gbJ/p
Ssg/vIbiUi3gMuBaqoasdIFWGfgRH4MyYEmYOKU0zOAWSo2bOvRsUfXD9qDaSAo2
+FAzhF1shNOp1CtgBHaDMod7ws/I3TSumYuH3vWV0GO13mHVlXc11AzklAk/GANB
OBTtI2JxqJb+FEgp0B6RhfZPMw517+u6Ql2LXmJCXY4G2ElrSybnstkGfms/9ExL
yuFzNcogXs8X0RoSMiMWtg2wtbJmTV0fPf/bWjMdh1+NAQSAjw8ZUerSyd1AUavk
uvD5TRj8uLw8lVurkTWfRSwvffQ+WPWlHygj2asOWWB0wsZYnGUjCtAWeO2YMOO/
7KIIlYzooOeU3vNeHASRUKe6dFY8JSkdH6zAXmpejiNXZsWp4ahIWEtTBfegtGeg
r0qgdkqjvmx215ywUktPxpQ4zAGzKpi3dctFAXu7zCqQH2RFMB55Msc0wBptnB6P
QSUHWPZbwCoijEBZtyt052cLfNPLH0OJYg/gBO1dQ/AkA8l8BA6aR9qmYf7gaN7X
59iy68Hnts6jMIlYEOmgTNfe/GuGiq5tiy7wnI30J8Lxi9j+GNp6ypR981eurH2y
tTy0bMeUShOLeNq72hKvZcLqAU5mXtdO/IWPfa6jfAl8erTHu3/K+3jGJsPvq8xQ
Z/wG3lm6qKotraTcXZ1+xaEWhllR7aOQqtF9TDL/1rMevcZjC0y+yssupzXizQMp
GdQ2FnfhzMmF9u6TsZrzyNcuQiXKU8vFIjUr1hmEgfq2q7qu/QXM+igIUYwWcH4K
IonygDnwy+LOWncZBToYOD6JVjQoX+o2LnZhZQ3DEjwbEZ0gCW1UZ9DKow7VRQlF
iwrUNEl+awxAHhSvhb/ybpxxySpsmzPF5roMKfvR0y9PswmR8iIs4Z1p0u4Dgo2X
8EFBlimOOPYW/+ySds/fpeCacc6yJ16MYf0TaM6XBMDYHLv554gNKRtQyjsx3G/A
gcVROA/GZRvfnb9bJ0qe88wUR/TxVTS3XpIqYN+XCh+Y55O9OfkFtz/A8IHq46VD
/mKq7Cu2BmyqxwvvxEWgxNo6sMME98hpvMKgLZWQLk6vxkcJSlCfAeCuSRv5KLA/
BfVEXGh2GaT3qRMCtSeuIVSMiFXdM0dJrSiJuk6T/PObhbNAxn+Hfyisg7SYKUZH
DwVtxmIwRS3yM8PqV5Y4ysQoWSd8MSWzp4k/x9TwDmCNDM2GrJzHDFN2Mdtk7LKJ
xP30cVOu2bpNQB26MotUKW5boz9dRICc+pJLEPCrDdYBHunrb6AhUIea3EHYX9sI
cbg536zAI+lqE9kVJpYtVzhfACna1jMi9MwSnMGJ6nfUAlCUSFNNUj/kFCPd8mxO
vzdunil3CN6CVtqO3JI4pD8UCO0GvxHIIkpKNmsbQZXaH31RMZE0QgVcK4+5y/XU
l6vwrXsuLmavsTJ98ES00GnC31qX25y0e3bN1ercGDjQDHqcs1YW8cHLqLuvMwtn
p1iHgKQG3eOb9cztLfY50vtOikfY8vvmlEp2zQhLJ2Khxw6hELEM6SCD7r8CnYxh
iKpUWlkz+FusbqRw8iD7g7NbZTiqfiNGLtjqxBoKdjQuyO7FIKWE/H4TVND4Zv4s
4KygZmDQhXaXMuObecwan87/gHK2kB7OmU+g7Csad0iGE5cTNf5UmY7esj8pD1gl
XTqvqalN3tJF8IliKOrPViBHsPsSdrqREa13N3IOmsWuCwXHjmlFRnbC4WcweOpq
QEFyhs7BfGInQFZjH/QhUz0SMDtMqL1Jfq/uZ3Xfi+xKxLMiv0uQv6q/j08jetOb
QVoRfA464PvcjRzfz4xlEx/W2eZsDljch2i9vHwVbes3qJ6mgyfldh8jkAsveCnF
n9Wc1iO8TTJkQEK8s9y9qm6zpyF8/CIfI6c+EiLiMCFK+vpmYKHwTegrCiB0cIHV
9WB1e32R6RDvpR6mViUYlHHT5fGmT9esZD/3+xjxJyL8tYxK2lB6vat3IdkS2agy
9WebmeyjhOeJxBL27mZumzX155uQQsCbxZ5uJwgEfRiBByOgO7whs7wRm4Q3dstB
UKGb9+Fj32zogXpA5yVhehLGVeZvhAr0+OyhCb9gIsu+JbmcRbdlUcF+rb74M4nD
mCZiEdooovt0rhEcauKGBX1FeIMASfrefwX0NWUa8k1MWsvSEasVo83fouHWAODL
xQljT7mtqGKMjAehtv4USojJuN3s9quaMtrr/RrJaStE31yIosQrOyuSph63FsW1
Z6fkv4zc9iOBTjtyEo1ARM/FzdAlxjydvFLclqaFW0YTXi+3kq1mAdWth0bxWMzl
OGs6FP2+JVkWegBFlPn+2gJFaWYjIu9cPsMPCgSsSazJ3ZDPWnGlbvNGoSljl7RK
PO8o8Z5FojCsKLP3AhbQGFHKwblZDgU2/rNFQ+qJn87BNI1GvQ2eD63LoSiMox83
gL3rm5cMYgLvLozHAtW35ktEGq0Y7RFk7E1m20VzwIcSzj57fvYYu/LDXZNJwZ4I
SLkuYH0lfA1rQowcinBTfmYnEE1NXzOYOpV2F2xdfFfkINSssbwowZuBi8GcvZjn
h70eJ9W3YwZcW3jUZhwuqTs4Zo7DvVVKSRCEIOjckmH2hJE3RqW3kfE62z3kPRan
irg+1yG88wc9n+DltFKlQXwtlGbpp3SNcTzM52EgxKBEwSt+n/AJNjbkxjhWId/B
dnoNxbnP72SJzx8EAuTOndXJs/Ajj6iHV4jj8wzcQFEv6k9OsB7wU3jp5cKB/flU
Qa5W9afGdXsnRxqUN0coRJCtdBLDRHZ1dLEO6/hC20Ivg9TnB2718sgdnrFrz8R1
wah3oHgqWDbeSfXD7QKkHBss3ykzLb0k7eaCIUkG2OWf8LdPJ1+Ak5MzXk9egjDG
zcRD3IBtLhlWtvKeXdBI/9hOx/XdmMo/qJNWiUMmhJRmTGEe8smIPARxqBgJrV5S
EPUY+kWGQEe9y9jQt2OrPHCJR/ZQnXx4wf1+W5lmxaTU76ZfM+WMPuAFZxtRHIim
pe+KLGo/Exvu10+dieRpvDn3qT6TTU83FBfx1fTKke2R3dhglUYFCD844BZVEafV
F9KWTK/vaRiDAdwTbw6BNaryz0SclKCkAmj4L7PYE502mEh4fxL/oEZVD0ZGWz25
FQyAnJMbhlX0gy6TkSgT0lFKJo0AX7Qv38/xiERpxmaNh4AicYHuGd4s+dXyR1zC
cGACoJWtZioS067b3TzVx0/pWFceAlXWO48dnDhaEE/+Uqr0dwvlG0UpV1T8DK5f
7daH/1GbXv7/dq6q0/Q4VCadZOaSBUxYUiVYRRsoZNTD6Xi0evwRdIT4kHSdfFY5
JW6lveWuSaplOuxF7rgp62FJZ1oDMkYOnyR9KGyEwtcbiaFtgIUsd+Ry1SzkC/Uo
iyThRKphzeoAMG8grWM65ySyNULKLXJazK9z7vWm/8hNAeKLnpXRbNMO365VHWRH
pVaiSekQRGZM0Vuninr7Wdy2iLZsmn8LRto7FpGBClPlNK6m3JmOMKj5VWRWNMRK
qrG3fV5T6KtF8rBDqNFJ+MXV5lpKA8Lk9W0GDZmT+dPkOMzCkYP5oZjgLA++VBUr
SX0SuFjAQ3dNtr+F+8t9TOpZ5U8XMvjzzZkLM4FPSTYHK0EOw8a7nClgifTZZD71
NutTvjQfXAeV94S8hRWLDbNLcQDztpUBdknpK4UYEbx7800f6zyhFvrTFmUIRqIy
QGLOz3cBjGpzVCfLNPYUZzjupHJrC6PEMygbi4HaXUGqPa+5bCtuzmdQIibhDou+
Af23buG8BhJBEq0xs2ncU/2K1/pfGF9sZYlO2KlYVAmV3PWSgj9ydcCxXPdqMVVk
9zk6uK2b9mvd8eKE7PvlCOR7Dbl3d2RXtbJxR/eGCT+vMK07zUqSPfThbYOkawKh
poeB1ibtN/eEN6gQhqYB0boPdorbflkoIHfgijI4VGG7t3muqCHFkOrJnj8YdwYl
ycZRqM+esrCRa1S6EZZzoCRG3lGSObxcckyneJn3K4DlXsWg34yiApGnBS9uMfIQ
TQO238hVgNlXRGAJLjLpMnMexvzCshkRYYMVPMMBCy+Pub0rlt8PWS70C6V256jK
QMlW2t/FVAagGab33m/ZwPG/iwZHldAeyyD72+TJBPtaZJ+NcYi3EWF2PaiJ2QN6
eY1AJjLlI5kVyv5nNZSUEryE0Ll7HfW9qkHM+crBDn+0+61/iHNa6Cuhu51P+I1d
dLF++Da5amRrAeI5/hW/6ZmqjVypxY1YNmDDIDpQSKlNBjiGCR8OhtcM8Gl7Q1mQ
g1IJaMZE/OuV+OFbjIvKFe3ss8LX7+ByfgqH9nYrB/X4ngDA7HzTKFSp/zU1Lpw+
gPprzDifDPFMVRGBr6tROEN6cHLwZbTkTiuKSjflDqAfeNXDY93T2HVBr1dQDtrC
Iv5Ow6dq/nJYQfDSbPbMRGkWPmaBgFu6fTkp4i6usRL5v8vVsrvNSFSv3Hmv3Fqg
gKbDHXbnmCdyKH1PKDxg+pPxt38m+CtzGNJCXASSUTgWvyP/4juYvf2zqwoV8YZd
PRXC794vkC4WOxFqzCg1m7efOWoXjyeUjQeiVEZLr7aqh1mBcnu+p4VO/NREqs2j
/LY8CeKzVKhzDdWWhZSJDBAdTMA/DqvtFF9w3DCbuzfNWQqR93k4NP/Ypv9GE+a0
Xa9ONNc8TteRzW6Sklvfn4JlTRbBfBSm8CZzG2wATKQH8kgIfsTWWPxun5GCuFQ+
26THVOnHgHOUgJYiyTrzQTWRSzZ6Nm+Pp9Bi7Q4S+sf3NbBg1WcM80hf3IJ1B0Jf
AmqG4bH2lCbjInQsTJ1lzsr94wkxQp7sYFoAloYbBaUFzllnW7YyZIGaIiZf6/hQ
PH1mobqYAZy79YbF2n7FyfkmUV7Sxr7XnofP9npWbCoGD3+tWAFecCKmjIBIPzG4
6JpQcpcKAyyyD/Dn5FUL66nYhhHdqdHJuOrKZB/6CAHMw+pntcUx0r+aOFqzFqv2
GJvRVQ4fZM/r7WVxJupz8CcA2QW9FsK5ZCZYgO0XDdDm/vM44u2vEIbksBTZtM8M
qj3Fuy1q6dIvIU7DGxyMZhupnW/2SNGdqeNIqmx8RUVx6OBeyuPi4dL5+QTTkcbH
S6LuxhNG6lK4JrjsvLXfTWTDiNSfQtPmU9roHlTS9NuzEDjwZm2TUGKyUDPWrZ/G
jk+H3PekUk2RI8kqdz9ksMui2SQsHsGv93KUV8hwrR7e+Bt+CXtRfwH6KPsDwSQ2
dnuvWwRSFurV4cunURaqmLcGlMXaH9i+4QrhKRSs7QLMk/7hBRZC7mPlhk5Nqd/v
V1ClBtvhkdYh+dqbf6SHakiA6HHLantCQgk4bbZk/Llhz755htn5Mg2npummcUMQ
WR+LKInVEGG9NJ1M/+6NI4C4pfHs0qdTuQG+Onj6DW8tp/x5P5GbHXdoSX6uui25
X2N5UYZaW3/lD30FyPL/K29jAUHoQd0i8MVt+gYlJs3TjbW+YFJyqcqlPN8XQdwB
r95wGA6aBsUirXgRn85MqkiJ3Wijt7xseDJrWRuzPnpQUMgjBgRH15As3mZ6IckF
PkY9ZwjyLxNTdmvKYlnA3/2xVFDQvedWPp1MvLsmiEc84eSRDRxpYAUtfRD4Dr30
FUQQyLwsYrfhZ81EbIhjGgR63C3rdv40BJljHqCm472eiZ3+m9a+77szZfLS60q5
5Q3Bdd91sDEQsoXxp9HZQHs/JyDGx82mdllQ1xoGbmMF5saYnH4g9esARwscI3XU
bnh6ta+zxxHR34Mss+I2+whUD6jtH7Fdn0clWA39wJ8Xd/Z3vICRKh3jZVQFVluu
iG8TsUo2F3sWcv+vB/cDp29fT69lovV/vcFIKpk7LMSaR2JyhfcFFsS40wZ1x92R
txBEPp+V/HZY75viHSgLI6j2DZa8S7U4UxghgZq6fzAmRi+KLwhjLRKe/DBeHF7n
ysebDWxQK329naBEeQdX8rycKhFtSzbLM13OanNN3kIvg3//kBPlsFnbFqTOOXG4
Fc/UBwq6Ga7j8tMNgFMcFX0ART8vOJPEUS0hWKGYDgw3rcHLmM/pxzB7ajFdRt4i
ToXl6oIHjuWPCAcSORVMMZInJ3Kgn0v/GFRrWHZ4dUi/JSwDYDEjxfizbPhRlSIj
cfrv7VYsCe1bI+hA4BAdHTTyYgmRYKcKMFaHORYOvokKmRWi/lrsVEL/R2YzXibC
19bo2h213jP3zciLqD+KDzHaLCcJY8EllwCqnB81tDg42wudLFIvh0qFKpCodvLG
vVkP45pKop3mUeI1kFvzpd1koiNOuKqJGibt84TGHdxpyODa7OTCbXo+9QqKaYJ1
OZMamYfoKD49Tarr5iMXhOn6L163l64MbNmXVpRQ+gGKucl38mhrdu9l1eEz1uJC
ETM+mvUkXrPFxUTHW8+uv74Mc0s3IUGsmWaGYdXI/umpjXJaoht9suw/r3Ff+1b/
Az/lXyDkBM+JQXXI6ebkjh4plk4VAgJM5Ro/tqTbUAvXxSvGCoNWjvaWuMufR1Cg
8Km4peVLzx07ZURqbSN/X9RBv88vALTyg35uBQEWBK+UsCbbE4AbQ+3pm99v7Mpd
XuxyTCsx60zxHHA+TgiiFbglm2IQsiSeb+rVDAB1C1yA4l84lzuPlhgp5wYH7ytV
kVPGXWtMtUiUbBKVzq6Pgzkc40eou7giuLaQzIYuXTz1GY7Rxr2kZLEvbKQosjrp
mM9JHtdJNh/DIBGITs4EIj/+mnGWUKw4bqOaCtc8RJYLgiNAG5Fos8iLeODgVJQG
H6UpZadYcOwC9p9DWHWD3/SDnX5D55YRli7BDT0dT7kn8VDwX4Gats41uSvqvvc6
sMr4Vuna09PI3ocOGeEdHAeNW6+DW4HJBI0PxsY1cvx7aCswBBlhbeJh02IDjkCM
t1R15NC8xDYJKvRRaeMjamwrXmlRnNq9fT2T6JOSParkYlzPq23ywmyFtz0jS5q9
GDOsGgYSu95+hixak0qskdCjZSV9SXn1bB3nyBtl+Qqua91duc8vc2Kp8fS26g3B
twfMvHHJO69l4DvJ/utPp4OvikLqPx6VSwVSEkhqMc2tIOXG8DUtzdmkRfJpJ1RQ
VHimdfZyiQcgvlFaA3DIjhBoEIVX545Kimnx9kpeNj82gVAQHeGWnE7QFncclCA7
1287wueXmqXzn9doH+IQdVMxGBGmLLydgvjTKsbKzlmEBzFyrt1M0RryHdhJgyJE
fOERVdQOS3DT3MU3/hW21XINcXasU4dmhYSvQMdEU9wS8itSOHC0Rr7WQb12XF00
EKZm53k1lUiQXXGfZbTx56nzJX2nACrz1Fc0Nm6TZXthzSf6KSXLhZ20VZl7L88I
pJHLznNJhVOo5CSNGgRY1ND9nNmC4Eu9FXRt/b27DXkepntedJ+Wo4+FO5wSD3af
+Pce/vcYYGpKnW9q9SLU1f4Gi609pujGFSDSvrCesBEF6MTqMCSmGx1NCfQL07UF
z6X8FoxyMg6tkZtgzNo7Vdqv5Hmh37naUCJ25zlGY3kpdLrTyVefH3ca/qRumwIz
9Av4xoEEDE2fmPPtOjHy0spgY6I19imHX5F4cqH4eRdKFvI9l7i25bKS5hIDbYuZ
wvx/SvO6SXD8KS5r6e6Xd5ac59ncxvrfzGf61N9a2fQpWpZKqxq2q+UBrMEYQCWh
lZLEZJ5d2AxU7gLsXpfk4aOGfjkDse6L0mHNkEZzGG0lEMfBHgs077bK30hLsIGe
MP4LUOB5/4TpORT64iN2uiL5KRFXIZpZKwdfqHA7BS2a5SO1xkkcMB4WHGii1CD2
SgK287I4xBEhFvQ1PmCPxqkISIwaDxtjmq0UDT477+R2diQz5IWapVejepXkybtY
Zz6gRribJwCQUhUDCSeB+I+9JiaMpDaVdrYA5TKHhZ609jGrASOvVrOTO5lO7bWa
W70ZmlZ+QGRcwqugt0N73On95UHnUUB+kT2MmtPp+uCr4P+cMa/uOWyL/r3Ozrvk
eCdC/a/Iz8d/ihpzJ/WpLOlFArr3m2IYNHn2zOLSqr+4Bpu/fT6PShV5XFk89/MH
dP74e/RCHN+IQt/z/YWukwR+wmYZPfWkY5oH4D88DVn94tY+sz5Vl29hbaHA4ZG0
XxhMR9syBAeOLf/KzAx2sieOZHbXd0xYS9urRHwGGXoPKw/A/zhhnuLLkoqljp7e
qGEYE/8cUkN/YVYGqeRGMY9hWa3p/3wP1lz9Gj3e9kkcQMY9ivmg/R/W/3zBary+
gl/jOEs0uvobNFYi5phUAkRmlUxtbQSP1bcASe9plRLD1A7c7QpyBaX2q/O5GyUu
4gJed/PITtNLK2U3G+uYJ3goK4zul/g+QekumquTXUpUGaY6TlTWdGDVEjI8AaG+
0BTbHDrRs4jWSnpg+PrnXY1Wz7b3AVeAKRIKpUMQmgqItWorghSV5JkTHRwghOqg
PQ6ppvHmpjMGy97n4kIqBjXx4VbPcKRBHJ8VvQ2gbaPYL/vGbqetiCyU3RXYi8a1
2FvdUGF3COv7QamwWdjozay46cXGV31U+tq0okvwwLeDP5jXZi32Fzb3hSY7WBeV
DUbzzHREKY/KQHp5F75UWuhZVTEyK14CZ3r7W/1oxlIEkrvOArqrg1Us7ISx4dOy
K1aWYWCLBEhMoFhAbo2MITzKu8cg1SXQ5x1fLlCJOg2We4TuCMavUUSMMuc2e1Wp
v7RUDpIBwb1uB4Utx+pujeJ+Zte5TjCelyzaUhOe4E4afiKBeALs3zGzF3YYvERs
yadODMky3+hY3x8Jhn15/6AmiLs+gTDVk7e6bqI4i7jaYYnjGE6Bbw09OBnAEhAK
exQ/Rd6rmvrEslccDSnWJtA/AE4AZkjn/GT8RIzl310J8aALTdEKzgE9dYBQ5aAf
P6ghoQq0YFQ3RdqzB4/YhhxVdIXeae/nZZFs33KMh+ke3tQPVr6mSjkFlrECVGjl
9EFMR13Mp8DdqhbDQjtXhi6rHHlUcjyVRvX8E8ZPOteyaovpoWa3pGDM3YaCbj0I
9/rhp1/ZQcWWiFfzpN1IK8PfpTbzr0Q0hUP9b1RU6Umb4/zFtDf/xsRWRFYPQkrp
SRNYUYcg7/6fdJwVLI+UMnmZ09ruqiQQPhhXEKxUIVPUemxTvV48v/xuU5/oqU14
Y/vXX3sDxhZJYUpBSQEtX6hxBhW1XIx312bSxVxh0AIKJCtQpBLgW0OiQj8B4INE
Tr6XiAVf2pcX+pF36s40sY56c84cQsKQYyeElsEvE6Hy91TqPSRFFz5Pg12ktWVH
BPmBMlVFu8ksCWKqqLOQMEpsutRQUKSQ8tLvmKM39m/bpbS74MppvxYqdtvgkg+/
AgKGZEOgRF3MTobA2ap9E1O/ebM9+xHGnt6ix1cwBWIDEsV0dLXDVnbzO1Oh9A+V
fVBNzvwjMtE6E413hTD+aY5g5q0bg4A8Gh/BePoyqmCWScONEkFexs2QtscqpPME
YRMlWy+808Y09F9mNybCW39zQzIvLJuPtVuxIn+g6/no0g9o9Hd/A6nTt9hjN5Bq
jBmBc14LXUEAEJK3YHOy82phcXNZD4lk62XeiUaQMWQEKwnUMTpbr/vMJ6zPyCY5
15sA6tsf1cxLMYcESug+DuEhq4X1byAhR/jGQtvcaY3lDFY9QCVkAhJnPJoGbWeZ
atBOCuvE0H4PLAJH+MrP3X/uJlJWD2aGx5uul3Qi84OJjJvzGYGOnWmj/avdVerU
mST9ZIEegBVef+UkEjnM8l2Xm1//3p3AebG8T0vWlUCSsvy11Z4oGKrMRBb3PSen
mxViwyi/vayWjori6a//jfWf9XOxUKt6Y2mUxNChNpebtgICqV5aX3gFMct612VX
fazn8nuMzLOfyoUBxtpYiQGyE/exsSo2lHdheB8gtFN2T8MBN8i/HOdcI80ACkMT
i5WpcdHQ4oBwAG4ZFeDK336c/seQpzoKBH1N8IiyP3ocveeP5XM0FQrXJqOG6IWj
KO2/GcteAE7fRAvHR+iomYwnr0b6o5oQ8VnkLa9tfOrAt0j9AzRSxdm9kSWzVBuJ
lSD+SvfaP1DrusibDWl6hqLIlmvFiq1Fv69dTQ0dpyqN2YSt7UAhtl9UsgKsXpGk
v2/jywOoFkwrYr5pMOXgDHxEVu/nXBSxyuClixogNGcnCGuz345OdN4tUehA2Hg0
P9a9lZIZo5e4M1nTe+FsAQ/KJXDP6KwsBR+i+R+kqxkd3CDfpCXJI/YU9nwqgcXZ
+hq6pNpeJ8SAfxB2R2ZG4FZIcqIcrYQPSpt7OJ0d81gI6vLlpXHWVaB4d84JWK0n
QPn7Bxv1Ez4X85PnEOD2fm58tnV1BfXKwtgSF8Rn9rBzFDW5eEWRmU+fggks+5iN
CAnAoUpIPgrIHGgljIjwh0P4SS13tL8PRJGW4N7BG4lX/mN8dXVc5+utpAhFH3lO
8KzhAclcj9M8PyZCPX9evsIeD/2Phz4O68ayv2TtbH7yggfQ6pm6lc0LjuBQrZHB
8Mc3aq6YBZ5mrnvjBFZUqUiNSRjKM3ya9Vv7t2puueQq75ctrpYUGJSBGk0ElKAI
qrb/RWicWN/xZLmxgtXsTP0eggPhais54NUhjmtnlrPJ1yYNzu4BDpR+9kkJu2c1
KKSereszu+H1XTlIN5TqDfaJhzyhzv7GfcgG7m8nYoT1miiUZM4gbahuTtk1Jm0r
Dc/2y1yfTheLPLsjIt3YT87+TeYo62/ApC56UPeOaV/ZoEE+C6ZmPv1zxF1c1i1R
VMwIwkjUUDjFSL+r8gWTfqGDCmOY9pQqFNipkMq4wLyIT75B9l/e3Irzrhr0c0pJ
r/RYe3yPRffREI/+JDwtmmv1ycct8pAzm1ZJEBh+dJQiZiNH5XVPtbxBu1T0JGLS
bRqVsfOOdyL6h6H/7TOmiwE43lGlw6cEX3payEBCWqFMNkDUJgy/tJbnlzdcYZWc
i1uSxgACBMQwBWRN8Airve93CwxeQ1P1aO6GbAflTs6Q/Ahw0y/ceXoMSWHBh3EV
0S0Jo+xOAm9yPjdFNeeL6VaLEQacfX437o2m79theVu6+zv5xH7KzuOcP15rzN5n
lMGIfoFXie8Xl1KrTmd1KLNgV4h944h0uQti6oIAztW2+lm5FITRkBSqNcyb9uXT
Wtf8UMy5w5lE+5t5l8L3Cdqrj7yK4XFEsRggf0HB7H8OKaDSKAW9L91H2sZmT6ql
JmD47Sis3LPbkqoWo9AMRfxOfOlbBSo+6tru0mQ07pcpBUEQGExdetjuf3EwfUu7
K2SaMgg8ARR8aU2NInQazv8Jhll/dp63uCJlS/KEn4v4kGxkgi9+bLnESn1KdFh5
xZ/PU8hRu3SwvD9L6NpgLmH8QqJTmgZHlQnQsls9e9s9EM/XUoZ3yBtFsnrW0fN9
2ibtQEzcRnxdlG+Veht200SMT5IC61/f2UtCburNq+SwEYB+6mhCNp9bmIYPC/4Z
UipXmBLDmvaNv2108iyIyYkSWa2KkVthxBmanQk6qdnYzQ0sjouuoD+UBelfzsda
gslTsK9M8FGUplUHCKLhqXaveP8PAG8iTDHZxp3xWOYNb7ekwAFSKUtHvJ1uMsHh
Ikhvr3hdXcVYNqjbYk7658eLEfXHQ9VWR+r2SpImPWINa+ze+CWJO6lo2uodd3rl
7YN/EhAkyXdwc/xA7AlXAj3oQx1KvWhfPgvB3K9sn8ESttuDc+2PxSM81i4ENGOd
CaiYNZfYl/0e6mUDDOk73V3hkd1x+XiCF+DD9Rhfw9HVzl3Ml44zXjfGWdoARyvP
quuVgqB0yfnMNIo7kaSrVHgDldmqcKcP/2l+cBZqlJUugW+/OqxWVO8F5ErHpraD
SneDt1Qor6uVDCPvA8xR2NdfAuW4T2NXFi+PiY8WeFp93y0mtOC2v7EYnEpuwqqa
pxnohsm1sDA8oEjVQy9b2/f+gpf8yTIdKEG/7L7KnAuWj57qhi8YQTR0spqP5yQP
zpFaNBf4TSXqzkeVXb6ZpwWetbLUKOUxWqPPeTxKDIrFWEbhEFwQcVQOa6bSftvS
SALCH9hMvy0M20nktdpuCukv2FPoh133rBHJq6SYzv1s3hvUKtCRvQel/vNWkPT7
Dtr607Cix4BmqEl/yOB5tZrNeoR/rr/SAnyc3iVsYjXoBU7vDZFjyPTQ4VES2EhB
RXE8AnytxhzDG3gmcZHoA8qCv7EqyNlYNGZkGoBze2EfEcSWe8xPom/KuIG8TzP9
QvEel3hgSuKeqQItwi40s2DTb9UoUiIuOBh7C4l/UR/u1EWr7f9ue7iQpq5QJtH3
gQZAZxKOEiW4zTJ6OWpZ6c39jOlniqMfeFEVA+GoqvvhpbHiYgRGE1z+QdA5czMI
5T9DqPO1c5f1wc/im6cUpHktpU3XFXr4qmn5u/O4fDHZdETKsCp+EEwG7r33HdyM
ZAkdSq7GP1rafztsDwKVund4jg7LkhR8pZj0SYOT8nYAX3UDzzdzPFQ/en0H00Hg
4sA/8+LoJaHEiWfjDOt2fKNdEqeyUOXzuXDjj02uloezFUjMbCryn5LeTIiM7hOB
ZW8PhIZF0CKkqDIy2OdXZuZ17Di0msUmK0Gg3oS/NLUY08wg+abYK9BW+124aW84
niLiTRXzxvj+diZqJU5FyCAYutzXZx890BImu/Mj0iA6tVXBaGkRVGzZkgX3OHXu
1+gVzBUxd2b552RiFG98L/Yfhs45c/Q/EFvCEcp2nQqZbk/q1pM8Io6QSyPPyWBr
XPHJimVfr31vXwQ446P0WBFLpzR1MgmItm4PE82IaxnElOjp2nD7LY9B1xa8ni1Z
rdYLrgr4naMQnjPkKb+ZLozDTFz62VKYITNpbQwYJlEz/igsWK+0MrZBiysw7K8W
EVvtH8JPxnUw1z/T9Eqmf7+xIkaUqiKp8SjhwErIbScua/oIon6NT74+m8Hw/2F6
VCeJqDg36TBB599zKadL34cswW02tz2IsG4xKzWucZfGGSNcAAkqBANO6foC5/4x
FFoGc1g/thH5yNlLo975o+/SVecIlucH96LBgQVUPxykfu08hJVbzlw1G1NQrqSV
FzsDSQI7L7Kqcz2mskUOgarEEGszq1SMqtZHnW6muar3DDD6NFMsMESMv594dU6f
PPcBQSkF8+mjqPRu1VyI+2jEZm0T7qTt0pwArACDP8g2Q+B996qH1AqP0VzSMjfE
VEkbwgwJhAQ134DfXvXWRDVwR4A2T+wgNUD0idqmdq+RU3Rt9MlxtU1hb++G9Bmj
6/BLlTavqulR5kzv8Gt8IXwaFEIh1P4h9zwXE8SyEW9OMU9W86pgiy22MzApzo0B
HFVVt0k65CaUX3iNu4p+0QYT5HCXpJN5gdWAOwcsdRcnL11lVbMtvHnbgV5dvh+l
0zijZseNUWrVan39s7kmj5Im0pc5lgs6e29IGE5+DgS7s0ZXvLRJDqjsHMtnxI/5
Cn5d81QGL9Z9JqU8hUdYWgCmXsYu/Xf5BR7WeyoI3qsLa0H4O6qhrLEp6hRMoqMt
K2owI0D5GZQvJ6tXby11J4Opozpkn2mv9V5k2wo4WIMOUyIzFOt3jpkRRDrKaI/E
oXkPC1hlzyYXo7QA/6NXkoRwuOq7yCSl7INvqaRk48YcMKL3hM1xeKdioHNMOfIt
T+1fSbbpIsIdL1lYO/wg6DOi5Ql6NUKvp8gPaQu0wli811QvuNa7SICmpmG8Snpq
3iDPjI07VKzvVzL94KErTgvYhdrPmvvQppJQ0M4Sp12amY8Y1Wh+P0BnAxVYQ7QW
mfvFnHgHVjClZXmHAqI1+QWyNe6BT9MzJ+96rMhO1S+LsyWAk93F3fBcn4w35flF
Ej19V8sJ7YmR5DvT7CNpnNDxsT32zvmIKO297MzsldeWpF/EFv1wMXbmQuTA4ltW
LIU/BvmWmxr80t0sKgo3Xv7nr21hdI6gAD//MK5OwkcXzHaOynF9EvfAkqtEVa5a
tZcbKE7HYC2n5503SOVpSG3Eo0EGZfc4eIsS31u84GQ/naTHxI8y9AUpwHwbkmDB
uL9X2Jy7G0CACAW7L1sBwZqE+0SuA/+Qpx19cmX3ngytciznTRhWfs1FSG6LSm4X
KZh6RBwpW6RIbFPewQK1Uzb3Ic2vgkGMEFXLH0cAVUCf21ukQVthW92EX9DUqi9F
231F/Nb0nYOgrFcdCEJaOtzPsmvgcppRbPPwdzufvikVwBUchilirbOXMg0YW2oz
+Bt5ffJY/SXnuaUOaqi6zrbsNo9qf3J8S0Ludyk1JFXh6+KsnyZ7BMxp4aL2lOFA
LYp7LDp9/3Ol9O6pOy+psO3cUfeA6tzfVdjTmmspaHYTjlLJpteT+ivBH43PMdwV
xEyO9ffaanRFxwVvpdUKCMz7n1iVnVZSkBKFeJIgP0wJ1U7+N3lXWjaon1ImDTGw
lByAL8ISwsjl0hTfIpIxJjzndK1+jPsO0ALutkcbm77NL0pD9Kblt4CP+VXQ8F7V
BvVjpa6YjUGIknvBZ0HZdu8/ErNFgT2ozAIYSFDUfjaD76GnF7oWmjmus4nmYmDe
MABHpt2ve3fyrHH8DBbrRPPq2X8WdTF5iX2mTS9cji7qlTIl21ZgyIADg+n6SjiO
L6er/4/EoJknSfhi5lL4rqbx24xoodYBOiLSnLTrttBJWfpBtu069bKPYFoie0ml
Z33eN172PDSMzaGcLeFwMa+moris54q4bLXSsfGW6mNKBmK2IlNV5aj5MKV5FjsN
s15HAXATTIihA10fqlOiIECSxdZhE/m3TW8ruY5kL39Dz7qx1/IcJiS1Ocxrwan3
bWcSSbxwDJhbGkMT+LATcy243ncA3YDLIQN+KctwEKwNZLVOXMpkg0eBL70RDTg+
/fLNa6o0molFyspjFz5mqfTePGpDi9YmuPM46BatT501MEMTR6vp7VH4oEkHQDcU
wqlO42ZZDk0BIHe9SwG/xF52jP0XD76IuIdibOPnfMCq7Ya/iZWrue41f3M9OdXj
15pYlNPuauSiLud4paLBQo7ESAShCJgpEQrHrCYECDljGXK3MpZypyZqv4UQimRZ
x9OHNEoro1HulCcMYA81PKIyQ7K6mcJq0Hn/NBkTe9xwNwU0ulNrUPlTKZiKM5za
k8vIylVI2lJCeNcJsDG8yQGxB/gLRU4uYK9yvM0Sn+eTCPbeQ3KTFChw9fGnnNhq
pKqlOi9n/zXYhIN87YoZPxNcgYDYbPCztJ/oZryxF/+OuP5HK/ENMHpzUq35gV43
zobOZXW6Hg2mes2lrkHpCoWoExkw3c9p9j8IL6Zwex+CBB1k5/5xxQK/zUOV4TL4
Zv96jb/XyccvPm+2PPhJX9S9nPS+xFfSrsYwOZab3g1ux9tKnN39HbL56PBVL+SN
mIoEPJA05Ip0Df5bq/pzg/QTtH7QsfYpC3cEQYYy0UhUhUMb37V0zRPRiWX5T9CU
zA/UBO+uokm6DruiYQ2nfrphBCJVuXMTZf2S/4J/X6givr3TKLFmekctbjqETt7Y
OBkG37rADA352TuliAh+0qHLLZhM+498c6OOJu8ZfWfxTTRzdr5YovZk6WQwUEFw
hFCMqttSLLN3MvtP8hBmb5LP1EKw9VS5LhnojLoQqXmm/n7RIyFkCiHYXhR4vkwt
weMDW3jxAIyMtUTP+QLAzOcz0fLxk1h7NDUMC/wAnJyVS5JxUkqlbyLWSoYcRzkX
Ue6vAOz7ppmacGouWTFb93C3FAwpY2wkrK4Vn/u/aoKu0N3xY+DfdTYKyvZ35tdP
OVN265OPqU4Q3QSV0FNEItyCIhc3TNvh8CK3LiQGQWeFWXUm73s8eJNNt9no4dAC
yWbjlmw0/6fOLm/LX1z6dMrt1YM2CUl2Ly6bPtUUbmA1qVsol5OeSUTnhzj/Wy45
9DsXp0IWxw2mOHfr5UazN9gz1+ZbE1FQJVk4OCOLrI35f/IEti7h6L8oxcRGi2ZY
gqzRuphnEh1842Kw2G1wapExedE3doiZWcMYwsdaOGpZuSmnLW7fJSUK4TcCYIrM
NHxf7vbXXov8dEd8RdnDpAhu6kHLsQz4PBQfnntlfdzMZkg0FovTP/3+38cYLkwL
PZmTc1wTLMASKzT00EI4/uoOW28bWl+FyGGHC5GnMQpkLuY6i7PnJ6kiPivwieWx
29MR/FuOADeTSdCAvaHfiYLBiL5EIHGpqCy5FeYSI3hwnV2Wc8GvykMHZRkrNPOe
jj+tMv5Bl58WjekWecO+hvAYeWMakK9oTdyAoGGZQ3JaqqOV/xpS+6nWhTjSUV83
pigZCocb3voBv0CX2Q8lD+kxz9VWPLtR7GfZ5Jw47g9qXpilJ06gXSgreQwQAszJ
YkNSFWluA+/fjg5WiDHvW7pIw/UPTgEkQUZVMfiAEeB2BHf9pMpqbuYHs4NmRN50
qC1O3lLvU9rajRcTcUzoV2/uZyRW1AfB1V7Ea+CkxKLgCAE0sTPJ1J5PW8iwCVrR
ApbtoyGD5tzPLBi2vyYa/qJPG7r0t/mdH7thgsZc5Nzce0L2MzCrIwb4wd3tMFrU
4BGBic1adVcyI3KUoLDIrci0IxjICfsyUNwIhusxObDEwGHhogtTf7lSfInPhLX/
iLoMoe7AvlviZWsPn4MK0Q25zNJBBYeYK3qb68lWFhwIS0mTRGXoLvBO/KcCnJks
v0aE6OoDxGYcvlLChuPWXaOzAh/SR1AO50n7qydATo7CH+S3VbJr2zUxVAOAsxfk
gGim52WrTt5cDiXSyDCVVBLfklS5VKIkhMaW2p3fMZoz8nVD8mhZcVjotZSYd6Cz
0SMHihTkece9qAbS7CEhyZ5crORxmSZlpqXdYfRjg3+rvLkDCLM31EgDTVJNlOkQ
7XMbU5NeDHKmnabJ/622CkfUfsZdvOJbjRprXsrti3XGb9hyrKKxJ5gYvk1teKyQ
K1m7nMqxJr5js4A9+iXedBTuVUZ2FWw3N0BtH3pXCpPGlBL+k+IiW6pZ9U4lV0Q9
ulYnm+ixJWCL20dzviQmDzftCv1g7mhgVMm7bR30EsYiepASenKjTfmWoSFBKAIz
rrgL/igjVbcoJhIWHTDq2ONa1P2OL3uixFQhNs68vjHBXzqWvDb4kplsOE/kA2PJ
K4Kh5Faw5d5dnnG8RJ0cQ+sdGF38vjhy32hXihPYbSusaOuW6LrcJwchPSHKqPk6
cpeiCWurFRVBtq8neIx9S1xSnm8CF0O8Mpy24SYK8+BwUwjGghCU38d+WrJUPZTm
AoiX+7vXB08EUYYjmZMtAtQkszBbiKponDh2zPC9Yohe/DYh4ShAG++4g4aCbNhr
4dDPXxGqb+CFRCTx4AtnCD7NA9bJnZb+zFlWKKjDLlrTDemyDiyDF03iyDpo7OcX
iPwzqQNzBlsIUcjp9dITDVE6yGAJbaebh41Tdd71huOJmO2G9HtZBjI8yqU8OMwJ
gtzwVQqu0xRUA4KQ8XdOCpVdePwesTlwyC9+yUdRx+yxwfaEFBTLkrszsAiF/msU
uWtoCK9543LATS12nPkVhS1btESTQB66emKNIs0fapXjIYG+LvWPQ64lOvFrGzf1
T6eIteAVyJeO1bzX8It3ZpR0k0cJzKhumyu+HumxA/A3Aki3jDFPqPtLKxpnIfWl
QfVphUdXIPmR4XTNFVO6jWqSE3k/j/+gv8w2f4Xjxej27ZakdEbJsJkYc2rS+eg7
rzFAA2dC14+pEFLJ1GM3FYCEV5IL96C0gqSprwrgUzLxxVusSiQjKT8fiYEWd5YW
3WJ3PQFZKS2icMOF4uoMRojnsWjUt2kq90heq+FkR7R9tJiu+bfdNAsui1CkFUbc
k/H/p0wRrvI4DMikCR7Kr4pAJc6dNnRYADPqKzm9uNRR1znDhe6vKyz/OcpfgKTF
9t3DvxdAr5qxt8Iqvxv0Am1e6yu3LudhKcezRBnptsoUoQylHtJxlMiNYuO6o8XC
JA8cHqsnOBUeZq3mfJQzbPK/dJrJMC/OLhAA0S7EKQTLgWIjRkw+F8Vzyj2gaS5K
pfjkq1XM/2EFbt1u8EWDuqy6sH/PXHnPV2biK4lNC2eLaXPTVYiIpK43nnjUaZxs
TPEqc4qiFmr41Ok5f2ULkXIkVMwFqvrGihAJL+QPYZMwzTuu7+LOcwFBMc2RjcB4
aQ6p/S19/Q12xKthbJRcvinHO7DpG/uBWuF9MXXLkeem9gqp17z/Chbn91VentJJ
LF6giLqBJ3VgOQ3r9Hyf2DgPDOKioSv1Wu/zRQ3kX5vHap27UmwuZ2nVVqC6qcTe
J3bF631zqLaCvl0R165BnmLfSTMDEXQbELFFV1FfUYdhzhwUTcopdZvG4FoBmA84
xziXhaPdMb8NogADADflE6zWrZk0pQACU8D3cTxnNcf2/2jAfConinrY8qM2ekRz
RtBwaQ8bGAY4qk2vTi4WaBdxRB90q6PD9EFltMHyJuwK5zrkQziocUvtZUW8H3UL
lqLXH8Tn9MgSYBqpBSpIcCDrMrjyShbhU6QyCtdCJmTKbr/9xQAtzrzE8uzxa4f+
5Y68OQBFR7ZXz/95b7HvEMJKbdHVi/+sy1d0B8zlummvBmZOuwy81xeEF0q0+wrK
t6oUq/Y4pIfaC3HS7NQteCSYfwfuRPj4tSPYwgCxBZ93b4ARDwpsF5horlqJATTM
+s+1WbZZHykFVlfjAa3HNDYEc5p0Vz2bUQg1M8bWRhRFqrk6FbBkeGxM9XXMihmx
bT6Iz9dnh9wHNFraRAhNVgtSFH+oCK0b0cPMp8O2prLmJgSi+y/4CIn1Q8nEx+rP
dOsja28umdhFhtkKm94OfK4rkhuJYNMvAB1NHCDIb7U5zLS4AZHVarvHQqvS5Z1w
9tOSVoladMAyzCK/Qw7cauzqyW0wwWVewZk8SJrsXi61+X5qiJje2pdn4FdgYxym
HlebW1PRQEqvC9/RiXTHKcpPtYOHq+H2tEiedHAahmAbdIooFa4saCuHw/Ux2T4P
bzXa0GnCCuDsj3XQE2qofU9cgvpCXFlvOY4dqDkunuFtWnLdH2kBU0vxFHpM0UtQ
NS8k6cJv5cPiJf6T3O9a5W9327FGJqrGDIHJ11hVaIRsxKVauJ7js7+aLtSK6Gfj
vum5ZnKfW1xBPndxwiNelVJXYzNeU1ZLehreV/3Gx9UaVRj5PgNaL15hDs6mu1FU
YQDSfttI0kUDwfMERhER7JPER5VGP4IxlecFXPArOQULLFQobit4pkFPVR6NGLHr
WkInvADdrku2O4DhgvszriTc+gBXxx9JMDTiwjZAHWuo3B6HstofM/Q+jWVbu9Ak
eOAx2Zls6xzo1PdzqGDkuzjiJJEsalp0uKZr3Yu/sQwPd9OOLqgjCqrUajMsxpSE
Y3GXgr7eoTZnKUL+WDgXVnaE6MfX12ujk6htBhdNik+6Ltqi480kQ6DsCE7enoom
B8sVBHniB89u+gDAXbKE5Ri6IxATXKLjAA9gt5RSn3WUCylgBwl1qBl+qccz4/xt
hDnHv+ToFJhMvx2tvagr1Ib4DsNFIBWfnoCO1Gm7XiTxwQSe5IlKFCldjXVJL3e4
OmpkYyxxdgCgZLKOjFrpo4MnbrMUf9TBM+UnCrjl7vM++Va/REW0UMb3Gt9Duq2E
orMY5K8iP/1CrMQp5hCD+GGT7OVytVjMLPB7sRHu5QUoIUjonaX3tCDracA1C1Jx
xSeRS3LmEJZOOe85QpduuvIfXtpYwywOBBWMk0uBirLP8ZBJoLVN9q3NfixXLfJB
9bF14mcciW1SgaRP0U/ux7MQ1JdfpWvHMsHye86bS0HL9CTYDsYNz0RXyr760Z/+
iAhlFIrf3dV8dFb8hS4UD+G6dUwJ45sYsidKCVhHF+dzSJYYApFPK1DVz0rvn0Xc
rAE+s/ZfX/hPzmuIYWSjENsajGoqh+A/T1RlFJiGcvlZbPttyCSnjjBQwYn0vkSK
Zx55eijsRCpMoCrQjqm7V23PYRVUE6T7NttopBqjJ+zN3TMgL15+ClY4jNz1Ud7F
YYyq4i5csxsrwFJRMRLhnLfhraIaqJLZzEKUr/10IeSpWBocLaYSYifFUkfkr1je
nuaLg1sZSIlMyVEOui/ossuEIEUrfEQfQCgDwbHQPBTNNaU5710+F5oOaNm89nyu
2iWrTfhGyrdNHx7M4iXmFrJC7RtSokkyuo9RbO4Jpd0NCCwZJ37YrNVu9ZE8CJl2
iublWwYYbtNYoc2eAKnUgs/cwpFSEHmmvkzJnT2vIHo9D3Vafwvega2qErBiMv7D
1fskW6manKv6MI5QaoD3SFD92mla8DjpgdaxRr5b7Tvp3t/qWtGZ3SHVPfvntyzr
6EGUdJd3lZQq+qf5cvw+T9JINQoeYlIAk+deG8YzbQDoE599OzjWtlIcuIm2q2E6
gVl0AqOV4iRgnhtagDfnWgfZZYjf02Sbl++sSfcAC7kVNg07/7MutAwji0Rl8ILP
vXbH4tihsOUcHHkdweZhpZkHhlDMHEmXyxxm0Zowjl8oDqqezCAdCBNIG16nByvR
PQhLZtNB+CSrI2z63ePgqG7kcaHy4NQjpoMIXDAOlu32ajbKpjl1UHdiukhAG+fk
VGCgwHkvfJE23zhB+2b38rs/arCLvf1Ef1lzbAWQF2aba+30o6u++lnVrdkV8CYi
5t66mbobR5B0VHCyTm9GMaoFip5FFIG9uFFtftxddDdGxDb7uoMIh6DXTpJF6tM6
HlDIbDmzBjZA9qtb7jyLlI6PQJnL4xJFNOVssqd/xrun+yPIbXXJsnVxuYHHdRrZ
k/EbnES9U1m7SAMTHX376ng5yTAcQA3YZPqjclAIpJod0YFzq5XpVcmwnvRHwpUe
i0x5smO719sIbr7YuzUspahaT/VpJYPJqRs2ouaSkAHrWPKYRkn+ZIKECr1CtcKF
xpeRcM6b4gzbS9ZavRQUKX/pu49arNxbSNe7PLzEh+QGAuqfbJbsnCxvjGowYKOJ
KTujpLEEh5RtJIzkSo2Hy8+IHJ/XDOrEcCR4Hyll45y/OHMv0S6/33wEozAiV1r/
rz32XiLySV0p7npcrra710u6sLvfXmbFUC1fcwbkk1pYfqMdc8cBNeyIl+UdpAOc
6KCjfDiQRooIgk/9tWLVz6Ga1Ymv+6EJtXt26NsLWmCtduqtzbBn79gg+xbZpGML
GHzrAWa1YdMwKha9mr1agrGGCMpCHwTGdrHLomxurNnSkEzr/i9orNiivoCJU9zH
mLly0tXPwoee2cLQa07pT5rAw6CSAUvA2dX02nAjmFp+pTM3S86E/kiafvLXSylC
1I0jWEArwwWMytPAPf4l8GsJjDANQn4G8CaSaqTVkah6ev0pN1MQwW5J4L9px3eW
PA6NYXX9A1LG98CKOG8A8dMTcoAMGy7BKvy++e1MyuWkMtOB84AkjnOjBPsDfoX8
jFjfJusqlBezOszWkRDqOnb13Vhn2bZ7aTIaNgZBkM4MXnU8riTfoRtmdSH0rSuH
ICak2jPaxPWbktNkBwmaQ3CMNdhaRRxkjpCzNlm70qZo+vb0qOyHgQI+JYzB2Bmc
RiHV/4M24zwmOcix1C4oZXY9wja4NDOyuh9SUh9RfFAP4fO0sK3Gn1I65swE4h3E
XfoTtqwjHrFxbYnVX4XYp17nfAxw5C/sZ8N+kPWI9EkXqs0vmwWKIj+ODFqIPYjL
f3PjU94Lrl1oOFV41HF2uA8SMTtVQOsdIzJbfrZe8ZpPLK3QmPD1L8n2wMzPFkbP
2ZQlUGCw5BycM8rMB4thwGb8UVQNB+S6d1dq9QDE1Om3tjw8LKJJzPIFjAvq0dU6
6FVSqEKVppIptMecaDYQJZMicCnXu1F0f3dlMatuvc1BeWonB2+rwbWv/NJNU+S1
Fb+17HpdoKfEmInMvP1YBy6Q6oPU3VivdwvgJUSuVWiUplcRoWjtD6Ev1E9+F+A6
//WBnEXbOnSzXX7i8prx8dgh9dn9+/YY12tmzU+3oYHOuvhBiII2GaGg2kx2Dsu+
vVcjJN/NKdllgn9wBrKBwU/qpXmA16NJiEsZRq2Kd2yLX+9X5J/z148bNYqSJTiv
y/MpOQ9XLjAtSdaAJJiJpBWxvmMswTFip4K2Yjm7odxct9/pY8cXwI/kmfxSE/F4
JItgI57jqSin6s8yQyMOkmrgPg3uNT0undpyRwvcVngSb1IB4tzyBaC76JUQ0u8c
6XW+13OTCx9Sxi+xH7CGxlaSQYyQsQ84TblmLTEPsAOxcO+WqRIYPsrtRp859+ny
VG93BC29C+DJ5dlMmmmAXOob/+NqjNhTliRSWo5DmmTNA1I0FpP0AFakPsZ+gUQa
48l/uNVlg4CMzm+pUmGDaH6nrL4JYpbHgCVLf9fikpUHKtshjyX33iPemnHsSFQq
wTL7bfIheqb5hPYXU0z2lXUP/XplgDFz+LXrh5DwBatOpjjDNBK2IB98Pl9XQv+7
pil+fDqPHFoPSuM9g45WSBjiErbx+nt2VGlAzF62pxHfSSlwPCSC/yYyBYDfjLGb
aVvR+qARpobSYXDG9aMEnLfqqYmnjF0fesW1tskscQ0sIAyA9ZkhhPqIt4RM6pMB
b7oGM5EoW0wtenuoqLwwiSn7Igf2nYsTuECUZ4e+70mEbHcI6CobwxE6HBAANfpw
+xT4qyHbMxHAPMyFasGa91FE0Sx9xjkKeXHUMIBXtWgya9LQBb5nv7nqbYaw0aMP
SLd5gBoGkwwGqAMf8fTF2PXpevIpixwdlnLyJaEtHF+GGlx7Rmk7Lu3DynpT57gT
XjkpNE+KxH+Bwj/ecmVp6GSKqRREz2i10u9q77jUdn+MHtUxhQf59228+yIvyZKI
tzJcoPYY53rtyu3FAbM2o6hPX+94kN3Mb23OWcVNZ1Q1h9yf1ynv5ydVJvTEluR4
7CFhe/Yl1UR5YXkakR4hPWNWBD96NIr8UYacchTQOI1IGE1/m90IRJrgIe4+uhIE
CKjeHnGYfHYz4P2TuryBjjD3KVZU3ztmK295dziIVb0yAMjygxc9oNgW4+n1Ern/
jpxZZKBDIFkmmQtFPsKjdO8NxAuy5YdaBXE/Gkv79K5+TKwdQY1qq5/wOUqp3nCP
DQ8TDk7yEjl57JgnKA5gjS1ZWqBtgffdUut9mGglhJURiSdsmm3yDAl8n0wZIxR6
7ulX4SfVlfV7E7AEca2XIqxnusCOVX1HUS6WcRql4GFCLMHNSojvTGqoiBuu0Og6
4gslNlPYBs8fCM73IUINGkUwT4UDDzywi7DQcXwgoBw8J0/I5Vxn8GTNVUCbJwLv
kl5B7IzlSCXImhFG1cxFhfgSYLTKNGQKjtw2Z+ZME3cwsBCoiqITtFt3WP8vmcJ8
6wHDqsq+F45+jufyBW6PojlG6jMqZ4mbFahQRfkt1F9fLW4Em31sCShXSNPRrDeo
D4JExv/TAbtsll5A2mid/CZ87uLF8wTTnK3NHAfsSvFzV+6EN0jSNK8P3eT7Evyd
e+NXOk8KnmWrAAghzW3BsbLdS8LIGu6jLjB3v4sAJf6jjehoPOdUtXDCzkZOoNar
tOGWZBS5iVOxbjGzD+aWcwHCcchkbc+/qnpcOSFuPKQOGwJTUOptJWNhzFxpcEaa
qAlNuIWa28qBg4vxzSxehYwwUVxHXy/DE/bCz7l6NT1ZCuLwHTs2Msr21xZ4P3y/
Qs4l+j3Uf4N3wrmX/CD58Xft5V8YjIDvnuHECTSOlTcHM0z1+thrBBL41u5F4Hki
6h8xUZPBUpZa7aFqWTEa67IgZEL9hPvL0BLKybm7sJOqNaX4s50MW4lJ6oyz2kgn
AstSKL70RWCglyc9MwTJ2e+RiK8SX/wswoVA696wrfzU3qnpt6584IL+3crCnz8/
jD3Pf5ZcybBMEaoJj0VvFfYcoXMdytO680dkvXgTN68KpzTUscHCh5ETbTJd0J3a
r14T6OdVLHNsgqw2lXCkftwUeu1zxBgpboKQaexC/QHgywtsnzKJjDPBZQZZHFhd
OT1dmc9s3UO4+iiLKUjehhr68Yi3y6cNCjLJ+X7sM/o0qOS6fEtkqoktglpkYnnA
FwA0h5ASy/RPppLWvRMNdtPf/WYB8EmGObHBiDXvU2Qi0psBdl4XuseUQS4CbRGJ
0VqQ6ciOysWcpbPz745XZAd4fm31TN1z72SpdehbM7ef3j5VpAhBfMtcO45EykpH
6qWMzXKgT+4SWX3HBIKpnrOBUEmr5Y37g0GjqDu6lE5C54WlfLZQwIM/XfqJQZEV
1bQhWPIdya9V53mPaI9R/5+L6+W4Yij/JNOYIiL3M0NomZIy5Hf33GNckyA8FQuw
+0zTDmqkgsV2MBurCHzS/bUkv36zMRJB+lxCXbACjt3NZLKB9cVdL8Q94w1c26eC
+3zzrAIEuHyvhC79SLUwvAc1MysUfAiRUrYckd7BKpSPf5HTPndLPNSKHQjEWUFI
ic2OxsfDRbIlD3i90RYoE4+5a4R3I3vIS1dHsclQ9li6gF+fZnzvRGGHfFdrDGBn
IlMb6kIOjvDATxoTMa6bbhpIZ0SxgX/c7y4sft+EO4NHNkUqUk0YM7Mentnedk7/
iQxHZE6O/yQAeJo+G6cOShqzX213WnBm9O+uYmOCME6cCUdllUkeDkYPJ5CKSzYQ
9jpKgMPlMvbznS4sZ7I79mHflkYmkiUwhgIjb1QnXdUk++l/NbzVaFZkDrw7qjlu
5FZ5/2dKK6rd8xTTNP0j7H44RBn9zCNiM4VLMLdYvTzmJ37DY2eqaGvGMo6OBGsm
TlUXevUYB9dCFNn/OwRPyjJNjzhG+RXZ6dJYdxIvGnBTOLEckQF3ek6pRzl6Y7uQ
tXGK0wh8o6ASa5wCRxNwwbuKqluea4J7VDiZs/vUKPTn5/4WAIe+hQUAPEZsVyvq
D0aSutuuKsirEewaxYxUJil+Htj3HdMmjR0n7YRAVCdOYe7R5UI4TXNGAbs5JY8x
PVz9GaiVDHl/xe03JIyZj7giXVbFCWVv+s0pagNKlY2UhtSprrGCp80aZ/x2wefy
ISxTi38K1WvPc33hTZDQbtUb0Xbcq0PdEJgPa5Q7mRj+0AjmWsr3KUjkakPwoz6z
p24y0M6ytrp/rr8H31Cka7KTc/hYibdmHl09tPIGxHo5v05hdvcjTxeCi8VXKRz8
9YXz+/O4UAqp0vy385qXc/rBlrX1iP3yDukfZ3oXhD7Bj8AhMUuVAotxDtdju3CU
IZD/5h2oyfFxIIdtOcKHPVJJVso7BPpQxzjr3fPb4PpYVj1XpALACasvSSrkkJ4W
8aOfT8x5E4iTvl6XNg3bvvtiIvk2IPa5tnBubBCND5+RkqJma7mZchJ9XExzTjAz
N1bd/iJVjPI8AsFqtBkJ6s9vGbUt523l9Zk8AefsUo/YPuNp+TYB6DQf4d60jC9k
/77PYIeRBDY6HZrrbwJcxazigKRHBoSpEZ6ReG3SbXwJbtzBrR1UzOkX/coLawqs
At9WLlOzObBI5fv8tnceNvbsXw2MQwyo/rnujl8C3ZqqViKUOgGbuFTcDtIFCL1b
8X4NuD9GZyN4RRBx7gxJpyMK6vpp6O90R2NSeRsKYNtkJuOKGb2uzHrvjcI9GBeg
ac/SWljER+U1rj7hcfVg5Dg5cRegR1u3sHtY5vg8dtShECGNsqphAY3fDKwdCGnR
RukrGQcVvvHn2bgMt87xZrqmmYyivV0ZjobkhHD0vq5V+X8ho4qIMEtNcujTuc4f
1mU4kYumJPhl/hVfkzQfYlZFQ06y4Ne8GZt97f97yqzyv2bWjydhFR7tmd718Czm
rRJ1gHLe+JD73WpFUntIi2e4+Z79tYw1DL8KnyAVcAaYKnXBCBTbr7hX6wd4hMjf
3buv4My4DCX34Nftznnu9Lw4NXUn+jpOSB4AcpO3fivwzxsQEmE1FQaFVDoDTxGX
dRzht9FWeLjKQUh5TqMneaVSTvQYplbAsgffQFX6lCjwi46bdKyKozfavjwMUJSc
Sy0VTvvleII8Z/B4Z/lrCFf9IdxnrifVMxD3hfjFrVUkMhqdInFSKXo9Bk6/HF/S
RgUx4JCMrCsreumsOnX6xpQ3uUSoYMZuW0Dw+uFKRr1aqRLZUaBzfplc0bFfVtbm
GIwPa78MLQp+bTN5QkDYJtEFeb63qzS2sGPvOa/0V06mhtjOBqDkSkPW2Z+XvVVf
IyKsQw8/0BFfiZ57WzDGryiDeKZH08CX/MCUn18bitM01fu8s0d7X5vEzJT9fNYQ
65rawO0W3DDuwgHmVt3wAEnYv9PMs5Gg9uXxx1aq8eHJxRB2F+Wt5M8O8rbIWE4o
Qhkh+LHhwfaZGS7XEJfieCiLRz38+KTR1KnITVDI0kPQfaleFealKobFBcS+CtHA
CCBs/8eFzhWlBRMyC0vt55xwDX9pOKPKrgHmAxplOVTUQrKz7EJ+Ik6zma9PfJYR
yUFFMCyDIPWEFjCyeoyB3O6teq9jGqUVPptofl0WPG56QzIrkviOS9XdcspK/rZp
pndreNPral8s5Ugx4hV3tSw9HzXsOQVPM3r7EShP1mcIqUU8p6hI/piI/aO5GQtC
k5RvfWvTZ2h4n/eicfEUCyldf5pdYMgledrKBiFw0IXEuTcpar/92OoYWeKRqFZi
zpcoAkhYl5n8iEPvJl8wIX5L/RUXVCO7EvE8p7AXmw7hkJ5GLXdRv5VO+Cxn/aoo
fSqZcw13T3tVJijg7iE9pOzmciegWXz3N+N3wg9/JH/0kezIzeHebFmY12LL+1Bw
1ZkJP0L56fLzw7IDVv5RHdhNBaEZBVsqPEXWP955AUOkBK0cye38EJCwPNqaPWVJ
29f9sLM0/k46a4QLtwhSIhB47/tMWLm8lcIjfdSP/pfjLgwifwYzE2dJMo7raFMG
cD2Ia+V98nCil2e/xVW38Gh5OPY20M8j0pxulEaKHSuZNIaRBDMMgPvGmO69vbH/
62KpmiMF8lVznqiVoUU9H5vsWOqGIbQdm/jmlWexTAP5W2pAMCFkwspFVcRE6vFj
76/VfD1E77dVh0i0mKmBYF6NiaESLeR0xSEoNvVWik/4Qvg7TI1lQgi9p+Iz+Oky
DBij6zshs/iRmE+qALpghHJ5AnBr38nJ1QzFcLfcrlQVtwuHFgDVBN8d5d1wgou7
7LWTeg9mU2VPphAiE9CnnuIeZlfI3FRtXw4VUZOhZQj3NnnU4IOljirtYgDkZjhV
BJO/HGh+fE1wMFbof7cd3gQCdmtvE+dYPqe1tSEALL6PFwevDF8l7aJjeSVz3aoo
zSX9mtLr67AWqj7j/QphePp5stuWfKMDFfWjCV95/2RtPymbmFqyMz2SyF2nXb7j
UMA3wcwnFRfqmnnEJcBDSBwvwxvLi4cv46bS6q4wczjHipOitIOjQ7BilWG8HoJA
ZbscGtd5lVQek96XhxIa0ED52WfWbohdfC6TvpLT5YkDHSfpkaSYSIYrbiAfC/T6
Dcttt7XhscuPBwSiSfG+lbuJDPZNErN7gPcbg8o2pSqhXv5FZZyQ2ns0uHN7olwV
H9nmXXyCGssEMj+J06kSio103haKjvn3L3FATrjO33PZ33tppY8IIUf2naU3Ip8q
7leU1M74+pLKm7o3AmUVT6DIR8U0xw66Q3mZ3+PICFm7TrsY7irs2DR6CHzwDXJK
2vzGupCvTG4lsugGdy1yeGpTtep9+x1Ww6Z+ZByrgd37xGwnBaNB9aS5ZSXw3hIi
cDWwXSyLZZDx97CAuIW6A978g361t8lfrPOdCGj1LNLEeJSFkp0LPAZfJy7fGYWk
+21MJOwVdmJZiroH9Tmp4eVY/By9blk779IWY+6aTD5k+ulszogVvGsRgE0UjOI3
ePSQhkaFU2BL4eXplWj7XHZ+h1G2cWuwU8OokbYvETEplT4aXpuCUEGjp2+rd7L7
gDwad/NXGAjDXBZqsn9+b5h5Fpj9bAd4SPEuYXoFkehp+6Xb6t2A+3Jh1ErOeJGn
EZacLlPfkJ00yEUg87LmkUOnQng4LaZ3axD+AzC/nTtzRZYJfuJmU9zKrC0Bxpuc
aOBXSEPmIBcNTT4xtoJIZya+OCa/VfkkvAVfIEFdDIrLDFNwdsiI4+52NC3RnoN0
Aopjqv/sAoMf+jfPsY1YL0biqfcB31pfp6g8F+QMtOkDIc586fhopi52yeh6cdb1
FLHQBSqPqJcy7uuXA1y81y9oF1FvohrlFdjFJQdE5jhL98blXx6v4mjCjI4bots9
OQSjP8MA7dZR98asQ2Y6CuiFpvohWd5sNgP0AZiEm0hnE+vRhYqQv9DOBYf5iBtA
2qqGJiVTHPR9WQCOU4UwkkwAAI8xqBvEsLLfj4DoD7wYrltppbTupcggPRl1vRTq
B/U8DdzRTgNGgXlVgABEeMlth7qwRyxUr45erIJWX+uqZmrf+qLDZLm42Os+c1Ns
rnuqtvKLjgbf9yi6ioZaUUuxOSjguBkCOKc/LHN5cHTx+A/WKxSHWVtiHBhLCM15
eBv6Bq6zEiJibzIiT1Pv2ZO/vJLmF/ETEC2iPo3kuvDl6SY8X43tf5/sFX7s1dtk
9+oH+216S1VlCWC0A+jnkg1IvgIurDVg2GlxuA8UlJMyhS3G201cW76R/y85C+qF
rHBxcCcCzF9Eg91n5nvP/NFcFEkB68g/JFcZ8LHlmD59UJana1dGLGX4VigmoixU
lSFwvfCx5MIw7xVIeOuFcal04L6ssfiEFUA3jDawiLH9y+lltyRJfpVzwBxe9hVP
UPy2HSvGNaSjATBcThmcnFhk807aa9umcAN38OEtwOMiLc0lLZpk/3E9f7BGjD4E
yCaqqiSv10meoRKF1RuG3MDz1Ztt1zx1xSvwHK3qS6dBfDYNNdS+sojmDEKf1tUA
0imqwOG4X+BOI6hi99ZahluKIWMbHNLgDrU8l2Aw28nwZUlLqGYESwoZsyJCclGk
rh3T41c1CBEUMMP9ZOFVwwsUTlsHimyFWNTNdCJh/86VRckyyQnV2ERR33/yBXLa
36DRaInOJjhgIMiL0xHjp2Vsk3KYEDY2JppLsReaWiVPOI5q/mm/hwUqg7O+D6kv
hlvLnCD76JcmSJBAYEuG49mnKQ7Bfx4nMmL/7DOBCkbPIJLptUqmu9Pv1P1ueZMs
QxfCOyRb6xiQmBwPnvVhWhyncIbP5dGi6XngS8V/bdI+O0eWEMKlsF1z17WuPa7Y
Jjow3NE46PlED1yh8DycjT5DzlIMiyFQUJyegqiVODD/aRVjqB2njKkHTg48ped+
e7O3/ZHYKKm0lFCouNnEO2lnneDQVUY7vu+sLIEiQW3NsW48ec98oruBiCGorX/n
GEO9SdsKgOrig+JxXj6j+3LbPTp6lVMqvGV4zr0KlTh8tXc1O3X+DZSOzaBtcvgk
j1gAafGufCkTUsXW5bV/USvV9fGPKpR3BuhUJsPR2xH+oqPjl5OrXnIiga4gsrUu
ih54gX2xTZeHAS+Z6+IkqaPi10JunqRs4SJ3Fvt3PS5Sie4/DhMc/QSdegDtC+UB
xpoLe8Hpk89oS4HJCb4LweXT8CxOmq826KOBDSfaLHYTuh+4Z+JZSw5eLxoYUpl7
bKM7ecKqO9tsi8zGFC319tY2+W5VETbnBNHyfGox5Tpkl/m7UxaW9yNdMHLBfXrH
FBfJ+P1CGfuHvxJ84CtpLKDhutajnvDgOTM4YxKNodAnrpiyGo4tv6rIXOROKXIl
0Itfg0a9s0RvYautpPyU0Bow+1dPiAjl0wISrSr1Bzok2EhxP+7WFMMxcUOwzIjB
UZqf/oYQkiaEurf6fUKfneFinFPcoIVO/pEQkiPZh4QjcYD+zxGjyAWCNlBaxOgm
611lBGhWu0P/bjinzCo4N0iwxE4nfhoxcB94F4aLiHznaZvdffIxTcgL5XCvvFm1
orhHvRcWR5e4bU1gu04pvJ+McEGLwzXQR8YUDkIEXAqPCOJfip0rLOL6HoWpj2CR
T6sE39/xL0yt1msityq4I/2rD/cslzQg59Vu8IFiyNgxPNcB0AXtfBorOIe2XoMf
nSHHVUgBx0w6WvZet7m/ZGPJhWx1zd3UjP4f4vOv9Hwi09Euq9OgOn7r26nbauPu
VwXguyk2e70Qe5fiTK6pHqyZ5hMBmssaX/xSFsYaS1WpdIQDeBYc1h8ZhjqAz898
BBHhvrbbSJ0uyZbBY2jfyxL3xzajA0fdZamQ5lnpWtNLf63zyAHnD0oQR353XtAI
vIWL8ZAHfByuCMwkLv9GAVWcxbBMX7oFGC0xOrRZ4dHYIAYv4l3heX5Af750+sHL
54S5Ils3luBuZ+joroAfzLfGYtUOsbCwC25bjx3cQR1RFd8RTV9dOmbkd73LFCc8
aKXsNeKZGWaaBTBkzmyrx0p+rJA/COEwDJoFG5aceM5cr8KxirQv0KN1QT9w1wHI
XRZxRCPBz4q/EA8jvMZL1dvhx61IqhNd1K9kBiUlr85Q2ei93JpPaRKn9MSv/6Qj
JetO4ynr67Vha5w5yt2B7X2+sbWQvBRCwh8VoElIbERt/xY6fGSZJd/2hFV9tRem
AnlmgUMyLBOJSAr5SEKaKZHM+MAkNL9lDUV8GW1cXvZ43CHeLYwoliFJyyC4Z9lS
2GJXhIQVTHpE6c50TtdcDIi4gkSOh+nnWVYjgketjmJ+/J2h8mR4jbg9UtsXzuPv
9oVcxxSF9v2J6tVM2aAR4y0E9gtf0QMIdzHiNlIQUHvr6tXwvTFlzXVlyfatrspd
ocZy3XtFx6tv5wKZ15axgblL3dcuPDw4Wsm+qPpRoVvMx7pO986fUkxAkNnGuczo
+V15qi+Kky6cocooi1ySYqWMgS88P+YeOFDi+zejMhum/GClMqMlI4hipde80EUM
kdoeHnXRjrYkkjNaB0VqgjVdsAuhIMxZ2Nhc2i4UY9IzQoZozX6k5+iHmblmuHri
1cWmitKVr9AQExEEnKdAOozNcSF3a6qpSCv8yE82bWqJ8nkaoa5Pi61FpinKUQpR
ALSgdmiaNUZgErEIWtVe4Yy0KBQ+EWRUuuhcWqFGWg8alIhNoW/QGab+pTBhw2ml
nHcyZijrUlMtST8TfA27Qz+NH3tlfp39VafZ0wmMwL+XKYwsnd4xS3vUETwZG3Z6
6xGk43UeXOdxfxgK+2t8a5Qog3ChlE++ofbJEaJscxRavHBYozMICnbixrIWDtSw
QBijWqYxjVXHk5lqaUVK4zrZLaEjAFP9Mo4PgKaONI7yPhsgl5G0mVZeE2kU4WGQ
PCJH8aqE1C96k6g2nZWuH8XzV/osOe67GazkaafD6h+rI4u8XNMgUcH7METMNBxb
P1XgtrI4mDfs+8SHmqJy+G5WrJfOIyzO8CLLAYjLOHY1nrOXDqcIl9eRKr9AJ8b4
XdA0Yf+KDkyio+SMJQJWXOnj4YkeotjrH6Mdz99feONZjaeEdMavXCESW2LjlH8e
wpA27NbyV+OJSjIpMy9t57sTcLl5pPtXV5s7bHXiJ9JBvfAVXq1eAxs3AaNghRZX
JUn8tn3sRAcumxE16xqJj46gumpqKWEFc6ZODl38Ybu06Ahk8xQviRMub7mFmm8F
D/XfW5TmCwcSGltFlsgrbZfTyZriFqlydsiySGeHdP1rOAVsgDxCN4OYYAqyY96X
Awycw85IS9mbM7EamUTvUdQtSxIxcxaUUj6EYbkSGw4wiw/jtMMV9/86rlAYlFbl
w+uwrQa7MG/jEefzequ9SBL4Bv1bQEMyTnhajNgBVAUPPGWwqEHYJXbL/JiLzWC4
zCtIkHr+l/d/KlCBvRkiFHbtZaTMQags4kAg02nViwP9sVO8/n8OjbtMykpcG6yy
An1DN/CQivDwLbSzQQBVaT7YLHreDDXlv82jlkntZ5jGk5yPBSd7wpp/M/76psSQ
sJ9+I1XGBmC+S8yobFH6eY1irfwfs9FYd2NtW8hhaBIQciZ7HVpaU4Tkg74KAHVu
h4jSTS4Q9eXjoylzeVpsNif1IrBAf787l2M8RI08B14otnn0uj8c96m05RTcyoJH
v5oO5S8rFGNG+zKf8Iuu9cWoRoJJGvMP1GcFY8OBAwWMKpw21ZqhwsnUIEzS1aOM
kd8d4iz4pWMH/Z5PCB9k864GWyWzanAKl8AHUIPoKyVfhAEVO2Y+g/xqN5DWoxRz
TRauEtteQCDFdWTc99KZ3CBkbgJvoby04YjFphEqzeI11PD0nrnYJNGdoqAWZVif
PpJKuObstH0qfJl0tc/FnzxLN9fPmdEoErZJDO15AG8qWERQMIlsf6IjdlfN2T1e
2Z0FtSs/VfxxgfRR+Xz2zyCbaFTfyKsRABUSx4JHrrCo4eg4tjQHQ4HSYPSQLKSG
upGfEijKD5Csdmix+eLifI+rj6j6jJ7/T3kBarCY0II3JISmpCA7k8hfR4svgKPr
xr2xckZyrrL44hMQ4XOdiJPw0JhMn+UrmlHYedHshCz7Pz2i4vtY4O3TiuETdA/y
sWNhbaluIF6qB0F5ho6CB1hXy/XX/LGIKm9SsSV92Vay6sDq0HYYknVOwhO8MrGt
+kuJHEBGHxXMPk0DFGwmq805FGC4urD65hpMrD9+ZaNo8sxbOaW3StiII0QxV6m+
xpWawqCurxT+mlU7OVQ7yedYbmSyIzgiwizf7/qYltwV6nT5zwxs3o1V62bjAwhi
l+GATwLZUDfrrEhET2EhQR4vp6VRvUNpSQGcde3c4AdvSUIuuOwgFKzXAdgzGIDr
z3Fj8KBkUELmMJWEwVCHWSlpmJAYG199EebUypss2AjexqYNitqC4wQG+nVfMErO
RzWy5IXScPZ7kWxBT/9X1FoHmrteo0m7PTwHaO+SL+x/1qTQyIT67mUgIPf7o+hM
3OQUJwpQzxjX1fxIyRvUBe6fE3+gaFka1Amxl+W6VqJdQCsx2hs4RF4lyd1V7yjz
5+JfHztHn+APDVdO7dYf1Ms1a+iOuPqe0UcUSs04xPLSsS113Ce7srvKIEMNBqt8
i3zOUbFCeg3xWjSRFsnLrnLaJNSGv2t7bbncW4yLadyRnyATCw2vwgeL7M7gl9CL
OZH7RRWKZT0z+jKjQwNvOiOtIwlFFedi9v+gnNXCjWWQNNl6zZFpn50k1tYEXfl4
lSy/w7/HUezaNKJ9QvBnf9O3Pclpp37mejgWqipS2rRBvF0LGk9molDm9x9G9yzJ
aPheW6Hd+uJMZuBaTimi4rahOSMjMQS/Gf7Zy2Von6CcpWakIIUSfVORsQBq61Zk
jgQUTcOYYVLB3KiXSuEPiY+yZSaYVy1qwDOxHUq/5J4jKBntmv35M3+/1vI135uW
MFXNPGzEM2Zo8H8KDdXaeIVh2dPlZ0EjuSLgZgsze2fgEo0cgn+/JLORkg0IEuZI
PQlM/jdSaN45Q0edJSnqCHsnde/zwKCZkWnHPo4EyKapNnBlaWMOO9gYzVrSUalg
duh3zYU4OL2B8Cr16zE3Djop5N3yd7v7Hl6rIHnyAbL0OV0JtFlZ/eOTspFOyuaq
v5TCQEwxUAwLkEFGwMqgeZDxHGVwTrALs580b6fLqqk0Zxlm2y+H2kezmU6LJTNN
PClVF/uugU9FtEaXssROYtIqotwaqUvvragV8cpWlQjN5SE+fqzQEgeI/xV7pkB0
w5QiK0ObeNbDSmw2q30l2a1f9T3mNgaZKG0KVAiynB5fbg21u1yMK9tvOF/madbT
7Hjo2zGmaBx7v4ek8vFUCqdRJQNix66qWR/BBDNR6ko5LMz7b0Yyno8v1Y+bUgRn
3g/sfO+Oxrg5cpd6qRzIK5MGZe4Pc+lvT4a0xeq4Nduq2g7QHctXvQwnVCSeDVkI
Vy2dX/Pcf8dgxNkIIckiGQPcRsnBaSYzUGooIP790Y/q1PU5zzCMqO7KQDo/mFc5
G+lK0gOe+QFtqNkZKUCld7s1YQwDhMQqwIpd3bKqTugVNWFPstJvyMQ1oqYzUmCv
s89dLQQpDY71MRu7gJGMCDFu0T/k52WpF4fYauLqYjBWzPg1c73AhtFEP/fPqQkJ
pu8JIaCUJHqPAekbkM9kiV2A7YfetwemBKWD4saM9pxcnG+Nid5t/U4LSm2sGHO9
kxHouYwep9nRwsmEScT0gi2F7xq0uuD1wZz73zAlc3ABU7fqpSRJpvS6lKNofBYp
yQaYCfxiSQ9unXYJ4EmBrdMjZa2Y17AgRYnYuc71kaVQsNhYQmX/1EDG2N40QsJ1
GXFk6Z0/ZEsJbJNqnTYysJRj1axqs0xLyfP/uCz4ADNx3Kmp8iFrgzj2njTXXKYd
HO1VuBkTc57A7itrIMe6Iw46yndUlRK5AcNb8Kuyo4GlGFu9Oj1KXwteIzfBLkhc
3AuM2gD8cRy2Rv+FdDk8Yz95/YGc8r+gPERQTyBJpo6ZolQ+I57jzhdmWMjRgpnc
ptGPFjL2ZGZMLP5MNezdVB81LUB2xaUJ1yMm2szOB/6SbvMkIOsWop23OGf5aQdG
GNdubXAp9TXJRthVwTFVaYHogP6Ype0NDRIH4VlWxJabvooocH/ZyclIbfKFcIDJ
1B2RXQd7VoJHY4jJn5RFC66fIflkni+qnbLKvl6rLfR2H7NgpahfvZ9GxzHRB4Wa
Xnw2iVnNKot4h1GEChue8h9XmeoUV77mdCdm4kIlRiGxNQc7NjxdOU82xCcsQY1J
uVklT/OpgH8yUQiLXWMjwCYCYm37cuc0S+iYvmcdznPL/vlllT/+g76n0mMVofLW
n/OeuOLfgXgTQQ1BqyJl2sQ1WDubtDMNosVtdKgJ5YBoJHgWMO+u+VFj1nc3QVJ2
ZCc7gQg6KABhMMyysPiQ7ncudiotJRfwwNKKwYjZYkSu27qDkbL0WECj4+dXFBYb
IBGlDhigy/2ukVCr0nku9kfCUphFkPow4cKK7UjqDEr8pVtB7UPgJIZA7buWrzqr
l8uTkNw89jRRy2hnIKArWVh0UyvOVLs0Xy+aXyx+6ilppqR/omZyG+g/3heyfgrJ
jQcKsPUEjQPXUE/pikonwr6Q3HcSoRoP1AAmH/O+VwDxxFZHH6m+m+QP8MqGkTbd
aWe32aR1msUT3f5V/HjIkRovEEUL7iJxwr053I91qL3jfhAjJSAvqo9p+n0NcBsF
6CDzFq4W2mpLr6trijoCxu/Cmf8Ip0MpFDYOGxD3ZyvdJ5HzzyCj7JTy3LX7TaVv
uNCNLD2N35dpVmLuoc8TCjUS0Zgu7icChdU/wE6J4rhO7PTq8ZDspe6C8eRYhs7M
8eD7jGP9c+xtNVrEzrRPNYnSqGpjrdW9va3KtPHldUZpZuOt7n88bBz83ukqzVtT
LQTypU0Jnt70Y0MFehiBZzkKbnq4aJfarVDH+yj0RZ2J6LCJAFqZrKAppYPwLazv
vm1kTOJPFj0Rsjthywnsegpf2CtSExfNRxhfSC1vmQDyj8nQJ1s/RnnUrUHOuBEu
hoIXsFMvPihXKwn9MTNOeDf0qrb8Fc40M/DM49FCOwmHpKkX+K7izgWQCFXkF20r
pJhzfox8J0jDUAFtMkprqYp8UPdD1fLcRe87S7zd8qmYyYlGtBTSAd/jPrOeedS0
1O+t05gf8tmum8yAhz1co+JU5fVlFUhDc/hAD2ejvKISlNov5t4yNPyL4PgR9xFV
6r3Koo6mUNIRl73li0YLVN2LyQXGdZit4Eh3O8+yJeJxPD8olXQ9QRwhbUOJLoJA
Ctd2amCNwXO364UilueVTZcA4OVFoAESExFm6N2WzT+Z7u/sNYWmhHrawHRt6lHF
0SjmN4iR8zzURF2tGgdIrGp4y9x3n8Uh9EQI+yENv28qelaXrjb255RNP+r/7rrf
dioylh4vwKvKV3DCIwtbbc1XqtpMNEm+PybI75vkgh/kaSaXzZoDk4VyhXSXAiaz
uT8ZaIpqTrK8BN8YSxzU2/1bvIPA1XKKB4yhYec9FYU9qHDOjkOBsSouEbyITaGl
zd4KcGPz6EPylh0aO8KzwXilz4Dh/zswtLZs6qgoTczTxa5+RG8wwjmOvzH8/Mxk
MbjWObcoMs+siQAvQfYkvbWLiPyjDTc9RMssrR36GL3yvRjfBoyYBZMLMLceSe5d
1iTGbjQLjurKIGxW2sGx3w3gaRfIKyfYQ2w4BA4xs+x+muwmTh9uTiXAoZERCpjZ
9Z3YcKwFQTfYRrWFXwVoCUZdS4Q17sQxoDtD2O88ds0R4xXIcmonY/ILITXPrYUV
TIPzUihLBYCE53ukWgWDJSLrUSY2zCjuLL/Y+k5KJMVGbrn4hyxzFFJjYMaZnJEf
LvZW+KDlE0MqFYPUYtKygpTmhpRvDnwfcscEp2B1yIatOAro3LhES7q/UdQ5yJCN
wz8idCGX1Zv9kotZw5ZxKT1bMzACpuOqse/AUzZNfE3wBCtSjbvvEM70z8Ua8GvX
RGxpjnDsOEJLOZu57hKUHVqvgpER9M13h9oKvr1OY1oB3EgxvJQeF21MhQNuPXeK
9uVCjPkcoJzfuWzJY51lOa4FPtb0j4bL3EksL7SMd9xX6KsIOaOzEZp0v1XMEfLI
SgOEU3yMWAYRtMtmk9rgbhuzXjsAfv0kTC79J4hSDHuAZuAAnyJN0YEZukq+EBO8
YvkNno5YaFBHARy70wMXv7JEqiiKa89//KpJx4ZoqFiIKaEQ1glBgAbtel9C0/MV
J/C3GOdfF16yChmzi27yN358W7gLdcMcON5cXow/n0FUSSZEp4b9oczmDqTFeFRy
lJJSnvlP7nkPgEdpCY5P8DmWZePO+coV/SZUXY1mACrPOEHqRLe9DUzMcAVNDXQQ
SG/90+KOV8VOYJihl7jN3Mb46aIqgnDpe5V8nSo68X0LjGeFp17r9q4qDJRdW6xi
uGwunPjQMEp18Nsd+ip8O5VcHlrvCM6dlwKucsruR4azYTwGXrEHwExTFW1esZv6
AI7PQK5OgNWT1QiBvGwUGIfHY+ZMnrlx7s2Gee+S90DFFVdKzAFOSKioAoZPK7HA
pLiVuWy3M2C8nAJRUZZ3T97ZWdq/7R6O/y158boGgXvzWv12GnUkGFK4ktvy+1a7
lOvZqCBVp/MLebsUXsW2KMvxNBrfseCAzTA8dqxOKlMKj77qpMIv/fkJr2q25+et
SMDnFrXbsOfhUik0BBAkmtF9qt0Shmp8Ou7+KkkdLaDXPX/Wnw+4qosC23KFe3Or
fwdVTEFC0i3im9PANFSP5/P8M7YtaLK8oBNCDNVjvcuiatnCFSYV11StW5Gciobp
iRF3ZGAPtku2Vvz2woOFloQ9I6hFDDVM9DmbKdYI1+Z1kU2Psfk9RRn7NBn4MGhJ
bNhfaRDWeNcouXxB226Nu/3JwPu2gm0XZogA8MWbNSQpsBqneRTgomhD9E/6nzuP
Szhkmgwo/YL3qIAjFjRINjXtDPdM66ipi0Zgx9l5PK3/cO+76/sipiT9MPEbSI0j
9lyJr3Cv9pRLQCpUwqOuEXH9afzZaoUujOCqZm/I9k9T+EcTk5pdMusgZETChEnf
lR7wtOs102fHuq3+SbjjwO8nr0yv63chcGw5r/1wbKTCss8sZvsynCBu+I77RO9z
hOzFwu97AgfFcDyeOqf1t7Jdq0zKG6ClEOhhpddCRwfnbmzFAI1rGk4U3k1/Sfe+
lb1lgpQil5lGkS66D9iUH4umx27u88nvtgG/m6RTKmD3sMqfIEi9NyiH6mxU2K8G
Uk/zYRbdaJAdKaYv3yWrM+kPlJXIOTuIv+kbso56V5+Pae27UV+Qd07w+Yn2XLb4
67bRuRd4P1Q18Zm9adSdSSCH9Upq3pED8ZjA5KMug6zlX0hISzygCyoit7ZL4R67
03ufSQt6hOyjSUCVhKK5gUlsmG3PXuTt+OKPDPMaHN5JLtEEEpzeMsNiA7kJoXc2
vGKNFvKeH8ff0fOL+aVfZ5DjBgVQYrDPR8RZyUn0RarzXr4WPXFL0syAV0Vu8PKw
zgRU8f3JRaAy+Rh2DSClN5JtxKmtLJx6W/Rs0RxIU9dovHBe+RFK91kU9YeWsHWp
7epFtH8RaLPyxFgSC5FPtO6oqk8XfBkG5uBEra6AW0nAxhSrAyKnJWUa5gflS6HF
h+PqzSIL7UgnMnFITDkwQBZziAZTGZA9+Tu8qhEs/2iPVChvP0Laug/HxPzKRpP+
toJfvWVUT6O0q5fY98jSyoy/x9mGZtXsIdsh0BOGLEp/La7pEKCcB3C5b8mLCxXC
hCop1CNQ4+GsOgHE7QeptfA2jJK5fgD+cFzwkAf4x81leFbI0gfzqg1fSXXCnvsq
l6eoWWuEOlyTrsii15RwcApSl0O4vsArixmIWZOkWJofDw6B6/POfKdjm6NfqUlc
epekSqv4Auu7Y2zhe3xgmFiFMacuTzr/wpsCXPYnFo28vjGDxQ4uUYfrmoRwqLEt
fLIvxLpGuy365w2Ly9FYFWLrF4IJDRwiXcMhU0Fy41TtlZmQkAeKl3H4xQLUIzdw
h59ljyUShWDA1sskLmpmehvhCuw1edP3CxXb/xpxjLoIzkWxIuT8qjKpJTFkN+Yj
xgef3D5ejHosFcHImOjgVIQtnd5//wwGsDK3D4PLkKFHLoEEVMcrfb+Re2NgDsK/
YyfCypUW9Vp1cLCfd9a1PAFXQWI2wns7WsSfEHEuby4XOd/dQjOTnwIYN3lPuvBM
H7FuC4zNn/EPKbFvPKUw6ltAaSh2OfEODkvgIwi1YB2Iw2HgRo5WA8WVBWZJTuph
92YYiXkmPa/tCJCtfr8s7LF8ahjIYcmIDuuK+FiX7JiYnScG5WYLwFeK1dxihMtd
AYquFiJhTwKCSz67BGnK6lwON041Ab1rjBChejFaxfCT8nV+APVDl5YiQY/MmFnb
GklO5qv4wDgNl+0kIKnJtVLQlp0TSWX/R/KRkpo7mrFPFbr3g0ZesLELW9lyiAzo
N5goSDmr4DcMmxJrTkQVt1HpEMmZmlA8G23hmHS8iSBZiMq9fMUudKz+NN53NwLU
Kxh7mBQuDTxIljM7PaoBOyVBfwMjW/6qDLgOOkE4RIt99r+g+e+nFxevLZI4nod3
E79iAAhyZ+3cI/cYqaEy6RyyTO8HxJAj0aL/tv0XP7DE+pc4azmV0XhWIEFZXDcA
4UUT2kDe5zDH578o97o9xZLjGKh45qSWMcDTjy0Hu1AImHKscgfMjzaa0GZSoDrs
Fd6BeH9pbHrsfTVjWREAcdBH0Q6mVEAGyeiEvXyRri0iEOcDjg4xzVzQGBqf13lm
cMoivPm2DJQUu3Wri6ZTgudQ9JRyL2MKSGl6jgxDmQrRl+rAF7eeMilFnfx9MT1h
QXv6t15yy2x/BLafb3pMVyZk2dJ9c7cF77y1RsJWgGnnvLfLbHZxMoJYIkyWhFIY
oCEbhfskWQ/Kg9fJt09HA+n8qlnLUuWg09UN1vRxAdiHtRCRPVu7mqh0aHkF/Bla
E6sSBx8ycgdsrdUpumyMVGer7ETz6NEOWcrOeojDQZ4EDvryD8gncE7qPFuBUiYE
SyJszkn4E2cGaIHmcZVxgW1LFtKTK8BwqfyuOc6RGOEGsw2M4fbeENQpqoNv/RT7
3D/e8rTVisdOasHoMkFPQb8PcHPPi9PW8lZ1u7K9TqxZdINHZc9JXv9wA7As8ZvS
Z2iToWPqSBcgYgn1dBpLCFWDXypQuswiL3wQvSr4ORSPRcU2/fp1zbE681ElB5Qe
jSyuGthFs5BesfzwVtiXvbzlDm8vNMCsmBaFUrx1l2y/lI2tMtKSM1PaDToIxljB
hPnzJ0FBajb4N/xpw2nMd8Mjq3QejR44LisvxId+hKsHTmLSM+k1cWYCRg/nPi2r
0cIo+XRW+akpoafRbJK9i10s9ek03CWkj0gH9pZ148Q+CraALHRjyPUISFtZoiIo
F3UyzCq9y32CfSXx9dpUYoODz+7e+RpkUl7+ax5cGeCvyf+tH4WWW0HWPgG+nomz
o7waIA6JQG9GTKoLtJwA17/F9wIh6srwP0yHExcGxGObV9jeEAc09ppz0HsWo0lB
1wzQWbt7qDvgj53ka2LmIf/r8XomW3VJHbO9eSElRjDqSbKvKpvia4/rsRfsXLYv
ouBbEvOi/KHVYzEPf/NUS0nH7YoVtx6194XqIkL9v7bWlRBAN69ziTmHUMh5h+M+
5hBLRk+cwDPwCq2B5IH0qgZIMnQYDzX8+yJPKA1yN49DGn7FJIIIn2CTfAZqxABP
hFCYXLacfcBcRbgB2BEt0dNsXAc8CtQq0shP+0AfcRSSsdlWYsyUHy64FyGQ3ikV
X/AQPSx/1U03mI32E/y/RhQlnd234tze7Q9OFzgyGoMiP+ucuk/lY+K4C/FXMtm5
U8sGkDGMXJAjRhLt6GUHjq3xLbtIIP+zdNyl3OyadKpo2ke0TB6rh1mQHtenxTiE
RSNu9uukYDap5HfMax9VGM0EltOKGgXnv5CNnnYSjkxdv2VkD79dL5x3QFzXlB5d
kzpuYIC9e8+OV4LSbYO/JoxFp7d2CVZCRsNLYmg2AollulRkT6IUUkWtYPfQvRhX
N3jQ+w44tfrgYn5Ovg0Uq6+9fo7AJbKrHPfj2i4bYhKaa/63dkKywt3rRRYI4dF8
fIhJ+2DrBbinghHXME4G4yFeLZs1fWaEB1By0aEoyScoF9GemL8o9HxcriinjHAP
Cono/E16sKm1HCtHBrOdp4XwGFMmE+gPT5DeHbagiOPVdmoUMxz2FOH8+XWJ7z9X
8xUPT7nxHTGFmns67KueuQrQFEYaXqS1gtBA0dAhTwqvVq+LuQimj2ZA4MD6jwTM
ZKg5osrzWiA+S+VQuvWUYzoLJl4B22p5WmIx1x7aBsC22atyWF0YPwJII8f7vNkb
YdbX4II2WLtvSl6vOHy/t8c7BOQIHhGOMJqRBNLONLCX557cBVR2m09ZmajPzu39
9QjUCPmX8UNR71V1pNEOIJ6p0ZAEi2lpGCItd6NEFxJWkdpvqBwWwKDLRF5nj8Cx
bA3XUC96IgzYDej9/Vp1sK71cHQ5hJcpA4KJYhWlOcGo5xoQRFEC8uXkOka3sWas
Y8jB0MawPatNh6X+1Iit0b5JwkFeGdHaTapzwYBI4469ThD1tAsOcH4Rv8wF0shp
hfMEoSHkEtWsPCl214ZuyOmqUgrvJiD28eKRSD1+E9R7ULZsY58fjfxx3DtbZ7dD
ybhSmPQhvnL9PYg5mTlOTaS8+RUNM9gRhJ4K85bKjr7DpOPbS0+5ceTFFhNMX4Rt
HWkjqkv9Yq/JWBP4vVx+L06Kl9A6WVRVutnj49AVijijgETYMHWm/+ida8vEGoZP
Y8L469vog5nf4pxY3bVhJQcdED0rnmGz/vWxOhiWm+HIP6ir2zikSJqO2iq1ZsED
E28bN1t7BxUkT0cUfWca6k2Vk7ZdtiFLmY6eFJtsIdzDOY5uhfSOwdyaJiGOoYii
WQKe81uXCLRK1tjbGs4v6d5RkQlVsU4KvbETGX6XoGshbUYdeM+A5YzZnM2TwY1E
VPetPMCATO+/q9eNof/BKJqyAIxoOgVXNSSYa0I09xGxL4dXmSeguafXc40ieiZa
OH7GAL8rnw2GDwLJB10A8bgtsfzUwwzpxo6YypqH9AMaCRdxYGDhhJkB7lcWAPcY
Upxl08EucTQph19htUGqTY3xqImO/V1BNApMoN6/IgL/3mer6q6SCnMQLvH95cfJ
0+KLaq0ODqa33hIqSiCtyqm1DyEf3Fg1eXqTVFYZ6bwRR3qndH/uAyYZ227JKi7B
aL4NhyeJXAXMp+fGJpqn09qOAQzbTdAGqEWyiTC+KPDMsHM8LhuYAqQHfr0QZ0nB
lU07N8dEgSEsF61Ne8MvnxAEoz3GtF/4iCIGNMTbA7o3GzpWYbZKBvvi3n59gJHu
Kuy7IX3yR2+aSWGO006M7DxWu1Gj2QlA8bHEe9Mx4I0IC1ITgsdWp4WVpJ+iBs3w
wm0iPhHASrvVSnRBVn7Mo9syGNmFXg/TbVvQ2beXX0e4Nv2noj1pk+EqrNrdUjlC
Beo8paKxMz8gbmolgkWonhbJxxc3pWrBw9UdvPuY40m11haBFyX0F8FUdyFC0Gk3
xBpGKiNqmfIkQEPICLSWhmdaaPVwcfU7VS34XtwH/qTvqBkLCqygUCZnlL4MR+pm
9Nn0s6CvUOtTNtxrwofTth8UbMqyPYf2U3SzmChnqZ3kvGXqbQZrsyHxnG1oBHEq
Lnropi0wUGAeEP4/0m1/f1WPUBo36NVS5GxgiTVzMBpfG59rcuLhC6TLiEykHfeN
TrG7ASenWVCKW4tQ8jLC6R5iz+J1g8GNRiENwNXxEN269ABl8GyOfMCXkvJ5JNyV
zywK+LBsfESQ51ida75ha7U5PqZruUJGEgJJN1Lxm8Uh7078MhkLyAcCuvwovuSn
57ukNmvulsagdRLOyqWOCl4PLTkESEVUZYz6y0bqzZaLq3BGbj9P+Ey5oNWE8crl
nXCdPlBwaE8oVzLJV8gABo2Hpnnw/fherVcwliA/s3rwNurXIjNQ89swsKZtJXnj
JQj5KxjyA6fZ/okhWUas/+FtXIfyGWBU8j/cxJt3vR+qhG+2+xd+9ZMF7lcVdzuZ
sJhmxKVHYIHvJq6O5Ui/0+C1WvCKyFQrRSxcwREInJkAcfsDU1jhCg2iIk18Smc1
GgM4TdPAZcgeNRJOEcmR0HNe7jZF8E+o2kbC28xUX/cGj04DB4WijD7nrk/bqy2I
kF+WITuWe475JvubShVsoz++1BVx7Fa0uKv3fCGsvqDHL5YAKwnfol5QRPQwoUxk
fg+8kNhlaLD+br+ry3urREffknmSc3SY1ivL5qNBUANJwbZ8nOqemVTUfSX/r/XU
sO92gMic+C3MwszLQWPcVrTwPuIUo058Ywk/EMW/8hoWPk/D7dg+EzkERTacpikb
0eX726VHsc68exC3qG+OHei3rjKdS/IWbl+u6p9hj8bSoMiIBjHhOvI64wvdGcte
/IgQzkXo3pJf5QIQQQnWszoLEVzTBCgf9cWJ4dNo0E+eFZPP/nYXZUKb/sCE3xea
NDS9v/f6YZLEJssDQoWuRCuF1iiebAPe2w2SSJbIk0YgPbx4wowk4ZBr8AKD9GQx
YItVFTbXZ5yo610H9mTUXNE4RRmD2sMTx1QK8EQwMBxsp8+J9eh8OWXbBz1oFaUu
XfJrR8pAGWxbKzR9x8rRASQ5w9vShYmpDq0Dq6rJpe2rWdNM2o2wZgICLnf5AwH5
bvOMJUo+yPBoBrf09aItnp2lwah/09rSw9FoOiPJkcMgwsXNrKpRtPI6qC1QKdri
lvs4AvmdEUROdQi5qto3QgmOXDN2MgBaJPalYiyzfkmOxjTzyjttfEwK+H+iPOeh
eWWyeBRCC6523+5fQ39nXc53mElIn0LyuQ9QWc789EWsYNhVPYtMK/ubtwhB1I/X
Kei1Eu6u+PL9HZG9SgK/4EdXxmHM7a8OJM5EtfdsQjHD1qkKa2GuAxtmRAFZSX3g
inmB/UhDLev/JfhlkoXf/TezGGnZHX0X4u/5jqLWMrIlDpgYDCWtppdRSZfWExlk
zQBe/e7i4psgSnNNJ5klvtjmPZPn6x9dgbDuaEYBn+PStU5m04UsIFIPrCvR2tiW
wEa4KgHGMLgZDhiO7oM0kAt+MIpNQQN624lazav0PfP0G5Hrmx1KUbBSqkiaeM39
kgqfdz/yYzDfkTpXz215UyGLAJ8vrl37lCBAOoyn+361h9mAHRq9JloJBAGucrOr
ZV9tq2dzsscyH9RZGY/foyn8aBXGg995VGO5q/ZluTt+al3rN7RBrx8oRaV2T8/Z
O7YVQ+KaZ9leUCA7IXpatKTMx+h6XQE2REMWgiZLC4gdJTQLBOiJbMwmCrp3+1lt
SEDb+JTIAVFXJ+dbYdh+0ZpcXEYSPyEkaVVPj5HkIgltbMtWXcnB2esSjbqUi9f0
ZFlb00QXv2aB4+vlH861g+SKDPUUCKol106E1IdWJyHA+ZbUdomfV1n4LFcglV+w
QT0a50KDjn/nmoWC/ooTnplc9QMkFbPeAp1Y4+MSTigdO9K/brUEuL1ODRhdmAKz
LfRND5XUW+qhZfeQ9w9AqcCfCSuHxpCBTKQ8SObe/Z1+FMhSlAWwFNXvV6keoCR3
AIDbXKZAUdJQIQck0OgAR0LVYqMBQeZwjolOxDhn+N2oyfPzPtRnq+vvbElssB1f
LA4lX6aLY5Vy5u/E91cNQfhHBJWo64+e7fPfNXELp9UPo8e3juxiZZgdJTrnM8wn
81xjTUq156wnDcp6VY97c3wznz9Aa4st7YmS2lkz5mwlRlam7zr4QuuCvLpANBZt
hDGKv3uIHHxBWJpgpW+oTL92JeHYBSGQuv0O5Oke269QeSbWYAWFljxdOPX2Qi8/
1N6v7t2fQE5ECrSgMG7FIGGZ+jx6tWwKQIv8ofKuZPH/+QakDNICZGru+3jAJ3Hd
+N2tm0BRBGwWPxfDJzEnLWzULBBnSbBIgPjf5duVs0SHmUGGcQIyHYb0WMDOZPw8
zB8YeBRCRhw5aY8Nz/7FuHaaHyrXg1vYMITepveXhgF62ePbpy7pvpDyKoje7ENm
FNTG+d3QVnM1hmSCi+aXAn/e+XW9QHh5dnc3BIzityzjsjdyG6UE082RlN/JrpCi
P4mEUu4yNvggyf40yX3GtLDiMS5rEiGzKiab/RpcuWxcj1rN59CcVGyhm5sxR8NK
W/81vyANZK+HLqIPP7vgomkblcuMu/H/3+tFD/BSjNuHNl2H637YLy5sI4nCicDH
kq+iB6dCqOknGmNTKNLDmzNHCEUWpqq1uaZXHVCBI5gBdXuEesAHIf10jZeFuS+I
4p8dvxZyEB3Tno/DiB6ZWvy5JgLO11i7JwUnYyG0qIXc+N3ju1abAOzxzD72f1rY
zwgrcQom1o9HhDimCNsVyScEu3Y+Cmyx5Q6DbPD8btloldiwYYR16wM0zcOWSy2v
K/qIzKUyf4uuv7afNqt9iT4/rS4bnFeZuXOdTF/bxCpHCXipSj/o9kK70gCO8JF6
j//QHdkfCJgyxdrUWehplTzwsIGteBcrS6c1XWkU6aT+TJbUWBf6GNuumvBjYJ8E
KIeeNQh3B+2ukFGfT7wluTzpDSPOqSou+fJNrPNBS2GiENxTek9mdZF4Z/xvLmkq
iywClEE0EyCMYcJEnyCGME1xZpivLcvvYBN6MJQuT5U0Cb+i9ipWx26eY+LqSDiJ
D9/mb1llgvze0oDP1crjH6vTIvxtNFBZjOLy0hPGf9H8xZlgL5VOaVsO9Sk+avWo
g//WqXMg53KBlHbllR6aYPaqyYcBO39XAMMVd3MzCXcX1lEwJFBw2La1EfXbXYMp
c3JIYyJEgBdPSTo5wKeeBQBGV92DxZBJ39ZewG6zeQWlmWXulJPobUQXoWwghX+V
DsdTDn+MfKdCHY0c43dcFcvOJST15jtIT073iMEiFpHhUW0wnIzvtV3XaqOgdPn+
RgEAFeYD9K4OkK94i/ivY+Ka5dR060sN6ubQ3xAk1rqpc0LcLnRdEJvlWhtr8cEk
d4Q/YWSTvGsxMHEWslVQwNPxx2q9Tl5ms1cgkCbWhEOftBk/GuaDUYmxg3yHP2NO
cjWpghaO7sM//4u4dKyKE0MXAwq3W1ADZwCiX8SvcVae++2W2vIsMVmwvOxAGC5r
duJVwCclaTNwniXikKnDfxZdmnQ2pHaH0AnXe7MiiiQxC6tLTiyQyZLiduGlFqDW
iwgRn/BSE/yZj7/sMWrTRYNY2K85AHlvoldfTXBN8Lc5LdqrFRCh2pj6MQud0aSR
yjsjB9VNQuxb5qM6gaaaZYqCOS1SJ9Wcj1BqeuhG5R/cz2b/dmUkfA+46mQZC2o/
Y5kkH98h8jLl8rMYhpiQMX5YvOoo4SYPz/3r8VeMiNvRu17iHXga1lvqMnPbeOV9
55sLYmn5cWNhx5MqXE0iUATv29vKeP5MU44Q4YNtNI+qYHrNh/C6LQi4+RfFZh36
1GPgFcnoadXPLNT3CiBi59obmzEjMgvX4L8YUjCdJ+K9ZszOFhTTIMM2TmOadvq9
beuSwEes+6PWjGzmzbfokw5r+9VnRyJ0Rwm1Rm7luenvh51he3GNHqotcVUwCqWA
WcYsmmekESJSvpZUOvb4BuNLMWIFVExnDyLbqUepuTV+fGx+F3ubol7Wz3bKrnQj
Lh9LURKNPoMcCesFDrRl2iw4diKDRqbKTgY6G/vk4TYkZytZENOUNwtyqkehb/tX
bAc1+HeW9m6fV3ywidPx86cvNEVSSrHwJkXoAsmJPu8gRjhtcWZl/sT4tjbUv9fa
VAUneBdsv8miYtWySwM4BA4i4J5EkM31O4ULKehf9a1mZGXdEwY5iZTiOaMXFiL7
NZK5u1g2duE2EoXqvfxd4egQdM5M2V4nUiM5fDKboHX8Qtf5CNjlDDpu9en64OQC
T8sDDh8tA4DII0LpOP+OFtD2VORjk30KiSrDJ/RF1FXwg8l7GBJMhQ+ca4mn6vUh
dIdxDOOBYpUJdTAxjYeuWbO9UnORNbdmKo2fUt98ozK5aUPo+EoBzn7QIGeykF0U
hZhZu8MqKNve7k+qyxepTfcDn5R8X+n8hvKZgsTwyvkqh1y1Qrb8cP5tsE4aoReT
wWqZFqauxPigDNLs0ofIcVSCXSoKkxoiaBq3vKD8SmyoChnDLeS3AEtGxooY799N
MQrGg+Esvz7t4/QAQNvZDjzdg3TODvxYDlF7SHFa0g+Vt9GbDdJxxu15UCmim7v3
/WpROFABW5ZN9XCBA+uGKeY3t/z417jn/6/38+B6JMg2PsHbRO4pugh5RpvZ9fSZ
Y5/60RZ2Bh+1Jky6DGHedVG5O7xEf5a7JZBtSNeMzBwm898UF93+DSRnX6fbSsK/
oIJSEchslPeiz+Gprm32+q+rB9kVVoWx+Qxi7999+OR6BDgipKyt08vjSS9jrcbC
mVbLL843EO2vIFM3K5Wv76FVufDv1hsogiXxBqlYSNaf6Ck0RBz5VWb5sC+i8TQb
zSDOehwysDsp9n/ygwhbhcUpBopv9aFKehlKdAPezfVcdk6ByXwRv6k5nhCJA4G8
K2Lg1y2Lk11WpB8R8Mn1HYWOMeZpD/s3mvZRk5lW3vcQvj5BxIQY8NLabTxuPQpa
3AQOSplVWS06IONNvk1Na1y3YT1N3h6e4b6qecIw8mTf41SN3vmO/tueO72o5ZI/
KuVlMNDRBxpI2//JwVy48AZViNwJuKWAi7Nzo7g52IGhfC0XTCfOlakoSJTn/8ZV
zT0SzcsY2E+jcbilZ0NWxHVnif+IMUwjVTSfRWI1YunO3FMXmlc/mxcEvJJGSP42
uK0zFXQLXbSAB0Y3yabG2ReseMBWYvgwP+zF+jIgkMPn7jduJ9U1iIPMoXymFaBM
MVwBK+89fadXA2RqW9h3lMIVoq1/8V8XanwAe5hyE9e2viOKOmw7AzC/fazUt2ZQ
/AeUZMqnqATJQLz8jMbviiPEj8pbFyFHUIHlAEt15KAMhJtxEkoxC/W7xqGJRlBI
z7coiKAKYuiCwBl7WL9GdWsr/KozAzw3ycXQl5lrmFaYbYhnsByIElJnnZ/B9Erh
xKFEw10N1pZKj1ee0sn89RLcJ5QwYG9TH3pX6VqyJNAb4GrCVETVaBzjUFksyLLY
wM+RdwveoShQoTByjDXjhfHdEAkxaqXm32RRtcPFAN5OzguTeGf0ma5oxQqvHltb
4I3VK+ATfeLRnIUrtd+O9/598kMQSX5ppmx7q6ZWMLbXRm2SNW5XIPoHyBe0UVYQ
rdwoM9cxToNQ8Hdb1F6shAeoAvNTjoxjL2BcBZBSE5+NkGtcBkD/xZ/69wFurECB
LZy8l4rjJdKcCA+8NrSljkoiiolD/qBLGjTdjH7HEcpi9Z4T7i0lTUW3/29akgYw
Y0iU3t/ee5o7K+O+FtwbeHz8oFpNp3Boyi3aWUDfjtpKVfeYRUw3Qg0RO0syV57j
Ah9NMr7DhO5+mTsgFMC+Wl1HvBUyXnshOsGyUvWP5w6doRlt79O+NKFdkDsEs7B2
leE+hItGbNC3wDRF2TPaCQE9H/v/TPGp373joy2/Sz4HoD6bdZU0ALsrUAw4mJSd
N2twQUrYWZGXAkkOuc1MzOljJwyqwNstDiTdvpWYl54aPHiUvaludb3bFxLYiyFU
THkkjdVKzKoBMDTfldSSE2ER4EMoCVBofIXJVhdabG7hmH/pmY5QYvcYLfwS+rAP
yjSCNh+8BZv0laSIiQynhQBTUN0RbtHLtMqW75noA7TMtOCk2w4WjkFfUSRereO8
lVc7fzHdRXva+5Efv5oMNon4myKbsqWCtz66FYLvrt+0EK9qiP9bpMgVrileApyY
yhf1zbR2y4Vf6gugIAiF+jpgIzCiYRnThW0J5OjpkQrz5S0KuRwPP7H3xaMUc2rd
LHt277P0dqKDmabPspAQVnnm/xo6AL5N6a89Qk7ux5vsXmZ7ZVgnVS/+eDzeB8ya
cCOPAE9ho8I4ObfDQ65CXX27rnfjdOY0PjhsjCnWUE2yCikBFfWRdsG+DAUliBel
dJ50Vh3gey4nng4ESkgia+o08LG8yQgsoPYi8SzXhaeRl6mQEJ6O6EuH2EN55dgh
ZIxm0bQmsge3CNqL3eWbmlzkjDEruU4Jn+q5tOVr//xqpbormR2pinuAwxMX17j+
ekcoKVpIM3vfCWAcWkkgKJscSyApvSVm3YB52pRDoBrDgBRtfyFuFGfS31+gBuKn
5JSoWINLV/7Oxf7FsNc89Wxp8EFLODBVkEzsndxXeifVAkl67sODEGj0u7IInDjV
rZdjSbHaTd8F2nxl1um7y7GSrK0sZLbYmDS/F/vC7grR0lNf2EdooMw19lgg5DJd
oy6qZAw8cyarsuaTqoGR2zZCk47HN4AcmZHmGGBd6QfknukrVc1+WFJT7Zb9mqDp
wSFULvejX/AjWf/2JQKU8jm91yve/PB1iZzQ8tXxERcUZZ3BnOIt8g2xS/M06bfM
qtSur1Nkt0eNZ+i+pRuQVlW8Mx+hI5WfRMgoXZYXSJ+/RCnck0iGXKJQsEh6e7ea
MGaQTTnI55PmWqPEAAGYCXzRHSqhbTjVhgFRpWzvoWJH0dZNZdIwn9uTK3g9P60Z
+vXPriTgYNYuJSkFD7kntgA3N5KEFoPIp3F8yGJtX030lKFoJlImqnjSjJuXnnw+
dHUG0FaGgGJGg46rl2QWZ1+ygVDsVealj9aRWX65qkPFkrUWjzjJtL+WajhARhIr
o+aMN8FQApAAr5w8psBHlQQPK+yOE49gj7PFtATOzFyeoCwW9P/cY6AoYPJTgWH9
4ZzR3+gi+P5YBxHhDD1RWZf4PV3wqKI6AbD/2FhzAXp5nCe/nhJc9Q4aAkzrZNPE
39wvwl2FomDxHMze4GowmKOhkyptjnFRKL8Q2MMnb7rOd+Fapokyxv6tm90bX/Wu
Ohe9JvwO7BiSdqG4KQzOgP2+3VzJtoXUi7MnCC92CxiH2JBNsZp/v5eS8kGlrcWi
mgW7lSu9M3WqdXvGNT3acfqmEPO2VkYuozXl5YM4KxVSR/ff5mMQr4aTqBAoigcL
s14XfzLk8clgmgi4ygwsMm09TxO/BuY8dId4oEMlbci4ss28VyOHHV7nhNuEEcYr
eqw+uHALgtqBrtb62Rd8DCjJy1PHTRnq4dU2xVgBDX21EuO5Y8asxSIHK4Xtw+DX
Go258SSQ1NyqUuejYuxMzPIkw7rmhA0nSPdOn5E+yTebYk1tdD9aHou61+DCGyak
N330I6ebbNm4tWk77YIv0wznBHA0fMTDyCP6VE2fMtq1XHTDKUgIQQqb+SUogYj3
CzZGUHBIbn3/ZPtovLAVqaqv+lfThSxSQCuULZszNTQks1MGBxEgOR/EH1jYq0YB
Ve5+AuPW/yHulrLatYPwqWIKi35G8J+6SIJxgHgRjoKQ/q70jBxAZEj1eSpYnnhQ
mgOgK+yV2lC//KAwFbjyIf4FLSTueI4nY8OIHpzxboWx2d1bE2r60s8huLAp84DC
nsoRUF+A19WNhzd3pjxpaayuBgTm8aCewQ1GEf33Ymwe3G2x4I0DMLdDiyhyJP+/
9u4roejrm2ydz2JZlcqtbc9NNaEOrweA14BtepKI6i/HG7YjxrVNsdQtwdlR3ocz
pTME3lFexk73bxPB/abNwz17HFxAvljvVEKXWiGnZ4umXDSNT/qA8b1zQ0yjODLm
afz1QA7eo6P9YdzWvktrJQsvVEbyUFHzkVNXoMdo61jwTaEAQXCBuH9CfgTa3AMj
Ngl9IjQYFUHHLu1hjbs610m1462fNvTaspY6mf9fVUNzcEJSlcINuSMmygSgiLo+
sRxWY4ieVTez1ARvbwOdOWB46+SUF3CASfhvjQsDau5TYwsa/aAwZV4OrAbkhiKq
QjaFxAWI4+C2Z+CQrlG2Ucw2BdHtUI+AAOyq0mvB7L8C5mFj/IHcNHiCWi1gHSBA
jpzU+XO3yopKeOih9p99DvQUaivBWxD3fpsZugM/wNxhAQjWF26+tK0d601yTKbm
naVVJieVHBkvuRvMljSQ9lRZAfBcJtq7o01PkeH0CHXtppX7EeDdRaa52T3sOK5g
j+WAj8mhdh85hHy6MrNZIqOVWfQfp5V1tVMYvtLcxunO77m3a9IzCtLSzubN6cIt
Ls4jnQlgoikBIRx0OVVOzpIoPY6qxerVITNepxy4sntRCC16FdOvsM/XDmVvtNdj
n0QhjFqa3edhq8h2MwdlUkn8LN/rk7PeEFCX7H7uaDGiWYrhuYLfibjmgnbUmkRi
6Lvy2hFBG1L8eD87bK+KP+XWe9zyhhRZ3sxFGxm6C7rITBqEeYGHITgd6lwjAYQI
NVN54a54dx+Dsj2koMTHAI3jNLtRim0moYy8K1ebtFLvHa2UkDiOzZCXQs+wThYv
JPnfdVe3SmxJ+zPCs3pHNXp47YuPoniUoLO50nwK6SYsk+2W1K9wtloPSgpviuaF
H2yTcHAa6pXLR2JJ+iWSdKhHaC37xqfMxTVYmqHyYal5b6XprKP2vINJZ6LUQ3VQ
DPfqvabECIJotW65xoiMdQie3T+nL/UnDkRrwUESDKzOQQo2LDa8DhNaORdf0Lbt
/TK5fq4AoWOqPN7e2XtQuYhvQdGZbGp4dmz5tsR6HmKyJWYRZCf88gNWWb361SBa
aam1LjEVJA+Fc3wVrhjBSfQz7R0PPGp1IzUgEO1I123jUG4WnHhJmy9W7ntRq+UF
mYdlHTYjT91dNEvKMj51jRUPregjLjp5OKixGda+bQ4+SPZ9KixakEKh6/gTeM2R
hhaXWmsdCYQqdWEdmsL2dFJCqewQgFLI89Ni6v/XlZYhZgGQsbi84TwwMtajSx25
90ZYvFdGcOXm89P/+AEO43ttvJ4HjjvdF+XrRXoWoVo/3UAu/a1X4Abqf/ThD4Pi
eZX0jxG4UHMteAQYaOhF/aupjOyXecC8NfNYr1Erb8vzy7UnrhvQbSrC6dNHRcEY
A2qFYOC8ESlNOf9zIL6kEMkUKTy32VVTlW+bSt7R6dVdYsIISxQmxwz2HJxB1KFg
HnPDZWasxoqCQnuAItfvaL8pSmw71jifO6CTC3258Twp7ABoUEOxiaXnrxXKlBM8
IM77BJJBebEkkjcuVlxYacZSN/Xuw0igzoit9uiFtGu6QehFvH34UIPKG2qvPo5P
1GwGSKqDB/S1MXGYMkJP5C2VZIUxViN1TOEg7M2jcdvWYHg0GRU+kxU829g3tBG7
ecBJii0QopkgOpM58ORwNncT5puUJvoxDlfs6ThMwobSunNBsd8M7sU8d6vVPySO
o3sEXOp12chUhoR336iiVhA3mnNaasMRWr7piCr+dT9YHy39pFBonApoqLh/f0wM
F6im4+ZtNuaIt6iE71j9WsDOIzD+AMIgKyl+4cK3ay3gpJVStoedYmphTGQG1xBF
WiPW+f+Jh33x6B94AgW3knED2YEdfzRs1HH8O9JIXKCHqlEk8g/lfOI7QkQgSFGT
9TLaFGzPBtiw22GpEQcOGUDHBy4GIXcLX7gAmezh6hqgGelN5QYh6Y9H7eYIjk3X
VduwBEsxLSj91ReUes0zm3NVfJF3zSXBOjWeBtzilEWz1xuqlwecj02PwHt5y0G1
2vRZfTd6iXqxed5FlxB8D94Z8sp7PZL7TnmCFFF8muBWn/phIzSTfzQlnIEKROwa
VXIqV/5P7tWssfaosfCYWn5kFksB+T9oVOfeeScV/Y4ZippfHkK77w1EgqN9wNVf
An4oyIV3CWu6ocD9sOV1ZzXWJ2viJ/OxEzupLlEepzKF1Tfb0wsUKTFRJFOhTRhD
yEWZYmrK26kGylY+/JF/m+kseuUdAXf6KIsBMexJLuo8cTRy2InYdI62TYQZEF+V
AEBJ3xGwRW8PXWVWseEJMzzS4EVCDE9eK4uKnx7pwLsmAiE6AazGKbFDZDg6W+ww
rEWAXT4MlRYzTNLxHcNUq9+WMGQXUUFyRa87mA644Zh5eNArC3SrXgZ6whzy+1oq
Aw3i4LfeqX07IS6haxs1bujh8g6PmWeMlx8gYApy6RZwBuEkVEjfI30bixDZCQJn
wCopf+TrOY2kqVVTJX0LR8iwm2xxGrOc8s1fnnaipcDMo9Rk0W/FXAalI1WN//S0
o6Nprx58KwzVSJ9BM6s/uLKNvsjrQepgvoD1f3bKpcUjBSKpz5ThK6sVU7Ktt4kR
IEUJd3MJCTEaCFJQjlQnfchLhymbICncrZM0b5NQWXr9TXeRC0hY7cwlBU6SW247
KUqEx/buLflstCDEwvV5WJmDmVumQjzkm6FOCNczUYq+A9mO/MUPl1+6GLAomiWF
Xg6kMyskkzo/ucLx0ZFjPYiJ0qoJMOpqQNw1aVHLWQbajvfRILGE6+8OTBVzyMmZ
UH/i+ed7oTy/hrZYHyWv+4ycCsEVvfl5C7ErTVcfKIeOF5PExr17VZFPoQ/1ZNxK
Cqg14NBonh2GM60YOhjgsjYkD0Pf/JT5xXFmhaYS8Vss/XEFSy7UnEvRTjWwE9+U
uY+bhhUM4e9rdskgkxnSKjN4OyhV2QiYyqC4IqjRKozKHB5VOv9tkdh5rn4fi+hn
H6/iHLff0mTu3n+9bF06dSwK+GXgVXHTqOmVWOhWAdme2NeXnplNSmiaO1Dcldtr
BQoptJyadhwPJnKlSd3QVAavXO6RXOxLexZgLhxBI051OaW1T9amMa09MipdOvNX
InQkkyG187EhiRlRj98XRvz4ARdXykMHqGm5aql0Bxah62tLV0sgPShu/YrO05sw
Y+32yYdVWbfke2AZfOqT8TvkIzpJuBLTk2lqfENFGhs/5muyY8WIAfwnj7zw+iWn
Ly7Kl8pmGoJosccP9kUIYSEBTRpBcfbGe5cbL4ka19ZvQtqJR5KfMupRP8MGN8tb
fF2DPfwhuWIgQsK/21M2Tr2OTL3bvMteyuFUsSxBocD292ocE5zsRnqySuGbKSCj
tNDj381bcq1z4G+qbiik/FtCoUkl1ejeG/VXp9fEXxOdVzxWx0fFu1CV5DZHLBi4
4dJSiaMz+Fk1M4sMeHZ0rVdyGkixRWNhR3J/AmVeCtzYbU52c53oZ29DTbvvamgz
jyuxA/nmJKpC7wbsHlthA3DgWKvt3avYHYlrMXIdP3j3wCprD+pny5qxOoT7QY4m
v9JCABLeS+XBCcxNeEAMf/qcdvaMAqsZalhTOlwka4RypGNZF0MGhpe0dv8/RoEI
dYHpxkpmm++0e5k671n7OQuGnF2ozCPKLiqvhZ4b6ZZPt+HrhTW1hMASm7XZijDZ
28QFcyBh/UoyyU79tmTKkhkqpsKjsxZCeWLE/CJO3RFk3V/CGxTDuQYsSUWxvp3l
+k19sAuTuZ/kcSjCN4mIlJGlFmx8+ekhp3ezExGt19AqJJdKzSp4Lod+CKlwbHrk
To2ISVxPX58S2zzGZuf8JATpT36yAumNzxkaGILtbgpdZWnqmuVondbN/mYfrnsr
ECaknkVDo845AgT1avFivPlkXMlteQJNQVIhnSWm+Yw9X79/gKZRFaAE64RlIlhU
BbbCzb7ToxdlQgjv6GIDwoZBpKGb+6j/tJIuQeMgs/LIj3FHPMjQC2YZsPgOZVoN
wnmTaZRcZKHmqAwpGZ5go6/41Sd/JIRN7qVDbwhpl2lWIYsZ74eceiKZpu5sdxot
HrPHkUvaZ/H7eIMh+7Dr/s3ev9FcnWAsxKkbrc1VmuryAddf0b22nEvmPO2bTbpM
3raxqBrL4gFN4dDZF8bavLq6U6S4bf5bQNyAPFBnmJ6UfE91je4HP8d3woh+0OFj
E4W/SRy4LFb/a64zY14Lwlt/8QlTzKrdaTXHuG14QWxCr9ChgMNsMxRi/kvNcoam
7JOhQYFfssm7SpSV6tJNY8QIRmsEAi7C6Ldp10yiqjeTBVZW6fMCdp0Wz/m51XDP
Xpm+FAr6P8WtSTKdZetZXV5lVjt8We/OR9s8gX1XC4547PoAxUKtgNikKrZBekBE
peS2bSwfiSd140G+RvnbBdsC/Fgde8DOeFFxvlHNndc2htJvlrmiF2To4ZeGpW6+
VrihId4S40QN1B8W6TcbNvGd92WF3q0ZdzzO/FhUEf1gleqFNLs1DI97YucMEcOK
BOfmsdJzpRornd2fdxYMoAz6zVupkXMfK75aiJ/fK/ayTePRdernCmdyt0A93a2w
OmqhV0jOq2bIeptSawqInCpiMndeYIzO6J+5og6DfmfV3XhTHp6CBXpmBq4OPXZl
UT+wMUPIJf3Kx/UNv4fZ2zqZJXW1Ht2pTdQemEPRjh1od+iYCZDJLIBKu6sLbqlQ
lJGNGe1uuoyxeaRKaG+i0Lo51HWv8e6FP9hSW5lJN67PGfsUEC0EZsNuxeeK5YTk
jLuqTfuHIo7ViPpqOqQJwvCoHron5JQ6xVU5GTQWucYn0Z+EhpKjNLxF4foBMFvY
TYwnHFPn+9QWkBUFsL7SNcpYBmKmc57Q+Q9L4WmNWoEcZAIuiPFqVv/w63o1ApiU
eyG239pAnVT/RikuT/6LmKSSCHQ4Vv2NqVvuvL5RL6n2pg2JF11eTPSVSFl+PFgS
up5LcZjrQaF4fqFZJN9eoScZPtjMTyFO3LgpNzMie01KvKNfTczZuYNyphFUkGa9
7YuAacStmI/TX5PzoBBCEyS5QXVspeD7QZY+lh/fNygLOElEfW7kFHV/evKQSJcX
2M74btGtu3KpN92kPdjJiaHsM4kO+lErozlq53011kvLWEgWE7j2mLPMKFb19bUB
HdGwI4qYP0Lyx2xhluE0i+aly6wU3JXna5tUjoWTJXLzmaD2l/F1M2co0jV5nPpp
3KEDBAz7Negq4gb4oRdUTLeeIkekwmCVdUP6AsjdsCOJeL16SKTza8wdKtIl1GyT
dpd4yMbEZUzbLCuOoMo7TCaVOU6AuR5B4fPl/Ky+tjXfoWZQSjmS/ibnroDFxpBL
vBv5qlGnZTPhjNJBTCVokJvkZEuqIFQHvTu8fCqKJ7AZ2Lwq6mzXorU9ekGjgkiT
I4c0ZQyNBNRvCbGDRMP/goit3/9xrXBLWtGU7XemxiuzI4GCcZr/0NblRrzqpEPW
0ogKvxlZxzbYYmkBRGoI7tBzgEAWCAzWN+llPgT6Qd03Vf5i6wvej+5wCMKNutS8
hsBaTIb0gcYMch4M18NrL9TQdnHWoPQayPkiB5o0GBwaUoUcgKGjXMo0Y+4n9gvX
rbdP/lyxmdRSawneqW5rEnwhKzSyjKLuwAQUYR4BlNyaGcX86i7Uwl0W2Oqp7+Pn
VS8gYc0pcWHHLKvoM1wRRIllnFfmnpvZTsD9thmwLkuvdzCkwKI4FsfqP7l+PBdw
tBESKjXsdP4IUUd9+Tr6B6Tydws2uFDGoB2qGxyW29/En0Rk9YnSkinCSNpQznfR
AW6Fh6FU2B13itqNsl3jxdJMg0OrYCOEUMjJilvhMkcaHkoAXAYpgRlXVBGCP2wJ
9BkK4a/QzRRWqLl/c/mV8pCC9TGvkgXCdzsO5hC1XChehJ8XBWlAmgzJePVO/sag
xnQHQKAg2dXArQLRY9+3s2qKt0/XhGzFx/iGbtqiFExtI13ICyVTUNVjKlcjp+mT
JRIdTt9lzpyjU0dcR/AAqFZe4dli4zpsMUV+pUg5u+vJquQcKcU5EKjQPJCpN7mN
RyUORMs9CKJZwcef60BWtvbYqdSmg3NKyCt2qEiBU4J2fmgpY3s3HL2iPt8hzFgq
fLotW0Aas9dWDJJ71PvuWxhZM1k+Uq83N/Et3VUfg1r/U/E6mO/KQutYuePbf6im
sGwy4kgrC9kCkOWPm26TtCES8LPqCQAB4NiZ0kg+mwr3Cy0eRik48EXuwRiJp0A4
8tXp7MzFmvb7H18GMq0lv9ruzb9TIREasUK0TdpyyJF7l/Lvuzdh33yfOSEJ8RzR
5JOgTtJ6PJWU0kN4YYFSRubnpkyKrNj/Kn6NdSu5BXpVqW0J/hrhmluPa2HO4cPd
yUz6umQTukvP4cwwTKWSQjF9GY0WB3RMLAVUHqlChCZR/LLFkLxlGNuSn/V8dyWt
xwo/UkfEQVeHDNhwbctHYwvZ8a2YPnZ6b31MTMVZ0bEiDfxY+JYndsArGX2u/jXT
tyZGbzV2x6GTGPGYlG17269i4lKx7blEI9jf4dAOBTNz0Tfnb4e7PUiXL8nZpLA7
1VRuaNfPkNnsEOTPK74r30RrR5U/SDLhbOD96cpAT0LYrADeQ0aC/CZDQqrQQDTt
0rAxoVPTTyKhDhXL5gfQFpmOhXmbAzwYTiN/w4ed66OWWZIgK/t8RbgMXviKU2kL
JvnmV5bhf0ytUde54QrFysq9Kd5o1VCp/2f9p9A31MGBXmw5wbLzkDKNqz+vRyTK
CiJvhxiIBNSndFdZ9DxgjTzyoqqHq6X5xd6Ylr0Kw7sTWEHPPv1JKdgvfyWPzDot
ON1c6YfALCVbPaisYNJwq0qEKYlDyloWFaJ8L6zikO8WhtlfPxtsRYaS1Wnk2c8o
365yPxvrg6bLeCVeLuCSsDXLyi9E6NPXdtpy+79OAJykUJjvk8qkWb8N6nofwjZu
cCtGpRxDe2EJe9xO4BAZ1kKluN0ftZYNMhOu+LyIhzl0FitDPu7OesxVsQ3DpaR3
LECglsMr4CxqXGSD8FRdiI7sP0y6dnC7t5Wc7wUoKyfiZWMZHom3f03Oc7lmcZXC
zI8/FWyBz/uAPskDUGYvouZnR3NIlsuyGtSdMKV2K/WTOFvgwaO54IVlLFA9+Gn7
SyVI09dUB+A/6YVLje8waUNaGvQgIpdp0OPh6vngnhbaUO+FUQJphmVhDH4ODYU+
1CfZspa84EtaDoqnjpDXi0O9nAphwIkh2dqZ3XXszGXwuNHE6vs9L0XWUdPdMFSK
NXWngCPASZwFkhUIEaLsfMQtb1D6Ez6AfU2+VX0gG2ouisljFkfX/DFrek8Bw4r1
GmWrBAemblFNn1xE2qLyT05MpCXPMzUO4B+1l1ACu8WlHJsjuVkzDqVE+E0+3nKl
sAvOOVLtcD5WS8TUDFu1PhBIdSVusQMGwRutHDLbWHUor2CWiSNXeoZTz3pwfPk1
r7Mvk/kX+i+0bJgupS4Dh+MwEIK3wyyYxlwtTsJYdPk2bdBUao82g7WbZcw556DM
zA2CtDeLmA/SW7G6EjTvA7tKQO7pbxXkQQXXOl/28jsqrCWPDZhi8UF9DG2ynhxr
lDauJZK33lJK3QaxKocniyuPbOIUazQPkQ3WznIhPir0N88ye8HQwAXU/6BhrqDT
dm1d1VdbqVTBYfsU1KFX3sq7iO4RWzhK3NsU3W3bdYRNkEH+5o5TW/N8nfSh6bce
NQqYicwMehKfKU7yZV+OCH70Erb/PCtjECycm2sajraFddPwDchverlmvzSo42RA
SSFh9Q+SiGE84KLBQFQehDWw3YMI3xGUDI/LZm8WF9ie48FfNjm3jy3hgukAl3OP
pbydOsDG68t7ksJ4A2hvnBDGhuseNcZ3slcBCNZnJXOTdOG4dPDF+f9epdJ1LYL7
5PcdGJAzXOEqX9D01zKLHfKbHCl+ZR7k95UL4gu4MibmAqeYMCo73R3yO/onp3vF
8bq0r2ZJIYsTIWaP6JOBbMiXtomeyJu5DgbskMut1Fsa7r26VLLPKoFlbS39WOjf
UWX0PtNrht4AHStSGYX27Z+cnDe9s6OtrTjd1ChHnLH+TuicLIwal24+s/p5Vv7C
Wl6buEHIEaSNg1CwQnivC+n1jeRCcWs8iKBkpKvKcp9aJNrMCunIbCjG6u4B1XTy
ZeIWpGP8wj7c8kXJr767DX2TLYdG0hBEG0Cras+I19Mcy5TI++Ttpm8IQGSvbrBD
g8kPh35EP8+yFgtL/mPOAD2lJPDGedMu33vHokZ0bkOpfx3oflMdfbI8bO2z+VzH
zUBOemfqa4UY2LQ/lZm1Vs77zDgLQ6fAerGA4wlCgmgf/e4n4b9n8VZlqHRYTZiL
wgjAHn4oYMHSobtLYTV8hWLlglrfGAGMDEt7jliUh5vj6IS0M3zhbOoeuw5Dp1Ae
bHYjq6S26IOUJqkhbPEidBYCg+AgXVHHJATMVZh7M5Il4Kc39nhuq8LKMKPtk6IK
IqCPoCN/FtqUDLJfiuI3qopnUOD8agbgeva2xvT7jXrs9LaRi1yyzV8G9r9jpPJ3
Rn/9csPnhdnzJsJ/VL1kftQftYqVhkdpB3VqSRZZbBvBoSjW5X7C1q78coQcxKIT
4VaH2//ths9RaEX9PERTkO14C500pEbCp/QNa3qqJMCpnW3rW+tjcCUH6MG0d1Aj
pnDvlojj7AaKG8hD9YMw1ScnUsXdV/DvxoIGhpcOZqHWKEAlsWB9uHUL1AdNd2LB
QPMAS3WIInEgxn+jqS9LTdtxUAcxedauiNmDw4arK0asGNVcgPkzksZb8JpBV6kD
+onUbxYzjGsf7NBVAwGNf2Oqq3kx40G5XCH91iruqEfsMv/xIQiIDUY1wJ2ManZt
mx296bKZZRNQdxu27HLek/j60nMQGpAJwZ+NjRBs35p85H7V3g5rXnGDS7Mnr5q0
Qrf2M0yIoZkzjofL7CBODtxnAOMhcDaUDGWTCOtHtMWd+uS/9yvYLTJO5PWQbO1I
N44/rNgYGQWExIoIJC08Irrxg5oUJmB+CUZ00YAiY/mAi0xQfMolEY8ZfirEqSaZ
+etpUrlXwc6v2B8D8xIvJLzCqPMJLUd7ZnHQHlqfRM5m6jVT6mDwsoD853EqKMy/
aGs85cXdVtBzntNc5tcDB2T0y3PKQ8Gu7G3QYS/2s13JLQjkcDzAqAxxA5lDTnzb
8b6kfzSwJQfWxhlBws4W0mxQrjzyU2NeVk2wmzPtjZH+vEBZcF1l9NlBPunrhYim
WN0uLot8PmvYFUMtUPTKvtxZOf4f6/rRInJ/SWI7n+gABCY1qWziCN3CHjujPz5e
azuwoIAWywOXUwLsSoXM6sEDVq/FKDwcAn9ybxBABby5RcnPeAhBHVnp9S0GOvh+
xU/nUCL3YVYC1Bjv8ru2SNP9PNvgXjtEklAJ3ANGq52FNVupPAykbta6b63NePtF
CSRYthUoYdjjAjv48Vw2U9ZxZsOoL65vw6pABUxc3YM9bm5GCUVFlH1R1hX48yyU
JbC/m6X3lGO04iYbzvy532M+xmOWul2/vpdg8v9+sOwmAoz22IKjspglWFgVem32
3cStXBnGsr8MFsdM04Q8M+7SMmOW0rhpOp0hPHklDfUTO41Ex8BONFnAAyqn+Xj6
SkMz41zUHYd01SKllVVKmvF2utYoo5I1IBgm7hw284cqVctEmOBvLyXgvKSTDcVc
rYJb8L2NNOihao71HveEOsXI+5iKnnZDaPuWsOaTvdnf26P3EL962t2iWZ+hNKjw
HnAzZPye16vdLzh04RqMERDMKlrqk30V8okKqBLCz+F1rQUmQk9FXDBnp2YWiKzK
KjFpPt76Y35nJ2mUgVejR11vb6Fbp98lu6Zs/BOMAz1a+PpC+Vat072v5SxZrbeK
WKgbNenIYUpBDo0b5N0uLpI8WAJ3sUeI3mSpZ5SRBhrd9ZdMuY4mS5PHV4iDcS7F
thGeTeWTK/uWTf383l4GRRAAF9lJklCia3Au2xTwwVpLHgRagFLPVuhWS/6M4SVK
xymXdDTXvQlx+l59UiAWMgYnS5HHfPe8WGGq+LIoEJK3P8OFZUBL+nXQHWriJvz4
bKnaeIYJQTFhKzI4MZXaaisVdOBor5uizrSBQEtXIkobrHN3oWYRMeqIrgAN6u51
ZW0wG7NTvw0mAuK65eHbKqeeYazJ48YzORBvSI4HaZBmbPCwJP4GEj6St36hF2Tr
2nntavHq6sY9bOhWo8Y9NDRz8k+czhUgqvqF7lx9//s5P6tbRA0VjyNM3q+pHyb+
nMqewWS7ohxFPCsDMfBBjwbqSJo5PB9X/vWmfRbcFaBHIOXurIAQ9QhebmZmC9tN
I7euVQgegWekvx7G0Di5LztrKgEOTc1aaDn3MtSsci+Ke6ItQ/1oSy6L+vw9AQg2
tjUvrb4lBU5KdlWzqnRKx+l1LhrDz7bc9Z1BrvkM8hHwH8sf2wyw58jFLO4Lpoma
Wzk4YUFn3Eh/hHCTgXhV/XlRZ/YrhXT3hXZk2veJCJS4lNRfC/3dDfY1KSQBs1Ga
44n/e9qEya+jPvSssiJY+JvJP3wZkFNtc8f02/cSQjBlbrAER/9GuRGL92UeHGQJ
j/mJaWjS2LCdzn3zq7eejQzQnJKF7p+ibO0p0gbOqUK6uJ2PgXV7CfF3o8HlTxA4
9BVMhWzwsj/D7RhEcoRGMXfrC6GRYSNCDdrlRUBE4u5ZNntzQhQu8TvfEO5wS++x
crAlgaB/cqF/EwgNFDUBIckolu72SVUR2yHtQlCGey0eNbC+nRziDrSumpslnX/M
vdKmkQcJ21SIh+CZptekKiKgx1uFk/T3brooJRv1aF1rPQJTM7jwRZof6/hxhM8N
eC/g1RwOrHLQys9+e1QxLi3V/Gtnmlta1FhmkCpjsvGUKCJN4TNrXnuJfiCqq+/l
wHdKaplhokSb6/pfV+PheKjnqgyaFSH4KehX3POiWQFzUxkEIpjAHcai2AWjkkQ0
lMMqc9ZIdDXK9MnLcsx5cKZKhr/gjEY6ZfIhYXsYZs5GZRFhnFdroVWlJ7o0kqrK
XayUj6lEK8btE5NCJMwYsdjRZlgZl5JpY4HsZ+oDR4C+C/wRxjUr95qJKh3o+1El
LQsvUkKrzpE9RiYiSRLYNZYbL5hymat8+t7k1j9nQOPDxO59uALn9Dun7bIa1Y/6
rpyt1n94iwZUpmlulGAAMsVi4nfIpTQ6WwUCIUfRljv9UGD2qGXlkRzXobR3XJOs
VkEUDWOtWn1UXJWjQs0MVk4oF8eVT8g9rvHiUPvUUdG+rpDkKNBbUdO3XmnqcygJ
GgzG9/kRigXhlPISk7fTz4Nc6tf/Vg8RW7GfR9bEWeCB8jhzUcnqmch5tTeVfzrR
D+NEBVY+RjowerYgMbTvj35HYY6T92+Zi5Ij2TsrwVJ6miDwJ30/gZHVBn/uz8A5
opvXToowaVqi/E2SHTwGvyUK+QPe7xMnqHn/njetiT9XWW5eVlOme3ggnT2Oin9O
DrmI0/1OIyXjE+TgfYM3rhMiqPuJheFHex9y59w7yMpxKlagrsvqw2ZmMSotkHmV
8zzKVvLJwf+xPPrFULUXwTTotK+OWC6r6q4S1kJNi9zcL/Buq+vV+wzWq3loxUGA
vnXHZlfiQqDzk9PJjTLs0LT305oCxaO65tox6E8nYhba54ZSwDrToBKEYuEcGdkl
i8C+F7+cFKGQl5kN51i6QhOjrXhjmdQQbXUc4ES0rgBpIhKIfAaPn3vG24bb6mXF
lXFAkU3YeTy/kGZ1jqWLo8VxO2eQJs2ktYCyynx9p366ps7T+UBvhCxM5il70S0W
1J2H7ah0/0ZrBaZVlDs878FMUWpezLH9bG/g8dr+dhXGZETXddvSYuXslhDVrdxv
+fCC9jHyG95U6FfA+4ojl75C/cwdsHk4vxNRRb26QDIJL3RZasKHgmw8223SfKc/
8svVzKfsN4wOl+Y1kpQ0iUPY0ihK9LrwxCZNVrmcMmRqrhQDm6nSHreYiH1xQPTc
beN/NLZRHx+MFl0MpgvdzgFwTKgR+V1aIn7p0XzWxhHC9WeYAvoqhiNE+O2MpyDf
dAGvDEMCWsRb1X4mNsj5LKKhpLv+zR0vB4sNo5h6HlAAHie9iXC2ecUTS1G4IZDD
bUxdi8zRwWTV4QMqUNw7sBZwdLZKvIM9U23sgrTYji96RApy5UlTdxc6t42AVLVB
1ETNxit7OI/3XLMq5s7bjkIipQ2hUzUIWAZVzBflaPMyQBMXACQyEW5zCr0JNG/e
UJfsaiDxRvNJYevjVfWj6iyf24FohLCr8J8pQP/F8WDgVpIjUE+q07O86A5JZQBN
cGS+IO0mcKlKKPcJ4XES0U9vhTcVZ4H5OIF2sDCGFYDnoEDEc9ObSkpCZ3wl/EMN
zGFa74dr2R7K87h66gqxB1LjIv7LNsaDRoqvBxJtnxdNcE7jLliJbvKCtSwb1Jez
xACxW2ZVWq8AK7Z5iKNzKivsZ9yBQYQAXMdiYPGuh/R8AChi8M5jxikJetyPzIhr
f1ddewVD0UuPXRR1UF8JfIh6SlXx4+j9wrcwGloGbQW4TcLu+p8j1fPeVBTayXDn
h2uTyCpuYTWHlbcOtGkf88sSl//AStvbVnMPGJCDTDWnblEYMHF0SK3qj3D/XgKh
AF7o6RquZg3EzstpOied1sn1l9yTCTQdSOl8Sk3ki1HxFFqlwqQ3IGaf+3RgoWLR
xEcUtORoQWPwuiOKzImJP0IpS4c/rcZjGnhmv4PpZeSPz92JYP7Fj6uVbSV4z8Us
R6t+0BgaHz49+6/3+hLnodrhiFocZNqZ7PN9cJHO4S+T+qMDBuWCwgAvYZZlCjZt
AHfuLRLkNWHvxZnZg/pWwha7uOJWKpw1b8Hp73aPY7chtbH6v+CGKttISI21Yt+S
tRnyJzBIXDKmD2bcmZpvRreir8k8iujaOahyDxmkryduUD0ptjSEin96wCfsBSbH
y1Jn18yebZTnRIZrcF4QQPFviWiF8P4fV9AmSnZLaOhj3ENqVW3FMMkVelzIRmPD
LbH92hHldaOU7HZBg/45ajP0H5rWtAKxND/NgPF6c8k/RXMSEnNbL0H/lPKc4GBB
c7tXB9wR6gHljISeyQOShH1GgFdfm3RK6Yb6G7LdROXzf4a6m+6XDH7tN0BSHI/5
MNtrbsrSOeEuhswYIbGRRIN18whaUTw8ijKcV6XetuMk2XHAulJuKsuci/eo4FG2
7Br3EAhfRsLm4l3vruyYWG10jZ50M9AOM8Lv5XCuj16E0bRO5xSdMIvaVa18mrjA
gwJzkZRYAonSLtmWquC3LZtLLZIbppPeQ/dQjxYq+NcBpoGtsCxNcTzUQhcuv2pH
XI64VcLMRyQEqE9aoJZW+A6qxgL/wvwSmSyIz+E29USqloXQxXYNgmBumHFrlnZ1
BqwcwkXsuDm/DCZPut73IOC/Cxoi7VpXDO+veiO6mX7d/I3d6oKa+kEf3FMO6hOy
My6XrRL1YwlFvAEr1yaFJrVyN2qKrsN0rw9wFXayx0+aoxXbIZ+6FwXfvmgQJR1M
e8DEnBRcPbWG8BJq3Sf08ZkDj1ZmyAB3u1qlIF3qSxfVC26LTN9dAkIXTVY0bT9o
qelOJZ624N2U4zk/igmKaeEDdkuPIFzihCdeZd2q2odtLOzPphal1XzRhzxrd1sx
DNYAGRHFUySpKD+aE4eaZMu1LL86kS5Bd/S44mQT+NBdBRdrj28hoBB27wn9AR2k
Ev4w4nyd8vPlQDMu9VP8n2UD2LKkiRwCF+fmkOnboUlzCkA89Qd/YINPkGnelQYU
3zfantdZU8VAPzF//lRAcJsOZdfi5Vq5DkqC4gpXkEEAYXo529dKMV3rzkgrv7NO
kDcBOxqXZ+gYj0c2tbMRhNiFBIeoKBn+PwtEW+lBn7ARZOVfmW71OeS7R8ehmgTo
YjiMOcXGqjx7xUVYM8yr2ZiY5O5T8eiSgepg9mmTc2O28Zbypq/Dc8yNv/hmUJm/
lL/eSOePDaP8Uq0qPwG3p287qRV7iQzxyijCePYplTErOajUYPc54VBv0FmZWwgk
LoQeTnrvXU3gdUFVPCupbZ/FXY+zgvM1szLG4nO2jYO1rXOInSRe2RqjLPtMIl75
eYBpQK/x1XgS6+R1gVelOiYLAjVMhOuTNkoqwP+AEJhB+authntybjACBhSY2zlf
lntDojTjwrlRNcNj8D56fiY4S8rX6es1Uanc5T0cfcG1PI6srvL9JWMoJTiAN6V1
p1SefbAt/a1xr1v/u4fSVv7dx3C1UeW/Jq4TVeoa5M9IP37L9PF5Pjcwr9WIwa+I
EIFVx6Phzd9dggDD/WrN0qrpYlexD6va+nEyNOhkVGIH6ZyrJncs068wPgCJRzKq
EAU9rkINrSaB03CiEmOfS/dIX2m7lcnP36lHmgFbhLxDUUFi5jaFWU+53Eru7rNZ
BeBW9zdnS44xXmz0A3xh+kCLO6m6eNIK0FDOXmPjAH+2e2ljxmrLsDfsjOaTpBDH
mUld4oy9HfFnZIrcaNMdLiEsVrZxo3MdbqFJ0ZBItQFyDY7hwDel92ZY3RMLdEd7
Bb3OiDIMgM7IShDOdtV883er/LGYO+mbilvWrl/Ap31l2gUXeG/NTNUT0RBJ25zg
qMn17qG7I/c8xOlERfx18ySBDKqgX8Bdbalri1+/2CBHJQSkyBuAOxmHG0oM6TOa
q6fIcJ0GPHX7B53WMGkUy9TH1nK1j/cWNQJQh55QxGz93yDyBSsZfIJwTZH0wUUJ
PgeGZf4ic2WmJDxVYN/O/ehKw3cXa+apCkVqof1IylZ0PxkjW+L5jWZs6Xd3yNo+
HhNkmEJwk4aptMQDSgnea921CXfYm85Kbmk7WXtfBJL3WDitTRC6dmVjKYwRG10V
qss9LKuDZBvua/fOre4JmWv2bOu+1cc4gZqpVBIrVbWPK0cZxoJIzqLjcdNnt79e
DjSW3XYVzy3gD17XDed2O9jiO5dV+ojvugvfiQ3u4+CCXrIzeO9yYy4fwirP5PEW
1X62IWgKgMUMj1BRQMc1y8G85lej0V1xBVN0PGPafckbL5J4aIlO4dOp6PZhKTDb
MvlkKC37SQwDBopJLQ3xVl7SCoqJ+HlwRhPOmE0hY0dMFNK+fqBE97qk1Q1hRQPt
uTOB2TP/6+WM+T1hFqHV1NoPFikICXtDTuhZOOn7hruhLhpValKCQGfLEeTicy7I
ILRxjfT1sYjEHXg6RX6L38FslxGVR9oRWFWNHGkKecHg6GOZZgUpryqwsZKkpQtZ
NmUHFl48cmA5GZLTQek7LuCFJRAC6XDNy109JeIzniXjNObMMJH7tF6eJyAkbStZ
nbnZVAjbM7JhnTVoNePpEtsNvtPL2q7fzFMRmjs4juGl3u/bxJQpYZFaZMa8GaRs
Y9C6FRoCE7vxk3WmMexdoHU8Y37Mtp74YXTylgYEhv2zaQV0bx1saIOKEZr1CfCh
yAYkJx7b7FTH3CnOt8Mi4IlxZGKpxqvNvhuWHRxDvnDX9g0PWOkp9XM1UUQCtj14
V93pjZwDhjNfsLUPt8t1WERO8TOrc3J/LDL2Cf6oOhWwcLuFWZ4sl4yn7E2v249/
nAnFA3ItyMOgqHZS1mFlVzBbhjbh/XBCZPiVjUuF5j1bjQ/4IHbJH+UoEIpMEhJ1
mKeaNTYDcsjkMJ+SMaObG4HQV3HSb+WRhhbo3yg/VF0mAzUuJjh6ebv1FXxc7r/o
D0pPFymnzw5yQW6o1TrbBHcBIkN9Kw4X0vgHZ4jgXDsAj9oZqItgR+Lkjbpls6xU
ivB463pzX9fMLCXPZsB3+hxdGawqhJaK6dInkUIsl52cZ7611sL4gnV6yEgVYANa
sMe7SCkU0hs3SFBwzXMEaM/sWXz3Hwf4bAhUakQ6VaJgZ1lWVwJ8eHSxqTaQAeBr
KaZp0GMeVOyMfXzUg5ucCIDF7LX00IQzlTsqcSBQ+MzPASDPrsQbTTRcDP+Z54Lp
Gxi0fCib7zUJi13rNQvtnzLjcK6CZdHRIj7ApQdqlLlgyaPNKxfSGAJAPbRsT4DZ
bdM9kMAJqo1K6TnXlA1Pj9TtZojfiX501i9w+O9fygXoMk/lVXW0fnIsM3NHnU6Q
QOIzJRBK0RrQ5x0RV5of40jex0nI8DQsirKahjP4P0U3NepobehOK/BCfNwpoYhD
aEKyuH9VT9KE2+99wlfmBcr+gUSvG7xPd8cUJHztU5AHtjX+ZpeaYmj8FDlLVv6O
ziubMDiRugYqeUTlRhXU5GSOE0aN44YOu1Y7NhY4Rit+7JLfqDF5t09NEpNFBjtN
Da8ifo8H23cKsCWPZ0wNX9ndMllEPu2KackuLLZEeMjN/x6Oucrk8CN8RtPk7c1f
tStkEaqVpShJ32NFsRGzFf3TDwcUctrdT/lnWvxtXKoEtaV9u/a9BM8I/i93nhqo
0pLwQKqRGejTYAC8JaUsyhoG21+DgzKcfgw5qwjJNMUwG2FMMCrStGuwAbRfGBFb
NIfeN8lBDJrkk0l8LubgDolmDJjBS0oHHQBAehzCH83FUgMEWPApNE3PRFEVJzwP
9PclAzQAX1wzUbwZeJhfyFSguGeX0TCjIieyTjTOvbQiF0uX1G2cLAQmzLn4SG9P
+dTFj+mRL/2wFuNVeodDvfcHkxV+jwU+8yKliWK2I3r0Bs5rkpkEDPr0HVL4oFQ/
+7Guy3vHh7duAP3Tw19C09hMfUfEjdWGNxV6G7+gFAnhOwdvn8+N0lIAwgCw94q1
nKd0uzwwJfiXw0KHGB4yO8dVm22f+9pmAgaBtDIH5uoiF7Y3hGlg59wQquE6IpNn
mkAO6ygTZvsPnkLbRlUSmN45OVVXUNIJdm2uIlzo0TG0PE6ZiNvRd6VkNwDvuCq0
UfZ3VQt0yGr47iyBdIXygW6O+1EdVuMq13QiIwZNRinmAMEDIxKlb5XOgN7FeME0
eeATEsx3TFSnkPIokvEDH/wQeqxHUJAHgeJJgADYUZiSTb/1BYxL2NnTY9qjCQoX
66zBsc3nPbB3s34R8wVv/xGAOsEcnjhZl6kXoy9/Ia/FirXVjoLu10sQ1pBaYq1Z
WWmaTTIs7FHMurH7C+OeGm8C3AURZBxqvK2qQ/01YhReFhdDY9hDHQMnIo8ZuFAW
N3USazReVuD/pEhQZ9Sk6RuXhdlSYTh9m2rG9vvX1qT/F6aARv16XDqd2dqKOzxl
vJR3jRIX9eGKbRUFyjI2Cne/w6KUZnPfTUSFUr/MvVXGaIlCsPrSjSV/ssvwjHpP
X1QiqPgmIWNyoFWq6j2vEXwATGPoEPzYuK2gnLI836pV+EmuhBOnkmlWWjG9/DZe
+bQys7R8HEKZ2hPXLGZSrgB3CDT/B5X3aflkKTdhZFu20gmD3D6z5S/N7Nuz1WEs
NDt/uImkIZslV5Y3IWZQ9sH4MQM5S/Gah4JRa2os/k6LmOmYBQbFCWxV2JnqG19r
0jvkCkdK+aPU052kcxDG/TucZ3f03gCFr1EIVDHohjbcIFUgYUCD6OePuiW9TAOr
QqSnY06W7aQwBqTeLqtYx8ZiRYdkH05Vk9H/C/FNVXHjq5iNvAgpLiO7grfRpNZP
MJjZeZHwkGG4M3FME/QGvheheNeqOKkkBCl3+wtBbM47KXUkKJYfhL8QnKmcthaR
F8qcl7PXi5kK5W1e6oKnGWghL2HGkL2PLyZBrllRI0KubOXeMkHmP8Af5zK0vg9k
AMqz36c4e6jJj6qsvi3wOS5vlaVY4iSZAAh4BbvIGnLCxlillyJrLqhesYshc+9t
BUhW45mIUBwx4zNYNdF5t0z5LBmOfmuPk/Mp3ALnrP6gZGXhnrirKlaw7jyRuT3X
fwgcqmEUjSMc+GSdiIZlyjmHdt8U7m6LR7vq9JQ7fIVhXglr7rxRahLo+mb2d+0C
QldhmlVK05hCPudhlX249lqYOYtBZIAh6dhiPNXor5CmLvBzYmdq2JKIiFZkkIAe
Y74Hvp2us8NW1dAWupsehvcvAhSkGEckAfBBaWgmJOZbi/pQhXzp6D/QSzgGeXvc
jOjaj9CTZAYdT4Uipr3J/AEdO5GdC7iGcAR799QI7B4Xk7JexQj3HxiBzzefp9JK
Gr+ksD419iqPK6rz9xuNNAA/3/8c1jZvsMYUdi2htajSBqfEsVrD8PAf3jhdfqyO
ec0pGPkhEhQWatObe4WFSTrOCjenfuB2hzFPQgBhL7E8UYpxDOTu1kXM4YSkCkpF
39AlCqVrDWqV14beiPNiASZ8AdXBQ4T9d7SiRylmt0NXPCKFHfjkDTvDFA00YKwV
5oZxNx6dJ4lvbsRHza/J2maG/c02t+sT884NF6FnIit5onQDEjRztTUcFjKxNoiY
gURbICz1YVTs/ByIEKptpniG40ummUmqVofnSRfJT0i+3MRF2Z1c8SSo93lc4khX
9EYD8hq0n67G7EGx8B9g3Fy5DpIv5CovkV93PTI1UUIInTIjXKuVI2jrRQnSaUTG
H2TbaDuejWbdSHh6NnpAmove46qlCG02hzfZCQVw7E2m4oP4WLA+Frechq0sufpB
5shEtzym6Phxuf0xuqP6BrXW+YKu6mho8kf+zH/D0nsDoKFihtEiJyw73xraZdrP
RIe12eMNx6NTiuQz/rhJJCp21Yhw07Gh5YtE1Iedm2tEDqEZpEYKi7Mw3q76JKkT
SNv5kcQOujD9tJ+gX7KMrWAQOftUcjD3meoBR+/Q8j9pZJ7w/XLDLrlim0PGN1wA
QxmeYJDnHjlS6IVrw0R9irRll7tnt0UODJFytHVr3WIjIgf/WOmQTwGFFE773OOP
Geprl+N1/OFbKBlmf6rLpq3k9dwYaLtV2fSopDUBXtV2ef6zCSteqrNTGWjJ6p+U
XS64o4bZtclkE6/b4RZUM6MXF68B6dOzvgoGk4kgLGKCYsjC47erjfGiu7GsCdGn
za0bRbIPtEMby5Yqvmj8Vhq52wm2mROUW9Uy3pW3ze1xpz7M+HgXMs2BWjRArvbX
0xPv3M3NMzzrjQNlw2Ww4REL3w4Cro+/v8VusnAiGFKrKm0Fs2dbcrhu8OLpycLR
ymXuZC14xcJSX3k5FS0gqsnkZ1LHFEnCQ32HakCXJxcptbUJ41IIKg5qhMI656rd
PaVMAtFpY0QhgwFJYnC7nMll5CpyiPej3X48rJq16VSN64mFWumKl+JaYOQdMI7L
nZmPjvIaH2tyUvncE8tq8OaevPGhaFYU4YYxOOcA8Q1uwKEIacryxHnJp13GAxR4
BJ1TOGekv17oDgssxIUXHgrHA19UatiUYGTKQt0EfT+1hJg9kN9k/4MiDpQ9Va8y
dym5O4O9cV5hdByVLLTrn38IL2irFVQoqERC1jpGZp+8jFUZMBlf6/QLV1PWPEKL
FmT3MHTC8xAVMFHwZjOIErcQgBJnlZkbElDymlVAGxb7J+EaQq4fGbWmybiB8KcS
NBSqKQ0lO2GApAYRpE9lBln6Jpi4zDHm8OcNNfXzEOgZgEkTeyVIiiIWoCz0fYuw
ECr9cxZ7ZY0dEDExGsEH1CcmFJ5TXyEjmYaIenJrj5/QlouyktJ/tjaxHWp4HyS8
FI8dB47ZgiKDH0L/z0D7LdSIgSMrbrk+z0Ii1/i54YnejjlmLAlepMvv6OuoM4S2
sHSqalimvgdEq8Oga6gE7TTTLaNQcm4kDf0L372o+hrC3FRtKC9U3rlgikV5H1t/
mN78G25MznPE2H9iIA8Tntxhu/W7wn2mLgk3xWpCnF20NxmQSt4G/RtMFcz3yKg2
lJ5cgfVjHF/Zj0awYIQgj1cLEEYbLaEtFf09x+n272wEnlwk75yq2iD1uGnQuPoI
QnbgtB+g3qPpyL7KdvTPy9ZzvTzegkDQLh0lLYG+8niBJRnPQadNPJv/Vkvg0MYy
Vb01rRhC47OTshzFAWYAMxU1PCGpHWmKZbKyKWWKJcE+MjMwSmkpBhhihRGV4Bkk
sdUVooJjIS7+akYi0wqhyeBw3jT5JvuQB3unxOieJvmj8U569PMRM4ZEKm1bmRIb
O8jQuU38AtxBTtCqdGXKUKidXBrmlG8EOyQ7FiPi19MFPmpnwH5DH7Z5/uhz/r9b
C2lZqXWM3wOaqggcPIXchkxChC132mdJ8hFRjZNt5fQWUEXMn37AArCleIXbLYhS
eijorvOjefBX+eeyRtQDJZRB+6kqmQGt05U66GpJzluB9tD+WUyYE1juaFtCBKh9
Y+JWMffpw/fbDvpw19+edGInUmZPOYETlZDX7UxALFNMPpKAk2gf36C7Uby00gSj
VocCSbPVb3e5isiMMd+ppxBR4Z5/ZY3FS9C7n1l+7swQTfcT+hw00qWPWeNJXG+o
LpQeROy6UQtQ+vkJ2DFGyVEpGI2WKt09UX9ZWFgWA9CTlm+aqjc/uUD+O6703bvZ
bdVAztIQVz+Gf5LWTAK2TvrD0taLM0IvIbZjYJNnZAUhN+K4g6JRKPE6KpgpmIC9
BK1XUMDgOZaaVWu93b0T5ptM64aFXKKj+om7HHxRW/DxV3JFx1VvemXJ3R3Tep2y
/8/gZD96e+KWdUitcNYvmKj75d22nLN0BbLD8vfgj/SNE5euSfp+IfVHQhrzBFJB
3q37AFmOPidM2Zd5JW5UDPYSThtc740O6w4O5ZzwUljFGGuIZJ+GHMhzoIr2BLuK
mJXIO0I7icXjkImatkAXq9Long1qt6SLCgxyXhY0VvklPtxzHplvp0cM/HuhLS9U
Hn1bTgdP11zvWKndXAcp5KtJogNF+acLGLClNlpLuovvtckw26rYNITR92o9YBqY
nU88EZ+Iho/NDwX1+vxqwSgFm86j+528lW6ZvVfRSIDEGzZwNRRM1dXxTKsRNADf
ph474A7CRWdcPJKRZ8uAvutxjWsT+/DG+y1W032WqEKrl4p7np62FYl3I/vH847Y
HB771EBdBBE64KHDQuaEcR6ZRZkaGd5TQfTgI9iEPI6+YN1/jK62ryGKnB3rMsyU
8aA2WKXhUC6rjZedO6qta7N6uKvvm2kYP82Y+9n6KnGLg0Ux0m2cvZoHek6KarzN
WbN9HW+NlXSl6LCMHigNEJ5AsiccUmY6LpJKyN1Xi9/h9sxC94sfJwWacClkOBQm
87xpD7EgEOajTp71F34mMOTazW/VC+sXWSZgBEdohdHMo9TFeW/pcwjR1OU7R6A4
muxCXWbdG0s8rESZw6yMGWO+qGcYqJ1MpgV5vLfAgdj2xqkeVqUH8nQDL2EugAdY
PGihR34EsqIOuFlPznA8x11X1gEFV2+BDRs95jRuBSz/nsmghGHq4BAv9fxA5LXM
bZZn2IQ+IQuQ/S8saSJbLorZoKlQySihpPRYn/LV/XLPuY56DvP7MohsfeWljbbR
cTw0oAKf+e1TNwbm+V10AWo7s1RVBXkib4Mrwci1VzGcgEv/NGXVOgzoBWD/fm9z
wXJDEZ+vjiUsIURwvbzIAXqQgnnuBgJpPfjxUeHU+RIz+3AIa/63J555ENWpFme8
4x+8dBfJ/xxWwLP0KKsVwOoOICbxnOW3tXb4+u9k5gAHb+di4nUxog4GB3DAruB2
qWbOrNrwazANtg4FY9PLfMdikX5aAUT/Qe7pjFINLIwScye0J/nUqh6fb7wdZugd
RlOkNrW7POfHYotabPt+RJ7I9VrK+OsTKXDZFPHe8zB7PsQS6BXjwAVDQR61+3+6
hRPp6sTS9Fot0o1h6Wk9+fw4XePk4VoY95GWgu25xL0mmxzsnpCYYZt55W6/9prf
HJNvYJW1gqCxqwrfvhBL97ghwi3fFvBJ2FTSiHoephbGRdg90/dqPqWjbXDqUcQf
HFp1eVHnLbyizWigAiPXLcmF68yHT1Y4kjLESpWKXpANET7lc4deFP/OS7gyXRsQ
8DHVxVze4SJ5DeztzVEBVB/ogC4k0KZ7DbEZPm+vD0YW4I3hPnQIzbmG6jGg2Z/h
Wt8qauO07ptIEMJPNx/8voSsAF9klZXn3ZGbt3aaMhfEeRtFOI0O98t9EFjKL7uc
KDMJeqsypSUXYEDTuWkWXlb5voHpe2jbIBS0MdwHHNo5aP7A4eX4YMPVLmavxTTK
ZIPePRiuiQzWfUTFIETty4gH5GAT+yQs4cRBqh6F/Fl7clgtD74LTnwqdbef947+
aLNqwSVtSf59sm3rZ6cDsK4y95zge6462Gjn/vClcnXK+4GUv8OAanOqsPedWYNT
j19gj33jsoFF/SVLQiXXabn8ySF1BfmwA35I0aO5qbVUa97d46/nFpcKT1pFUT05
FkOnwQwCmtOJo3dY6Woah5ixUWJFXrwVquRREhADqh/YrDo+mufDFp7dqXijIHTF
smoNhtsyvXVmFcRAlhlg22z8NzPwO3Z5jktXl9IyrWWCf8AE3bgYbloaGWQ8KhwD
5OvaAxv6tg9p8up6EHd02EPRuSN4qs3QEwOX4xc1wCTYztSXM04+QEu0eNBoCy6O
DzW/MTlqyE6xx2vd+ZLbY595AJKLfoGlqSKcrE0R2AamCIKSxrInHBK/tKxaTSqf
8e+t6ehmMobHltgw0ABi+VdaWNh07JKDXUWNIixD7qxmMgDaXcq0r3wt8SzjZ2HF
LvzHvG98dFpgA4BCe1i6t5QFk2xyq3kDxVC5ng1OXvlGkVmjPjRIDNe9ZkLbdKuy
OKyf1REuuB6+qdCiD1dT91UNt2vs3PW4JbsfAEI+3/l9Gr8XzAG9kyGgsYqcyhOy
regyZAmqmC5DdTt9CoGuEJ3TjjlYlCtl75Z4Y/3hNjgm7j01rnW9fIohsGxgQpkc
hJYOyFPwSdRRhcl5orJ+DmAPwivYqCJuf1FKMnotkV9eZdC2ZaiCMY0TNV6U/tq1
tSrCHMJ8qaqKN9wkrTPZRYQqJiTtxE7KTWm7haccftFYtGB6z7IGDXYOoBnBBKOc
9lkSUExJB8iXta5Y/gOd+YtCBQ6rgULgMvCo9/duQxKgVRvZFvEHSKntKxRqYCa/
VdITExUYgzaQXlX/rXyPQ3awGHIpdIY5gqRRYRYECzfdDak9X7IHmPmSaiyh8+BZ
iGjJpJF0SSrODRUc9qAXuXOFf3m2xNeWP02KzqYVSvoHAidoWDIekG0vEKDrcWuH
M0xUpLEcLRJFsDIZuDdHbig9hKxyN4hWCSzzzJaB+UE3frPpRWZGdgQFGmCfIY6z
lDorXtGBCf2hcbUP1XImkCHdUb61+G733AHAw8k1i8WUg163VoP7XxUg3DRZ3JPK
OST8ag4sPNsq/akqyh3fgmKlrSsDhqyy+MOsYrEXoQAfpPJe9P2qbIpifUiLIV8f
GTKObfOO1UytRybkpPqTEZnQaxAUgyRmGH55+rBfHlrUpZoM/WHW1Q93+B17sHqx
MD2ypbFbp7RXvg3VJXENYL3dolJXnH8tS7ndtBbJDRSnR5o+WHBrHMPDGTNbindm
oFBL9cTzD8pSpWvKmUsimHzTSZqNOUVWsLL9FF2cVRr8brC9LqFj5JV/5h6HljjN
hvmR/GVC3Up6Nw6fszqnpPHYLVxE8Eyw11SMQXY5Kq6YhY92EEu/mRp+/iwnbIJj
eb4VtIVRi6hxWhvqPpDWyIwyo96lp50WuAx/ODRnhgu2TOBsDnVjky2luY9nst5H
4fWhGv9lBpeF8mCPA72gQC2gXUTFpGibDCPqDGTLFYAfEZ0+r4/duQ5XwFSRBVWB
F5L0ftuaEBxELB566qOvoxt8scRChBJ9nEzx+Y2F2vJP7DhTjmIaKSbkUSQsDOzp
17V6/PrU1Zc+3pocTjGDlnL57R75Su9psDs/1PffmBZ5n/NFnlPYwNH/Cs6XiXuM
R5Lkqap5//aut8MMMHeXYQZB87xo+DIAJYz9pndoCO/j7YQNryjxA+8he4GL72xc
Le1d2fIGRV4LcbE9wlqgKzfJSwTgwM5A21+Ai1JUdBD9X6vr/GAeWLT/NeXrfewo
VXwuL5yRp4aviSk1BHmOExQUMtMt/JaE0dMYmdr77JS8J+B02mle7kPk98+1XxKl
NMtABpSbWFkjQroC0W6z19gkgHQVul/7zIBwsNjLaK2WKZ46oYtq2Ji6vuTlQ+zo
p5lwMcc23rjwn0C3+sE0BV1yxGutHlS9h5yM8IYWmycw03hGjWAJFLK8SQ/s2uzg
OsZsvM8nFDRBNHeANvYH7dTyDKx99rYEIYaXcm/4Vm+qg5IawCSNijkLGyO3CsPj
G8jWmiN05paVcCkV4oGePF9of/JykZP3Et7x8U9N/5uH5fFSx87wFiCdydPf+cZ0
8Ed4kEYK8wyhsufQCBEbEtCNWHJnmd+yOeeCThr4Jn3fCXmhT0MAhZNXLxLPY3PH
2g/FF+5WXGU4DFLe8MbKua+7QfuqNJtMtMq4dEGsy+BzsCBH/GVd2UQzndNBQ0wu
YLX8fHtqpvvLvsWDJBnYgpq3G9q/35VDddgA3orSj80p5MFM3abLQxDGrrckWcwj
ZHxt33bJj/cwiDq912sN42m3tSwsVvEYY8tNanB3RKPgM/4/sismFydrzQLJJbpx
gOca0+kcQF37son2sZ9jjSFzh9ib3Ht/MbCed/IZ0uYWB7dzQRVg0wI9YCAdhjO/
fkiPOshAkn9J71fJCm1u2MhGybm78KlR2xjSq/SZLMzfQi4uRRhHkPKEUyQvcaEy
vAULki6SYHz3A2zWpi4gm+cjxn4OZ+N9M7IH4r9+NN37lbZUV0CR5b8DURAkDuF0
MH8faNdE3q3onCMP1q0a5QgStf2Tx5GjnA2c+pZGUK2VEInOD6GQuuCqXnkVrgkl
ezVCuezYLa9tpJVJBxKnyrl+Y9FBOe6tAKBnsyOmnbNh8QP4074wJAbNP7Bgjzum
GFOwFng/3KbRqIMZ/Ao901RIa7PJGOF8KqQI2lumFQ870q1HDCfbQS62SsdqDblA
3ybJPP11AEHrpySjViUmXJlIal+1J1tm+H3f+N8NMzMi6idtyh7RSksSqxm8QxJO
2+sYSzgiLRI0bhssOLzigY4VX1DMjAS1qFDxUXsavzK6d2QHu+aA7zQ+aZDClZge
eE01nLwF/FdF4qBOhT3XOiYokSguQHL1gw/2u8k/E/AWTnuUv6JBlQbyxswuoERO
ZfRhhKUVy/oeZ9hhAED5+jg7Yl8+5iubfnuiIV/rNnMr0i7jBDDGWt0DlNRXX09h
K404GdT7xmO0NYYTfFZ2eVCQZszoKEeHWs2DE4CCHvWpMuCAon5JADC7ZGF/MJVt
OJE7XV8etrjgucmB+rM6w3js5O+j2DzecKkveFI5fYowVJeNA4a86kg3HnZpq9Qe
T7QbXkK0fc+5h2gxDnS7eGz9YViDZQVQQiMmBtH9EMFsnea4gBybJM8Irjwn6txg
Ti+7qp6EqqXUkT+xOND9TANS1X01ZV9woKhZw7gKZ0t0jrFl7xaHyzCOnzakjy8i
rWIWVoJzZyr5gthbuMGxOTpRrq+1/M+m0ic5iBGiDRRPslBWOHVUl3htmyhyzObz
/ztjcAdoAJR4UIED/2hfanmo6vjSi0Zsu6UGtGTOeYLs6QLtWgDpXQULwzeS+y2T
gJIa0tOxkhmvwQ3fsWr0UWt7881s1DfBneI8mnXwkmccYrxNlC3O0PQQbsULgFJL
GOT8oP0L3DpOFgucBaPfSUVqaFW2UPEuKLUP/SQkPCfYREIhzMUoANM5pqTPiTMe
dUtlklK+GQLX8ncKjUGLxTAHuvbeuYo7WyIfU7THpIKLj1dqWIVdxdwYN7NJTxLt
sOQFlMVWaeneoUnVoUM+IDEDlmDDOSieJkxfbr1+1sWYqSMtqGjP2oSjNgNFH4ve
wSluqsMZyxNP5u8sVQjODGvamxfH/HZwQBsTjxRAFvdEEYPVDBmgLJ3KBqS+Zat9
Gi4JaO7Xg86jjO4T9ozJp4/VU+po9IOZFWrRrRSEuShCclzh393zXkt95y8gNxdY
gVUVPMlKZmKiR5gCnVfV5hi3zAQkJJ5USSWSrf456oavSGGmd0bLBhGOZ/Wce8Xh
VXmCMfmmmZs6xZPz99lhZsXhwHjLw62OG1wk9/rmie3e+ZTLWfMB9S62XM14J0Wq
AneueS+i6J7lmuheCMdRAUcSap7j0YbJZOIqoLUJPbR1Me2vQ77889O5PjhtssRm
VmA87XaAUYAXmcOL7RUoL25/kWrcPgEQL9OLY5TsnMXD+YzxvcuJKd2bHaH0vYgi
a/Z09SzBTEH3tGdIOg452bAUTl+fKm67pT/FZ3NsbEjeO1TlOhPnHNP6tczyKnq9
2029KrwYcFyAOa/r39v3aJ0fL2USwiUtclIuU3y1lyLrGSsctJzS4VefV8aSSeGj
m9dt4KFjkDUZ/sN9k9G5C4rVf5OwkVKlmf8hyIoJVv7WbuTb9RlCJo/WqCaKEpXs
pg6hjzeg2xyfYT5pp8isVajp0BE/WpfSdhYuK5NZ1JylHsgTDf4KocR73wSCpaUH
UnsOTJVPhk5hSjYOsCsDHupsGNbHRk3/U774VXy+8hC3gmH3mwZQq8R/Ar5UWe7l
wO+lAzwYQ/9OXSN6XQLxFkViC7xYEhwO9lBByUsVtAVAVaoVRzM1hTa8LRn7GhAy
o2zTJ+yvHEXn/XbOLGizH1V58/IkLorcId5dSTiCFeXFCJKnHUYuslW5o3ziux3G
gcNgCfW5KpIqc36tevcnh+jKmR8H00ocsdPW8QJbbhuY0spMBjqztBV6MeUgS002
cBL82SngMNjerJ0WI1t1xQRx6NbjZ5WS3juc8k3hoXOhq6g6z3kDEjAWuPID4KUE
+TKlWnns1pfDRXGoyMznf2NfTeOUxHfoU0rVQI5sr1UNf+y/9qahXapkRbYVl+mx
vR9n7rhOv67pR+qPl5eVvoDHNnBCf1m+49f7hH5T0Ccz8bQwL8XOgQHRkE+81pf5
iRTm88dAiN5bOKkoXvIDtYBqYRXL/R7MLydcJ6MeKB2PLZwNwHkvouCzTQ6mHmlv
xZABV+eQQykp8Db//qrmt9EtmDzpS4DGxIgkn2IuaGzWwzfY/s+75pz7O1IHE5Aq
P3Lk3ssigo1+eMF+G/k7IBx6Yk+w1/SpyWJcIYhJFTkJO93B8soqBB1JBOn+paKU
RZg1upHfKl6KV/tUBOzHli3p/ycdR+N+7Z6tfeRrNnaizb075BRXoz63L4pP01ka
0ENknCji2B/EOzASXk352+tHUgt392AMlL55OqpStakLIT6lhoI2I4SDoufhWB2o
nVXZAolKEnDgbou8VkAzqgnV4YXER3yQWSTX1hWSFvJmPnJrtW4b16hgLttIc2x6
QCs7+H6vg7bNsAZDaj/Frzb7vrfLI6qf/lwRQsZ0XI2B0Wtv6dmJsGIDX9BIAXS+
N4g5N1s+bmRfyvK+pvVJb8g5WNNkgDrKPM2HHpJSJ6ex8oADN9oPYqe4tj5YyUsk
fKIR/GZcKjkxql1Q2Czz5LDNuj9DfaTJg+TWoxA7GOktfam0QK+dq9F9mbzdYuVs
qn6Yvzhfudpq9QB8h8pQR0dqODNYYPmZlaYRJrpVgORCytMOkr5+6J5NzCSc0DGW
GqtVIZ0XT8K7i392dHEZOJqKLgNTJ97iMZGCru7Rw+EXKQ/Bt99KAgEl7xKR7vz5
RY5WaiQnsEdB1CZG+wsXlbXmEfXXhSVIe7il6kyij+DF6FqhW3UBJ/vtDVgPeG77
whP3LE8DzdJQHylLgvLBRUZNQDYRIIAZ+g71YYgTMkfDMjEiEZXKEkU/mfw8OfPp
TAKtPIMGWodq6yakNUEyUrmQIEzWhTNm3GwTKs/54rLRFXC55daNfD7QHYrjIfz6
rr0Tjbr7GZjvvRKomJMHbaw3CfxBwgTNKM76gGh41yvn0Me8SOwWEGVPbqzJbjiu
6gcyIkUWZ+8DdH1IKZEW8vCHE+Bsxg7CZbN+lciP8kMR1zyue/BY0FjENyaGAxF9
vIN3ShUAZtulaR4g4jrQ8Y2nRABp/hztJAai5lMNd0gHF2rvW8tgBCpth4kGLMTD
Z0J6np8L8JyI9zwRYnPtd7HJw4+6H/qzdljfZqFET+tBDgZ/I//DYlYwkEvjmepo
qNlCvcbgjliySVpumvuEeDvUbVJpG/uEBRfkfcVqfszCI45JD0xVWV42G16ARSWi
xDJ+70fZZLFcPpj3u70qy6YF/2ywM3b26q05ww6jKK/0Sd5R62cQzZKUoef/uoNK
FsuKiY2c2XlU8DCLnSX3QZZefBeDLURkrgnPHtSImjdnwnfDvoLtQpVL4F1FllII
NrGUiPGpX6zBQn235YgqIMcmTSs4UJu7CPW+AWpcCjEl8FrwdiqG7GQlhtUteHdh
OfnDm3Ced6Fsar3/623fAW24S3aTzWHPUcVCW76G4q7lEaW+xFoDKykxv+rBgJxq
UeJ+aoAn9P6alJPkm7PQKxGtZs5GlX/+dcv/2L1+Y3v8J/nQtnHPV1hfrYMWSso3
y90jYo2f8Q6gOMcvytGPn1GwChkQnTZ6GLdXMknv8DkDjaXuE8m0ZU2/S+J7tV4t
3PQj3bs6AM2VywawOzRtPazwnTSsFSgYyZCdWdtXEjWEufnc+N06jq0G633+mZbN
14pvL4ok3IWZHbTyNmhnwghk1MHEx2Sg9T+UsjIY84vjKrwf+IHSQVNWSXx5sePq
hy4kHOVbXS9x4IDx0TSY1auS/oIi76waw8iOcEklSJepB3XiBOBzTZu12vdMNCvJ
fmMw6kDUwRrPHqOAhAbfZ4A8WtFHhkHj+d9FNdHcvgMs9Jmr4mdw9r9ZbZoiEGZ/
/ldLWYcea+6YHgO0C408YW8k5jKao206AbOPxKrRDXelfHVWM+Zpa6iQbC3ArZw7
bsCaXcs26k3Hb4b8nvH76paEtrtb5rSKavnOx2TpDrPKJpqE3o9gGLvtj8NhTwNb
j0vLdt7j9B2kVlYCLmxGoC/JiQcE8Yz5HR4Ofhu+XwyeKsKsrftaCqbnbViD0bHd
8nqOYflfuFxUSsYzon1CRxmv+eYRuuCLT+dAFvb0F/cD7q690YooWVBE5ZuUEmkI
uKmw/hWUjl7aYiq/aLUnIwq+NlIhis5c9NKn3YnrfEf3PjRTcKxqIfgjbLg0Cn6t
Zl9G3dtv0/MYwJG65n7xuMksCjHPkdSYlJIQMjRIlFaPfIL2h7edoQM/78Z6/ptO
KVn3Ga/ubDFuMjwydD0ESEa0A7JRQlEbgiV0nAxV0iVW7pcFa/TPbsuFExtIzZ6I
3KysO+rAgs5njfBnPtQ2wTsirEHEk9mucYo+JVQ8aNlMt2ap3OdwCGcvYYd68jJX
cD6FI4HsN9/IIvH9hmcfhXL+Y0Lmh+lP0Tm9WdYERLH/jfnaxhL29giqk0A4x6mg
WtyvQXgPIJQRLL3YtZNs7ifDqh98zz7akjjD7VLZUDj3bbeldiQB3Qz4gvwsJMvk
AWK/YziatXlyYgqWC27dx63ojSopFF0sjZF39howDVEQbymyvR/jTxEtT42gzD2X
uCUBtYnA2vUmo+hmIRKlq4GKlRsQnI66EyG5PExI0wwEaGYQiwxwDB8QNRID7Z/u
ePXJz8snrAlGUnSLRBKClkcFx85GRGzaasTeq82B0QHDXns0mEOqPxCdQo0Ji5pw
NHrDvtp3V5bcIttrbl0b/8D3bJ0E0FTzU+YnzMclEIeBx2HSfG6eZP7w9OB/DUzm
D97TTdZ8CL6dsdM4iyrQ4gkme1cejLMn5y8LzMiLoPcn7Em1YLCFP7qCBW3uvaq+
R0mRFOhR2OCzfSAwbOu3ydmkdxN2p0+ehzUwPaKDwX9dGOvvw10s3gQTGO+DswRM
btHlD6ZpaG/41dTGn7RaEZpPNLqWdo+CyDFUaErcu9Wa9gjj38zfMtSgw4VFZszK
/0go5+DVtidNETvh0HnadGiZPbKBn3nrqAg547vKJjuFrpiGrjHmSBGeupD2yAZw
S9Ei3Jt6ZEcYByjDGQP2VWXD6g3rq2bgSVLzQ6BoV821a1L/pCei30i5/hcuTu5b
f+1FKvMYxgn6zYzU0xUH0SKVHOfZMvObtFtFUU2KJX5wPJvWFD4gi5o5x7oMprkQ
hXU8ic+xnzDY7sulFKVHVwlt4B6Qy4UxRDSpRNaEzQ3WZk28CEZQsUbXAYZQyFvF
blz37fWDEXo61kwMbRtRQ53HrSAtbmMdk5NPtd9n6g/mOAu9KxOjlm33vz/i0sQy
T7O5gEOV9tdyhO97/iCsKXfiFrijW9ro1HsvHCfsc+ETWyKASDU/KO9rCY8PvElN
xJVkPA0hsuzuBP41VstZ2S3w5mA2wd/haXJ8ANy2aN4yC4PBZmeoDeRKpo6Au3U7
F8tE6PfKqwYYD8hHhfUbhLPlV1r1b2bwUXskt4p0syye2KBgsfLikeT0OjVAL3N+
four37eIbKUWmyqxPneWwB9cAlRDCioOf8FaFxLzTzOpMmv96HE458faX8ymgW6x
cbFpgoJc5RkizNLMg6KMJM8r0bzos3CacCc1i9/73TApKr+IUOMhR3HBcYPZbzvP
quQXvBDizNpAvJuMm/zW+Lwh3alDWIrMdpPOd58F8ZwU9j1lI7Sxrg8QWPbl3NSR
TjdwYxVBZeMp9VB3byKxve+Ks2ojWf3qSDvPu54N1ylwGSW+61zRviM+8F2ZMN69
3znG3UZHCKCJZxMRbEjA3RL8Z3MoFAfvOR7YkmedzdaMmLUE/FbydWQThKoAA6TN
3MCrhlzBdDgxmTuN2ddCUMdEKw5al3k0X13fU48VXMWnydvzqIy/rwWv1pqnEsQe
E28ho/+ab+tA2qKNlokOASoCD7jQqkSQyyRh3RcbRQAI4BrO35vcApnTyAbJTeAW
K0XZI8gBpXj/x+QLYMlHSBlvDNpCF7varo/XmWE4905VH/UTfVDSQfhr0lpeTK6S
DWyEL7zlSxRuCNveeTPT4SnfW//bQdTx4afO+zFe1350JHJ6cnWlXyF851xaE8R1
ugxoncmeDCYMwGsl9dmN8uMCQFVsFpfaFT9Gq01/jexo/M/x/tVXIKGSGfKsM78f
2+NqUkWds3zy7o/N2eKZOkGPTuImoywDW9sgluU66fKB1srVVhZr5v+Cz0emCYe7
cl3/jPLFFOTZK40Y7quL5cRSNVst1WTWknfT7NDqPb5wMlmJukkGSZwK9drYj75+
EwP001Z16fBQS6vyFKKoetqMZnd9MxxnZIZOOJ17+dj0zrivJTGmzF7LGFGd0tqX
RNMHsEOtQWOk6emaFzw5IiHAe8QiyOmd4mF1Iw9Mx2XvsaU+gESHKETn5tbbPU0s
+8U4m3kQtul5PC3F8OAwoGmSS0Y2FqkBDh6mNWWQ7W1WRAMqpGEksaPoun48MI5C
akLhxqVimAIuA2eVtiZUhsxxnUS5QUnHhCTTzFMha8aUn1HLtANtWKqmM5DPyGWe
CohzyV4EjZrUCY4XQUVy9NRxHz2X3o5Wt+/wMYxPRz7g+azfWPpv0kQ5Ady58xgh
W7B64Ay4t0R/X79H8of5ifj6Y6XTaHHXukvX7G4W8H75qvb7rxmzR0zgkFvg50VD
SjycNrL5+wYyFUypvxOtxTiLBIPb/PxFIVPzidd+H48laDZf1tq5r3YufPs0E5TP
j77g1mk+XcUknbzZRpOE7Rh9WBHcMv3ML8ZgS3l9KDoEWdtj3V6dmXLBarCd0/vK
KnEKzPqyMyY5fGO+59LNhyg9/SlQm5t8OmbRlinFS0sv49bGqxW6/5fRWJkv7y5U
zda7jXCJGdSgw2j7CgTIXIi7xuCgu11Wo6bPLdRlEfRHYdWZ0nnrxWrHcdEXkBe6
oRwxvHqR26yNpshQqUtxuQcxq3dtbB9nIPfKCTf9E8w3poOaz/9IWemXfFq34QSD
++NUDmhvFM9ElP6uh0jnmWJsRcXiX9tsySbSD6FbSXNrZ/BHE5upDaEJhgCsBiuu
k7bsyvaV5s2ISnujfqN75O1n3pI1buHfD21u5mltpOPtE3pyYDbqZXZZINpm2V93
SnBunapb7PlDVL4QLH503O5QzpAdKrhJjcEk7a8p/xcK3FP20CVx1cs1ghe/OMDJ
cPS5NLtQmZ/QzRyBn+0jJvaXMabPoqXBVF9O/zJJ5WRtVFQ+2K+Q7VcSi7wVXahA
wSTobZE6Xdq2fdL/EAXfO2ueEvuMJouNAZMn98x8SeYSjDbcam8zGkC/kV/mJ0jI
Pozf0EgEkpcGkNYwzp7vZ0tkIfROwB8aoJkMG+LQLXlMIVVz8EQd2jb0wNRBGK86
rSpt0EuNW+NF1vjrNIAGYGf4AMc8Ct8ye20LzPxx32RqslQ+8QEKcRKzMpbdeIAK
UAfx1rTPp0cXgObGFBQEPjabePzXvrJNIWI6lpV40WUf/CrLr6rC285TR/Zic3SQ
8Tpr1Vp9SpmDfQAJMFzEHSiaZzHhtweQITJzLX6A35KSHb+8kkkhOaEoSBPumg+B
sBoShpWDL/wmm8RLy9K9t4q2O+QAH4p5qHOYkBdgfjaWgEpjcVZex6991UySY6MK
ZCv45Pd1yoK+CIyExp8j0xffVUq/wynlzCqH/mc5vo9bfDY/LoLOMYA2tJZvPEY4
MO6AbHOPuvlHKJwV3FtVX3wrx70aSY4MW0Q6hQyUNXLWu8xnkMMWCoyn4sd3uHO2
UtWk1eW8uxxH4vKuoXJRIyE5JhdPo7tuX5nm7/eIlUNCVm8rEt6GVBNOUQ9O4yKV
EBPuw2Gfm12f26aBJB/5ZUoVyhVly5veyif0+qxGBAGRe5ZAE3UMHA48xen5HkNC
CWvC85NzlvpJ8g5t+Y3qmgVc4gNku4LFr1FCL1j2dbEw/k6GJOoj+g396UqxNkom
3KwNEqML851CwU7nyIAPEdAAE92AMRZmGamEPj+ptCGoSOxPMrxFi0E0OWcoqQkr
IT1xXbtHPTYchpmUi05MxiX6uKXPagQTCm4dQYBgi4LeCOhski7BRaH1T2Ez+TKp
QuzEPVi7VMjGxk7CLszCRfzLzsd/fmKsK35hy7RPDq5X85Wl0ylVrTsHTVAuYq4I
mmFjrH+xZTdnIRcDfrf4o1dYOcF7XrCo6wTO63KvPlkXygl96SXOf+RLsT9k1QaA
Du8pnHPsETKWpQZ1A0qV6zazvGek3NB/U1mhSsAiKOG6nQa6b7qptShn3alZujlw
13G1RiIYYjIK5vpA96BwGrwwK2lJjKXTPFLeQaS9mq06KCaA/J9fpte8G+HLbqz/
Dku0mvECbuge8rAVjnW89xe7SOEYr64RJD780U9OZjPxH/N1T1rerq+1nYh1u5b2
4hbTIX6i5K1Gkq5nj/Sq8KjST/qtmOmKQ33cMBoNjY6x1KvRUiJum/66KzY9GdO4
majQs9Mgr8qNVADTpymFFBUZUJ8D+hwsU0jtgLMOZG2zfH4BrLrsCmfFz0Wlc7Wm
SIqWCPESRsMDUq6GDzFwUS7bg2DujNdP4evkI8I5ib1jNpP3JYERr8cA2BuetItI
1KDJLcXlK7qRH659CI6RRCqvKoaTOI6utLV+qdJVVIc8nqou/vdMH6iD2gZPHLAQ
8TWX60B82AMsGBTwDRoVtGM8VriVMmIt6GBTXsgNto2Ij4q6RmPCMLEoy5qW0rsc
5xde4UW+tVTbV/T/+OTCdUtxgJPaqB8lG81pURRnpEQcXUlsFAJF9GWvNJd+fiFu
4l/Ux2hB0CtmTM35mIqQCJUy/oy4w+eAGczkmVTtZYE5wOOv7/z8AiwFPgC13d+P
0b/e8hiL7OaUmpdS0Ax23XYf2VTpK8SPqBTjiXpni4H5turI7XjWUG0Ai17t0qMP
oCx9m2181bhBlvKLrowvxfM/PA0slWDeGfDRP9C/zhprbF51Tf2cs9R+qbMKa9zl
3OtOOMOXDSJY+JqxUQYlQLo5EQyXYsCl7vys4/3uQWBYtTq7TJDix+zUovBCaCLr
x2Xf/A0Kivccl1ft4Mf4VcPZnw626HvTo4Gop0wPLsHSoR1f8PlsdfMiMg0dePcy
0lywXecixsSDdgX4xMMiryQ5Pnp3yWuM9zIcZ/o4z3ePNyFqOMDgcANV6pTHoJzT
n/x3Bt6OydT1D+aGUgjokzOknbI9yp2KeWNeZmOi4wAy6ngCVqfnsPyobitjfIw6
TUsOEAbWTqrBoPyvfKJhSeUxsVLVkIQrTO8NfchGxrdQv2URv1PvI5GZGCq+Ej4g
WyRF8MgpniuxY7qaAThlnRQj+Avibtvg//8ppypPWIe4gb7VmEHNxloAJhrHvi67
/kB9KGZtQpb50K7l+WO0ekUUexAXcAuRWik2zBLD7qzmAh79+Keu9eYHr8VaUUsc
av5NeqrztXhlcpZZiTRpw7rdVHTwyqNLYrAUgTh9k9BBNu4E65id+8etaoWzkBXa
uO6dVhUlEU1jqqdTfOQCdFsuA3TV7htPoHhWDvcHDNOSfKq6ZcSmBSj31+PrU7hE
r7ZzBYCluGeXAFx9EKThA6Upz3BzGaNnNuMpKIVp3DFY59GizbjOEHc7mzgTpYKw
E+WgkXBHRgCFiTfiIQ/zit9jhwBd+YSsETVaL4I2sXKNOia8MbS/5c7+/NL2+0ZK
Oms7SzFVkRs743H8xTO2RolpVoWUDNtsDZSkmVwueRIV2z6cFTI54SSIdF+QZ+fm
pGKYzmPi6PP7NhSzKMNpklgtvelxxX+ICClbqe04qVyV6z5UIFajJ4cZ90wpvByY
S4BeKcPJH2sp7M7NhzaPXo7XEZWVYiHf+nLniHJt37kNb7rcEPmjaX2XtxR1Fr75
xMUuG22m8nlj28HN69YNkNzWhJhMMpIdU0mCAVGiIBZFMQPKxqGxJE94d7CLwHp9
3iA7vrOhaCxFn/tJKxL8oPs9hd3/0Z6nTpqBftewShlYuwm+HG37G7DhngdOSC62
vn/x1DOpkeCzwQEe/89FqfDJzw9eQ7DjcLGYvBgGk2FnS5YcvMinUvnSP7UizulM
lwRK3OAlfKF3V3zc/T2jizYPQTgJSVLQ5QL7gLKLa04aNpVLWF1wjR86OgadrBXk
7vKJnjZEQqJbEv1On7HbVik0CK5wsEanIUXADPfZmy4XuClUfIOWg+xL5zrLc10O
TVx6HVE57UYFBgE6xEj35LOg2SJDRt7k5MIePoK7yZ7hwq/xBLUPECitayM45kvO
jBSa1/yjBZRtaS3ClJdd7Zp4bHBVllU1g3m1K8GskkDNzQbp0LTZ1RnCsn2HgX+U
zYqMUaeVNayuLlAhKTJmaa74A9Y5oT36Qt9Ai+KOpME3qKwmzeiZ2txKmWIm4C2M
hBjtdmAjDn9QbZ4s4w4jGohNZYaU8KkSJJ4EBduqAz63sB22gpKePzPhOagcJpCy
2rizo1nroDacIv861rpRVjrNZQ6kGCeKUO+KRSIDi56t7HpzjBLodEwvA9IQMYe7
aLAjf51V0MxFgRPda5VGTLU+qCD0sp6aZ3yFNjoIa4Jl4EvIeDjtxUma6olhT0+F
zNWzpudlwG0jE7EcFGhhyOQfDxnygybnQraBxwM0lWo3uKmnbS70AtsxJYQcQaAf
ybjLanRBvDzz0yKxt23lE8bVmpxQ6wKrn/AFAgwK8rs5+jRthIxCch5goJ3ceD/4
S9RXYPUZEinRZHvVvNsE6eiLDSn8F6NKgQtQ8qHNDfmdoac086xqRQU/jT+VtLky
keB/Q7JE7tNWdb9TcZq56vfukaXp5oBlS/i0/+VCzZnYYqgP15FsTpH42JPzxDfJ
lFIFkCbTTQz3z59SgCGIDYFCnHFeqBbkR+Bm3IP8WLsJ3Qa9II/nSDcpmDbFkd6B
1hJyUGPoH0tRSGPOiTDErGpjcbY+5abC1+P1Wl9bsMGjaGpmUHxZ8IFQf4bd1sSu
GqWyDGsm1ytb2U/H5rYdXDEh0RYusM8EjJfUb0P1hpn/+Orp8Vttbj+P8SxzJ+0Y
ybv1nltF4XMEzZYLoog6m0mc6lJgzcJhOpB6KhYDB7lIU4wp8eESCEnBfVsTfiOq
rlyaNxp1j5Ojq+GjPBJv6aVH8OMaLWtV7CKim+QaoGFL0sNKZLnf2vYG9OvOm2qq
SRr1ZApecVBteDa+hqfqbDPJ6+B61XF/EJCTVuznPpH4SzrGiYvN1uCtjubkC6Ql
MC2QPKPnq4F+r9JjfgZOFIQmKsCgfHXbdRExNk72Z7KrzxTB+noq7Pl/go/gZ8nN
cNbcuKZNCctmop8jR5Hf6uHLgGABjuyX+uRi2AeO5LDUQBO8W5xVjl2d6WWcC4Hv
JKeiAtZwPAaHQni3ffsJcKa3LGeicu9336trV9WGkrgmUhEUKbNudfEIQkxxSma/
0HbWYRiRmKCjvTnby4dhR4mNK+rjKDrTkcFbDlHzeexST2I70c8/gibtiOXCJtzI
d2NJ/P/QlU9J0QXkfmytgnhZ4T/Ogl+8e+3SIZWrdRER8e90p4Y3XDE5hnMKFKnu
8U0EczXuLvc0243kBSezCKVPrBeWXznnIkMH0o0nklDOuo8CCOjqEffI7L3j8RVl
QfanGmHyuLDjrlkGsFTgoL/puxG72T5yKP23DJkbJbv1ldZ1Tkodv5oUpjAmgRqJ
EkPPvY2Dn26HvcdgXZpe+p8ClGlh3P5po1JcUUZ9+qsuQjKDvafSk79fXEGCmRT9
zXqQaQ3s7rnSTJo6K2rgnBwRwXkt89R5PzrB3MqYrGiQG8higFQK5NJkSi9h3FBO
EMa0N4UP70PK1nqH/djRkomcxhqQPozLCRBsrys2RiuAv6uOMo1VREfUBrKdjtdM
P8IztZgS9IsAQLgp2ZhFbd/L3jLK7bfwU7U0Hq0axABeF0xvtYUDQQSLSYOVbXtE
Ng70XxTO3x5KrPAryurDoVKG0NjrWTYkxx6cjUD6UhACRDsucCaVxoC7jdU/VoA0
yEia+w2Y4Fpo1url1NWxxOXiRfPFBqPWOFeHoj3hitM3tNCpT3fNezMv8c0NkFFi
I6C4/b2lyAaj6iW2Gxws1D0UfxGeZe9fktasNyFUVZ+2cgD/N6DxqOm49aaGBMyb
Ao1wCh+DAGjL/bvV8t1pERVBHFOrQyGT4B6RVIRqamURWzCGE280N/QG1dODZV8d
H9VMC9ULYu8L2mqU+FwU7mPW4l+l9AiaNFVg18Mk6GRZxz4LOFysj3M/9HrqkARg
gn+Ktb3AQOhnVBv0Ni0D2OmXqXAsQWrxsyfF9P8zA0qsl+lxabI3DlfYIbAtvpT9
UfO4MXFsEMtF4tc14cPZL2Z1fUtzKUXhwg43M7bMtgMZxwjpzPc7deu5ORBj2jIq
C0q2GpH8ix9PcF4sq6J44L6CCtqVxT3afNx3kYvsYaDDTer3YBaLxSAKmAcT7qsR
SGrSyCYBZKyzE5eZSyh1EyBWBhYmPLFbYAqq8xm+UKg6zy+UvmStvZQUvOGzt1Jk
IkExqPb3LHvarFAhYT84XGUYudpVCvEqA+PVE/auiSkgxRKYJTfV7il5gmVLJX89
gvYHFuDQtuuPLiPKLY3h8diNMu2V5ocVV9naZVabCsXuoQYGOKTJmcRF2/LDgS7E
+qYeprsHsX3dT85fHBW7dMCEpAIZ85IgHT0o/BC35m5mi2n8Nlbn/Hrf1fpwtaCW
fB30qeeRkvau+VBzXsXofn9oxlNsTCIIrMkP0X12onFUA8Zh0rophyloT1B7ItJX
vDK3EhXzy9PBq/+DAo4EYm3u5I3Q8uJZ5ruPRnbnVJaOKzhKCQuYhlXAdFuCGgSq
LAFwLYAX91FkLA+5/ZKEdYFnqMdb6yaz98jB9UtSnoFNfbRrcnOTHMfPsKOcoKq1
sSlf4cAvFEA9R0Yhhhj+R1Y0UCrQZYb199A0DG/JJBlo8nH3Eo2GFM/jnIGqd/yR
uaRKMBdck9Z/SWAN1Aslr0wqd5PSQiA8rrXMPHpUqE6FoEQL6taBuIStPNTSG1yv
DiH/wHi4AxC9A/r1+LdOyyTyO2dbX1enl8hT1HCj8B8tCuWYukWoRbBr6TP0BiQs
Vv9WCpyaFA+tMDuBlWIy/gVofuHT4kFYWQdGTv+MqKmQPYLdwMG8FXPOzIpVjrC8
PjDyicDv6reiYPEuIvLuH4xoUYNSrbO+evwLYGBYEs86w/Szgb8AJm/eImmjhrWu
WS9eCSy4WUmGR4o+KN1yIosO7YtfbRrzZq46mbrEspj7oVFj05ZqDjp4nbr3BABs
EmqpI2bMjlSPL/NxWYzT+9X2HxFVhORuoxvOEQ1aAgOk6P/RGOzCZf/7BNDcnIBQ
2PfXd6ZuYKrPVF0+I7iqbwn0RBnsQ7PRL5witakJCew0iR8tww/LCaNVQK5mVrGi
pXvB6r9EFoJgMn7d8ehKvZ1QxJ49jhc60M+Jvcb9YQ76SyyvmKbUEQzfLk/dpZwt
WLDOUj0Bqq9BoBbr2RRH7kS1dqzMwV2GlJzK7JXwx/J4Cx+hcKWH+hezumPsriNk
wJIMKtGy1ictrpy5iR2NT2JTjpVhxHmciLKubigvdX2sbNbdAbuDEFJvgvYhRDGZ
HbBigugg3JdqBxbc4AJNOeeVh/yz7N8oHb2YOx/jjpBSqxyu9eNNTxzy8HpbGHaV
f0DK1Vu0WLjqhaNo5WtGn0LmN3v50DrRURlzGPSMkaAdqmEuJIEwYJCuarPprJGw
tB2LDjbtHvOerrHm0LBjvtjWHgYUW7eZKDmukqfhkSw39jZZM/YTzV0cEX0o84Yz
XuVbtMpLLkyfGRMSlVT0hHvMkAB+4mpod8T7xQZ+ztpOtWW13A3nmjL5Y+3zYqg7
Jzk6mtt+2TTQacfEktXmbnfehfeDGo647sQ2LyiY1mjuW9TaDkSYmWqFZPPgEr15
aKCbPXCnrIzA4b4Ai2MKSdgVXh8NzR6uZ1D5HXXNy/L/O+MKBosJItG8uRMEd2Rh
v7tdanb8La2aNjBlG37qeKMsGqLRjh35C/0bHFohb7hVRIR9vnFQma4lAHdPrCXx
Reuga9x5vo1NZJnw3MHFTZs2XyjswGDxLtOFCIjydZhyGzCbDGpnTR8UHezbBIiS
kI7+ryFhd4Fz0dhGNqSp+oRMCSK63w7yaC+jh9v0WbYgxBs/3pTWqNR7IvRBYC1m
y9mmsrXrJe7sCcDBYnhDfIylr7xT8+1uua4xKT28J9dzO8se/6I798AERbSTzP2S
oWExsYtOMoJ0I0UayApLFNYd3tx/UqONgcm7OVtVM3OTOB2v1weqmSAKGIDHpUPQ
r/jPvbwI9Lks3hVdX8TP7oWbJyKWXsnsUmm0jNR3RAGD8cIWLsAsljGyNZjaAMFC
PqzH4MsZ/gYU24y/pgeirs5D0FyzvATZqynwcefsdDPVM1mzzU7+rQWj0HgPkk9P
zhgfSQMV8rJh3fh/OgSOP0yldVIEz1LDmU0z57MtlIsdb1tZiCLQ1QyNXJFWNsSx
iL0k86OYA90V61P+WLn7tl6B+rci4WS6OvGVTD1nl+JkZ0PWSdMkZFqgQ2D5jfBQ
rokqOgFPHbjCmptw4O+fUzeCA8+m/aLUUsLvg5hvAw2A7woL9pd6HEl3pK5zYAJB
oH0t2pZOWsJ+3OE8oovu33PM0dtcSgEV+RUU+RkhxLhouKyV8PlIcrr9I9AKR7dR
IqvCSUmlGL8KmMzWZ1msMmhTBH/Le/u8cv5U0yjawaMb+oFj1gYzNDjTepkc4Idb
SDLYVvU8zwrTo5pTiso588uyIvHHbJvh0T70w5xmbbsmQGkL0FvbBvYlK4ZgS5G6
GNGd/AhdKNu8ZFIbNR0TuuqxVx4EcrvLx2qhxPkgxr/E6MMv582v3jCGcHz8IEhU
l4hxnFDZTmXdxnmd8XgNzVlzCmDJvetffXSPjPQ3q2+m9wWjC0c9/iQoyGoZ2nYB
+QPFRHf0dTEQ+RnwPjmPkPmaLzkk/9xg0TPTMqKykUUSXa8oWbe6ezcGkANou6+J
iAwfhe5oROpPUD3+u0Xp65UJCEA9ysNFEUNo8mqI/BDROnsiVSaJ69vguWYgg3da
qauWx3urKWL3mcmaBhBLVFSFWasmv97lf9hs+UjpGxR0PTW7S9dr/p5Idmq3Upgg
uOShMQaneOlDXe+OSmdD2KCeTV04u7YWFJtr4MOqHcBXys8WtSDE2pN3l5uXRJ1f
8uk7r+NFD7buga8SE7lqyJdcrmbrvVfKmygM0JqHhYDdeFKHyKkfPwUS0EtgEKWY
3uDOK88kgVlrXaxEF0I+ijnHesF8vrTKBjaYyK8CXJ7OrrrtTL93AY1hUEfjQuq9
lEhMV+3ynEqqzHD8r4RSCC7K0ZLYM/fZuqWudEM9tneXfjpv1WsNFlusDpCVx7Ux
1H/RzaI8whKc9Ak8xqUMheBQ4336kFTwvo/DX7BdiND97WhoUGUWPJMig4AZBIfv
oXWql+YtzRRJ9ZhYl5gN56lInx7BU7NI8fRp3qckJGwjfTyGKNTcbYfJD8e986Q1
c+Q9WHqzcAhyTyKq/uJdHcDAHVhXxjprah0W/X68PdoeYtujn0lnxf63VPuyruKG
uqyjb/kkPVI5NYaZZDQZvUOqtAGH8IZpAl5kttdnIFa7iesXosPef78BDBOR/qVk
7lygD0ESoO3mi81vYbXN7CZ3V+ROYKNLy+gf1b4bXroy3INbG8sLWQ1qYtu3YVkx
HF/NzcdiJrLWFOV4onVLrR+guZtVJj+OI040/BErkO6rkgWfTTpzMpQAwi9MdteP
PwegbGZli/+jGsaXZFuQUC7uYSqBJUNBDzXj4J0oo9aBz6O3EwAnoUOTIvn8vzW/
6rM5uST8wSxFCL1rBOSi5F3GH3i7mcxBDXWG1jh1FSoHnqghvGt7KkY0vwa9SdAp
ZefoEEDUKSJeUtmB0TMsPNknXXUnhAse9L3n4iHlIaZhO6IzwktXNUGWhX1Lkygc
0qpucGHFZiZRTST4EhI2zIZSb6HYSPnlKUnzJ+nW3rCT3Gl/EKp2EhpnM9b+m+N2
lO9PS2MyH5Oq+4jby6aK1RkC+lO0XPFpi49lvFbVTGePi5xfhdnVBYzLpAGZ10Uc
/QCCL1r9A2yMiDRcv5W9pT5+qJFyTmhMbzH741LSAn3JNSde1qDCBOaCtuHo9Rnz
omnZQY1T+dyZmxChxfOojqZUiWbtx6wjYO0Fc+vnmYAnO1Fe/EYo/Z0Lv2A2bPd7
oqawlU6fXk4MZYH1+vuX7O0PyvRY4KmNtdRF047ABJar4tLwxNZ/eSoONpNFlzgW
e4VxCfjzRRYqICBeq66Lsumdc9RIVh789w1xn+uVHuh2Yov8vvbfvbi242IhCtNM
CvyIyXQpflnQMDX57bjp8HLsYz8GH8SEPBRej8IY9BZ95i1O4C0d+/KWwz4keILq
f/dhmmoPbuv4D4ka9btxWT6PsSb8jLHXSPrUX/sLyW9cgcGSB8rT9VV6TYcXniUr
HELe+jzS/mlDe3KlVurg+YEvx1aEP6KWbwpc8CNhWlU+6gcs0HTocUOjkVMUPYT7
eDuyNpLeBHxURz1stb2Ott2bteYwum0VZZqVAPD1qBPCESCeMyAbBP4Zvd52BLGC
ruhhLk70sLOz+vPXcjwJdH2pbfd/J4q0jPkSLZaI5nzjRQWljVzIxPz7vxddzFyE
RIjIs9wOjKtwPj9x06WKh6ibTOY7Vh+nJA0jbSEOMGamGpeoBzbLMkvv7QNs4wk+
VkVY7Jh/5lskSdKUi7L7BjUAkP7HEZepLPey5BsYyHR6/TBL9h+coPfEv2Dy6/3N
jEkILLRzCG2QDa4ZPVj5csM+pB5EXfzGe3DiFREdrLMyIbLoP0qRa1RMn9v3RtuQ
/62+fLFUbYryRisZfmbHa9I7zdt2KjtElCP9SWFaPNNrfVGaQ5Cv09KWddronQpv
Mfh0qrPy/LViF44QJ4YY4BDG9K15nE/V0F8BWPMJ3IPb/P+8hsdh5oienVP6oPzW
JJ9InV6CcWXHuijucoeRmNKBUF3zZZdbaYdXhwMhbbx5MVREuTqa2/ot+2U9/V8C
CW/zQt16R4lQUgQGxuIxeraz/rJv7X3j1YIuXkqNIYu8DiNAz25g0cqZUjaxEsI8
oB6m19JM+aBHohzFl/SFAqEuFkD1c/lptAjEBBje1fQccqdvhF4yBjox0/4K/5G4
p1MPh9fhayjY1N8C3Gm0hFuELA+5CvNtTg0upD5NKLX51Oz328lcNc1bsT3tkYld
WGGxetP/yohGgHwF1HmRlCKmMxZ2mDfccB5VV06+cGy/K3dD/UInW09ztjkbvFbR
`pragma protect end_protected
