// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V0jS8P4VZnkjQrXmcwR5VHFpC1iyXuRrkzy/CxSQS0W6Sb4ns7nSKZxXSRqM8Xl/
0B4GjbbYk3B+qjXXsqBkVpOHuJr5f3fbrjDx9zQ3OKM0FtfXfwIMBNcCGLEtR5lb
9N/juSmx+DgPrrkW0fpv2JbKmwnlgs2KLeEYOa43Nb0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21680)
upoNYZvcGo3MedeJW8BRuvze4nYVjn+Mg8wB3ED1/1NCkNpFm6zDilpMZsIRFjaN
zjMHn9XY7hf3e1jqxjKFY1VL9JiCKN7z+Tvs2uV80rhsYZYfAZ0QxPKhIsIbDyZe
bG4rHefFKruYxIT90h9rvSv3isKPduRqeISMUo7rItbUxlQtjtTs2iYeEegbKluD
quqnSr7XfrXAlepFdYTS9lLuIrhDf0CAhl9fnZNMf/bMnRJzrG3P6u63o690KykI
FNp0VqrlNjSoJdqWJ0k8f3yR8YjNIGSEiWxRNqgAViJPe2AFbozTX54vSJ99QRX4
7Odeh5sIU9gGcx7ZXlPk7/XBBmh++iy78Tt5sBcoxC81sgVk0nyqWhH0iRTMu748
3YN/c8SNifmqTfyoH3F6S3ndGWcxgHrufoAFeWFv4M7u0SZDOQ9BEDsCvvKZu0ft
5Y89ZK2o1C6lYwOPvjZz6tE0kmX15sPOX4qdMv1cDBjEPAmQ7htU88//5UiKfs2+
AvKZ0U4B8ewd/XW4ugEYCWK80jXUoW0U+xLdbodySCq0zo7591x0zNAMmepumK03
2oqM12024jXNwLe8v3QRKfBRDCoIAfW8rSkUfJ4hyz7L9Hm/Kh9I7S+1ZRzCfE0y
vHQAmi9xQzDPsgRJSUZjgvtaHN3vGp8q7uwt5ZgJZAWqsUYRjd9dB/6mPOAxfIK+
t0GaMugFgi93d9WMu8j30DglRg8IW/Tht32EXkgYfIpNf+WQsn26j6Rg/Whtk+cq
deTnxYrX1IM+Yj7H4u0iQ+quHxeKKnXXqpKScJcsWvw5Mwu/4c4DO5fqpf4nLqBT
Zfvg9uQYGYSJ8j7MgV3+FAyte2rnXKfG43zcT7qwtfo42nvb/cTULL4IejLdgJn7
RPs+l7sr3vm+hxG4C0WKaf4KRXr3NWlbZzABKJ2GEafoDf+nU+uXwK6LH0VI0rfi
ACLD5YpCzqBDHRuB+m+B58hfjnfFBGQ/Ais/KSBrSdtYZbNo+qbfeBshfrncbBXp
U6mB4qhQDZ7AO3OLQ86jmkb+jH33OgAMc8V8q1N0MvXGphrwv/FU+5yxBHmuu46v
gN/c4/lkPbA+Ds64b9tfTOtXIjw/2Mko27Se8dAKQ3puBdQ2CtPLBWmyP6jHRJKA
p9zoJY18z9lVA1gKOVKEIbniBBFg1khvfYfA22AsdkRC7G/JawIw+9uBrjQPN5ds
ESXDfqbuiPIkrEy0V8BW/iDuLl2tMLYReah9StzToCSlr/jBilnW4/DChH9VCGFI
mPGIlZxbKXoYoEBxTZCjl8+wkKSTLZ9h4J84kSffgVzvNoBrEbg4uZ4nUgxbrfda
0F91jiIWbMrpZzj9kogVtqTNbDx/UoIupdvkqOP9Br8Y/jPXN4obxxFADe4AJtVb
O8VBBDdJs36hUrBJ6itFBWlQdjLpBQHTlVwXC0Zr4g+JuKdMysbHhrKizh7SgP88
QrbK2l5f1zCk2SIMEvVBIGjykP9PIpgQk2pY0QdSiQL/ZSY/gnyOTBqBR+ym5uFb
oXr//L3CD0bZaw8Sk4rPvVP7JF0fyeQgiTsMmqUFtqXJj1FyVBAbRE9KAVHQ77f3
y0+1Q3PG8m7owXpBKzgCfJg3Dqpn1yWkQCBdKHiuB/MNsN2PHOfGWKpR2M972x+w
aFVZD7GO9apTrjMwF+oqcM/xOonLm6GcI6El5pYDLG3apJqgxXpEBTxjVXMtEAbQ
AWmaEzi6Ok4bEicpkOSIPTIDw3QgjVlkgxAFgSxDQBiwrDRW6kNqZyMe6WztvUlz
TgSuCBGhdYgcPuwbFSoTegbV82wm/lovKLUacK0f836TG/OPXBMfAtLmAGK6pv50
IZYPKWt60eyFKr6h3VdTcNQvccxbgqD0USPQSsdPKp4rwkggyvSfxPmbIH5wEWEL
byLaYpHigXpW2MVIEQD3tULuzGS1qccX6BCJ9xEpfSP7VD4iemy8QPohW0Sw2ir2
yu1rCwvQJuqQQCqMop+a3WHZVzhc+NRK/UkMh+up0UMmEDSAEHGBltm3s8o2JhOI
P64XSfX9edTU4Dpb1mcJn0UD7S34BlqlMugjL13Bt2VNGJSlHe6b3TWjze8l8OmU
Ru2jtY2ZiBdhKijsRynfAGvqbuiCTfCI6oGQBZCxid3Tlfh9QLhb60XIMQheD/kX
u+OAmRpFsku6FheTQGI9CjEbwgIa7acoDF8yAwfwblFbPIN7AM9JNINhKT9aGJlJ
VyCYpDapRfCTJhnuZXUciL/Tj1dpaxZ2oizkhgq/VjsD5kpwbnZ35gjIXSxYma+Q
MRU2qEUSEkf8602OmRCxcU4CT3PbyUKAgSAfA9+FapHM0ab32w2YgUebPVwDIaDq
+/qyk3hf/A9bbXWkrIukF53Yz/qJ9yS2Ah+hC9bkoJXWRb7mWdZ3bcuLRMj9tpjO
ZbR8wAGNef4ITOGcEcGpceHgsfm58qQyFYfn9Vij7+dR9Un/6uynM6BVToznxlRM
cuCe7pmGt4XSnmlmmHyIlqdmV/7DWj2jr067NlhHiPPIYbHKOQ2rpEM/OTapic45
GfBZcKOwPiAgwDwW0q7tuAAWYYm1bINt3mNlbLBh4SeDbtbS7qjsh4OlK/U4+tXW
Rpm5pytErroGxgHQ4pWTMYZqbEwEqAYUCLnCuQW9oO8VN3eqR53E+wVc1m/y5GV8
L0xL4DPJk5Z6GqA995vS7zMpfiVuWL8QZzRqsoJ4ThpHZGeR20N+BSfD3ly0Uw+/
yXP/gK2Y9UibGGPDgxPxmzSOBppJ3PEyAihiv/kLInBvCROl3hbmLmk7Y3XhmdIY
vGPa0jGXIvISpyPxtauunjBijPlrXZBO6PEfsE8bJzTmJ4/OD0YBKiOlA4BFUbhl
bN9ASD8uZLtusVDMzhqe27DHQF4RcAdgLcbTXag+STgsARD/XHrgU0nWxN77KouR
pFWDvT4aOU85PWPUGFck1DBfbRA6DGiU/DgNEiXLlqo6+U3VgTpiU16vqk1DKEy1
xEDKDzVq++xaEIBVIZByieJOvo8ajagTO9PnuL0L9lJYUWu7kjomjvJDyH9euiqj
STIjPZLM//QNwLV3prx90uT/ymZPR9cmo5S8WZDITW18+Y7xXISpv2KdTrV3kP19
+w/pJpFhMjgWhBEnFQRcGcBa7fIEV6V147yOEYScU0Uj1XTsI03IUsuw1bEWP3zL
61N972Vzn96CRwW2LDtABlRW+fDLlN65v5jxRTvTPpKmu8lBBVo4H98CkqlGRLbg
VT2xi0ZZXz0/fLv5P7/Urx68S1Err0mtQFngvPnxP02KMzfPgUovBTdgD3WnqfJf
6nynUtb/ea/pCYowRlZMSUwkZsfeyanDw6VU+PzKTZTSUInjrKBOupT3EMBR0jms
TX7Jnzsa0WuhMQL5Y3cZ6owck1OKQN5i8neNRx9V0mAN+EECTgD1bkKEILVgXXYJ
HmIjwKAlPgvIZSJA7bi/WbD2QIA1CiPLrSOnsu0nMxEFvI+qFXZywOr1E1mWJRw1
RO1wMsOyl4CP804YkcYzDb0UyXcO31AkhUuvthOdiu7q/IzuojqNhl5WafePXN1n
6+IfvXrpmXLCdzzN52/W8DQDgWTrZxj9wSRha7AKqXvV1ppEthDEQIQnEC5j2RTK
fiz6kwk853uw9X92adZ/MqOhxn89qvCivHdfxHYuzmG4QbtkWHmrAfYYu3KmX/UE
mlzXaT1YpUOyaGiO/l0KHSYeBqsVX47C/Nk1PJv2nQgXU2BoJhzm4gz5hLjRMF1m
+BlCUJIcNyiMAlrou5DG7lH0X6Em8MCho5C/pKMkjft4BMgL5uEMsvdqghg2DG1z
US5tDtZQvzx2fqpMLBMrFrjy80vKqGJY3scqgRdWdx+YA4KCQjIaEXMsYWcEPPrV
q3Uqz8vhltXD0lgrhKSRL3CztOJsJMKeEjxX9RzP0hqU4ERAidPwph+d09hwpzXA
0JTJLhK/gEAo1y7DKM/+nZjxe+jbycCHJ6iID0JuD4l44DfMcjrNT06HMImsw/In
fw2ihji5PZo8uhPh37gyCQQI09H/D+0f6Ey8/dxf7qSvDPnW6McGAP538cxHwjmX
JW939mWV1Og+60DKvfx5bVVGzJid36KJAXnOAUZmYgEpEPewwM28ExhaQY5Vw8+y
IDlone0aGhe16uhZ6IkhDML324xSFyt82oDtFgTl1gdjmFvFBT3rxBlDDklhOwgJ
wYsQr+IucWr0JP/PURF3l1+YL8jJEkh3seh+pLR+igg5zrKnTmeqZq5dhog0y7Ft
iVYL2z7aXP2jq6CnbTLLE4VIkSHCba9tcjJsPSEVervdq7QCt22KkweFzcnWQKw3
eDbTLDL+weZKGYj9Of9pLqDxxlPJ5jM3k9mhxdaLv/ggfb63EeuyE9Q6ffDgpJFJ
mTItn/7+s9+u6ZGJDeUwI7JmKA68SqPL68hczkI+9ZC37H700DVCy02sUuw62ygL
XpPnDzRcd+ouPKW05dfsKWViRS3KMd9ADelmGs/lOrAP7zTs4Cq0nV3LHifoqZ0h
CO/y+afIpHYF9z2oQRcWmv55j4vGxoxeR+j0NX7GWLOPTHf2zowYTf557qF4nPhO
RR+jjlruuqjkeQgrUvoBSsxRg5FPOQS8CQN7QvpLBnbKs9CJGtrEEPaX1KmeoTaO
KEkna0soYRjAalK9u5lVmoxKNevC0PNQKfvG6Xk0IJPoPYJ4QLbykOmEtKOkANtE
5NHBC7AccljlTeZsJRVUlDBVpLwC5j3mZiLoBpgtG47xkLuH2R0Zgn5PeQ4v4CVW
imh3I1O+t4sUMl+GA9QwCQMuBisp7B6JonsAWj0YzGHW0bZNUtaQLxTsgeT1I6IV
4qasxad1dtNvvycEs6Mz9MslIqNKwTB2xvf/lx05rNNNg7bpzKHFQ+Yvls1gASJQ
fQ2Eg5L+WjiHyZpwtNSaE9rORC9s0gqBwAonY2hBewBgaGnK2M8XYIzdjtKcTCav
a9HP1H+UiPEaYEZX5h2fw9AIYWfeqJTu43l1I+87Y8aTYPKuM5wNZiGlVwzDJPHU
Xoe1Qt7E15plQPL6GpANMreeuLoLr0qSlt/B3r8RJOKiFwJM9rEYF5vgCVCldzAN
1QGZeIxKseModgjCXEUcjqwSQeKSHgRTTb6yDteV5HF3VQ7a7UXKnx5qqA53QTCo
GB2cK1+FjJqR+i4ix5ElRIrBCaBoB9r8cTSZkfHlJmk7dJkbSot9zWEY5jr5M0DJ
cWJgFD3B07HgYtxUyI/FoaKO/VuHrIDYb+LcXAomHlQGz8JKHblfm9IaLneWDIFj
8Dgz5+wHSrZfsMzTniL0k5DrSPNCydwiPS+mzqCE89fHE/+8ILeaawvOKSTQ/+dz
o4RDGJ6L4DKai3m8fLMX+DrYr5qglwcQ5WfnBD31lmIFCUJJqcX/O/V4j2ufstJ3
xDlKfjbdZUL4t8ljU01xJf9n4roQ1wkIeuFdJTqmvezDIY3xel+WZTmLreY6cmyW
DXswySnZfUZViFDNOYZzjjNzzlTZVzo5SXAMMsRlTJoPLmC9jQV+TLOOaF1mh4ky
b10w6jKw55Vtg7epdTDWhgd60t7NGo/QzJ/U/FhRn1o5KpjPWK1gyPY4NQl9xXd8
iMDFpnJNFb8nIkftkeRSLB6ddMaVi5FdfnNLnmCh4gNHZiNsmP2EcL5h8Hn/ZlmC
1xzltln7RHBR1GdalQnNHFvnxCpd241Hnmg4pjKDlLPOevNiGKsNmu51p13C5tkE
/tbbnoBj2jnPVr1WDxMsAbZLx3vIZIuLDNv0X5aJwdBa/L+csWPMmBjOHqvg8bNH
jpfdcBM9QdcNMw30rC3xqJQ27yYGXCZcqvPUjmacgucEQo+qT9WxR61em6wfn+0U
vlDEdjRIVLutiAjEnWqt6uXtRvS7r/w6EEKgAN/7/nbdCJPNo8Zk9TZtggRy313g
7ZPM3+NN4PPRRk5TTN46Z1wQPVe2dnRfIodW4+/Cgc7hEMYt6i3QLv6TsB/pWbeO
Kd0fQRIrLYXrVk3JoQm88Bcy+7yfaD5eime5S+OAnLEno4vT+71RdlJjJbi07oEe
ZpkiuKSfW+V2wM8vhAaKDEffHZ8msC7aEQGDRwMg+Y1TYl3Pixque7J3sbklx9N6
Juwf8x8UlD1PuUpAbPFwzkPGM5Fq4IaZESrdyUeFnYVq/EvH0fT1mx5M2zt/ZMup
4zlrO0cOKoNOljSNsyPwzLJiJJ3yoEAnzXp/FNOE8hCrSYobm6wkN/H2iQ+fX1bA
aOUDfv3i2yZD17BC1CSn9H5z+3YFsx2xOV4xMGvWMi/q0Ow82xDPaNjPGEF9bbeD
Cg0SX/IovkeE9qSt2ERjVPqZ85uQGIdK8qEd/SeeYaCQCsXPv6cyyTQhSfj1g7Am
e+EvQZxpVrMCxR+nVTk59Lo2miQqjAtXqPQa2lcTevsBEooWWzngflPimAuQd6am
KIs2k42hy4lh6H04xLpC08AfiaOABcv4r48Z5rFYYorGSmHGnXSd1Kh1fOG1CJW2
N3ZBllossA8A6sb2S8AqY0lwOX19T3AHKxkyFiiqAGM+bPZa6MhsgprNmLO7sop+
iW9jjICO7Drs5Idj4jTWj7NYkHVapVW4avEnWOSp0nzHs68lFKq8wRt01C5IIfti
91DUwoKQeGMHs6+lpakCjoIy+QyqdQyGXSHhiQGHYMGGqXUKStcxwe4hcCNxx7ZC
mJmkgNolwt4MDAPMuNYbo+/KKXe3uMQn6zdmHBuFhPId6wDd933OAUzQyfL4Mhpd
8O+BEuAKb39pRrTuSSwKTVko78Bh8URnua7qX+X+5CkDZtEvHY38vOa9Q3c0CJjK
AiEcZItHwx8py0z8HHHlQapvW+zmKDJ/dpOE7+frDAVwTd4+56wZ3mraVXCEQzwg
1Tb6yzsMWLRrGfW012z0KPhCcJwiDQ2WT0LTEkDD93sGu48V63kIyoMAaXpqY48A
CTguOnUGXI+tRzqehXeGV7lDEFLrYIlpGWENMVmHBzOU8TavaKiaNpyNYboAjmLz
6VSWaqyc6+fJBDB7jHkCl8PN205XT4/jNDDxGTpyi3buuqzTHesWIzpPOH84fopK
4olDHuMyUS9DX4xEhfFrL5JUzXQYaYsvZepKyqzXnuToufUKftXKqnRhkzD18TBM
NlKfWbhAGhpulb8Tnz6lh0sK3vNlg0s28RPPdsHOSKrN5oVUjDjIaD78DdqauDQ6
ef4XSauxEWxXLeFDtb/Ee5qH5CpVPPhOjPb/58sF6f2ug6nePtbL4IKXje03kKLH
QEGDfxeq8Vs4Go765Tp2WRtDyNGRsf9VpIRrn3LfkXjoD/SIQf8yP4kfhnf+StEn
KG66CFbrExSyEBYz6L955kmqlGLk7yJ0zq6f1HBvmSzPGe3+OpdJomfj4RWLzSoy
0MGXKxWKG45pIuUlaswZkmM8RolyDFd4xB+pZGcyW/Tt+Nam86yTmHHrgWjOlWMd
NNo5Tnc57mVmTk8aWO0eCEBIIlTfsC595MHSafsBhDnv8fW/e2Bmv8tolyZWCaAC
oKUrOyYYtSAcbtswBvy+RjJVSVjD8bACYGTmplDVMZBzC7HYllJ/gPptHCO80bZe
FKnC8GKoOD3LKEMTq7pWMDrtL001bwWd45+uq4mcQGdEsakqO4dr8+Cg2QJ2hoxm
GEEY7P3YB2lCudZPLHisHwnYyjB5FFKgguwJ4YU3RVWRf0u4v4nw5shI2JJ7wQEN
6krKda/iCkyCQULJzrY268GGX14jwN0Vyx9yGITT1Ws51GMff1MTZWzTRhCab9ze
Ea0GbQDSHupmAyBvltvZM/aHbe1nbPsvF2LA0GLp3YXaRKAJYAIHExEoC6g478re
58P6oFRlqQRZcp/m0JQ7Y4xw+Pj0pOkFPrQDbt5FM7oyHKr5ru+q0UaPL2QgUZjj
xqeW17iXc19AmmDRsxVtx8R7mGF8xGtO3buEIStla2ivbVHcW9IWsYLsZ+Jgql5R
Kx7lv6MDkTYRLC5opKorykaamJtazj5Y/dXpXyM9y+JroMtrA1CKBy4Xnop8mDQV
chg7YkcDlV6VwR0ucGrfff22luULbJkbIgM32zK5SEmzOND8m178CSZSbRNr3ACV
7jddQ65Q+1EIKW0IaYMnCT8kigE2JV0u22pKbr3QInHChOoqfFrqsEgnCXj92T7E
5y5EkVHUHeOOq1WhSwuPmUCFnh5RcikDJerRixMp/yXFnlNsve2wJ70gFfeYvBo+
2DV8ZXiUUVpwb0ZPzYRaihgeJFYVP/1vJJIlejWoP43d5a1WSf9iCAO6OoPFD+5g
6w7tnVaJgPqO17uyVoTDYftUW7MKkSd0QYWE3qXQsd+D8Li0reGBRjFeHNgAwlId
PEuYtVz1cccIxw6rHAXFiWvGbkaiRsPBe+WRUBViWd/17TxavU2s2qnQDd8HQt5p
zd5wrAqiRmPlOgmdwhIJzaMvdQtox7ISmSg7yWOoUyZ9+0+DN7s3CPO93UsX1c8P
JuoSGOGuuuRjjpe+286m6i2d0LxMwXa2IadrWEX28IFnu9ugLC3a0X4VsLhe0EsI
d8bnnAZbGHsBB4NxffDEwv3Hxr1yFTh1LcDRuhkqMK2qbVqwH+lYY3TMjLx0nn7n
AzjtLTYW6DdIJAKgv62D9O9Frf7Ehuu18BnFyA5/+SiTVzcrRVd+u0G9CZbPwXmc
3yu2CrORE1+coiRVc0KexCSTzZNS7XobjqS76UuSi5fd5RasyNL0m5RBgpGwLDrQ
DY8ZPD4Pp0iEvAj15CPz7iKjepH0K99+rJTNUe6t2uD2XpbZu8FwLzeqh22UveNo
XYCe11GVbN4qN/cEU6d35gBf8VST8TLwRNrdc9KbAMuos8iffrby87Q4DA5byOxr
8U9E8waT8cwDN7vc2GN3415fyLALOEFxwbBkblNTOTAOm9zuvUGSorzPyaU5ykPM
QplFlHinT7B7ukQtSnCeBa1eAIZS4cCMaji4RT+jYIbUXudNYhwpmvxRwHsC0gSx
ESCPE+kJI8HzAQT58fuzo54zAkwXHyAB1qBDsZ7Kfj3aAARhTf3Lya4885D+vIzB
xmNBLRpz9dz0Y9zXc0QqjDyBAEhy6CAcP7mTQc1WJCpU7/EQe59aaTv4LT/MHqZX
At5z5tJVPuem+4BI3hBhrEajsBVoo3l/pp8JWWJI+TJVxW74NTQEKusE3a/dgnR6
S3mLYXnpRik4SNxeurhmrop1Efslw70Xup8jXd6I08TKemgolzLVDw60Ip9nna0m
KQWC7lpjiPwsQRx90HzViMm//lb1rtR+s6jdOxKXb53HRNW2YyFxB3dayjaUI20Q
qZXpL4kdlxI1N3dA2JzBPsDjbPGR3iVfJgevHzlkyEu+5ZuyczvfcqU9c6HLFaf2
HSgHB4s5NrIlxuLob0oQX/iGaLh4dHOvbicJQhtsKdAVVXHkfTPGRojKMucQcW5S
xbfw27l/U0DjEGlsedb0MvGz/xwxLHQK+CUlT8Pj5bJ4ViYMEDFXGXk92Gz8fNEF
zwhmkLvy1AXjkuKvKGcIO0KNHEqRLbBAUrVKsj1nblIrUAfCgQfCTO9InJ4Wyket
q84SM91aOwX/0QnZ7Q89GJQK6w8MjHxqZlouHKuBTov/HN670QtNu5jBaeDRkAsI
9zm7qek1RqXzX7Qglk5+LNfgrE9jBWj5/IrL6Kz0G1lWKI21S7Jb9PiwT/AdkQTN
lf6XukEfZWy7mauFDHB27oSL5qM8lgRl4DQNQpOBxbPjdfpVsAGcmjnMNon88gRF
iWuh9sHmcxpPH3/hORs+atf4lNPpxpBL9J2DvmQP0z8O5/YCl59Vwq2Ir2HnkDbd
qU8loBz3vMBNJiJATOaV5Y1l4uZ8Idq/KAzTixSH9bqWrTTNFPNOWHesHYJin6KY
nvbGq7PWVy6iLpQfCBCO3v8iUMTYXUagpNCPTi89HmTmZusniOWoymDMvGtddUjw
OiVgvt1n8a/LZFQJm2Vo4YuYrIkZDKsSLelxN2eXt0JAGDAnd6ZsusPk4vis1YIX
X2k8HTKA8BF9Mwxnc5GGGBU5fYBrhFPrFNoy+aToIe+IhpHLA6pS0bQ0hoX65AYL
4lik4gqpbaWHmApkNLaoicy9wVyqp8yQTNlAC1G2scJH+d/BJtAaeTxZbDkztCeb
JvHMlpaSR2ER7kgxsEOf2ZeD2k7kBPCgBLMeX2KMv9bwK7PS5BHuHeuK4ObKe/6U
2OP2ixnD+8FBEY41PpBaUoT/pkoEv6rG3f4+cLMFF6BpxjzwtGAdQr2AwdlUbmj9
XBiEUIefVBk2mJLBrqGdEVQF7oc5S57Tu7f0CjclK4/I154ZUq0ENAT63hm3XrIy
lZUoMJhnMuLiAgYPmmMjb5pLwwNVt7niqZ7gbpEqalB9W9Wu2mDrXVbTxAfUr3M0
EePBiGxSy7RkNbG2FaEplQv4uao4mBQ3LaC/+2UyUFpXIf/4xngTmeBMkWAcCHZf
jgG6SxeEdTBjTPKdZSqH4ygffj4bkepljvxDNGPJlRZtwmHM4q9kXTL5hWMV6dK6
Wl8ksC+ZfK4050o60d7HwmA73bs7fH6JYxsMGRTe1tT448xqkZ4DUtdsuXk1Xz1I
vqkRjMM84To3tU8abS5+xaDqv00z2ihL9yOwOHjQBConoecl2atMWhVEo/vCKfvG
XcEH8lztM6lC+g/rENFsJd8YX45UlHnHu/1vL9+mLiV7JWVgT+FdfNVrXP/pLAmS
kvvuGuir3gjwX23sXaiJ588psP/dI11LfOTiBK8epVGJ0UCdW1R2zO1LXZsHf1aL
mLbxamR6zRa3+1b34kOXFcH7VpAFPa4fxVyA/UlHw0e9MLo85SjMuFt1QU2ua21y
+q5uGcLmMRBTN/pZiFyDEesVhBtQ9iqNF2jRSrKXidUpr2QLLmAEen5lkGfdP1tA
iLm82JtSA4BEWsiGqLiKJvVvdkhWq6k5TJrLce4BchDVAAIQGwCzWf0YXVzY/mAG
ym/GQTlEDa2T3016/WgoIX4ka/aKS54rrZ0h/jRNslOhmrU5KdXK6jxozYc3tIn1
2Nm0uapwyI8x58Ttfltm+zC+OTaCuLxekyIYC4adge6FFRSJIcrdigqWNhkl/wM9
DgEy/k68qOFwYY32Q5qoZAaDanG3tG0ugrpDBwwD3/Ya1mC9atYG1L+aE7ncgKJp
JoT4kupk1oEYIwHdTtaZR1Ng5NgowPIBKj8XQAY2PQFL9jX9n86zZDbsuEgy1k/C
rjcxzrXknBXPzIYjPP3/Ebsm8KVG/TL9d7HkrLIK6T3D2jDcXY5m433tnKEstRC6
31p/R5ByoznEvP9/Qbev16Dxy3cEbNnNxIpB7zraTHc2vbP3LJ3HZ7RZEMTHWWuF
U3PwHju19369rHlVhUVENw+4B+xkVD+z+B0NDFKIRjrhqWadKnU6lSyak7mykdyk
nhafaPXZasySaxIztrwynY4C8NW+y8R50VKnwXTHTkmqCxdFspOxyOzgagdDO3/s
tb66eB+ZkFzK8zPGpvZG8HwobI5cncNsPOpH5CNGiy06SqjhfOyVl6Af9OABi/0N
WDai3+pMY9VO7F8oRtRU/JBR2PCpo2hMWdt6zsPcUB5RcglRJ9nCVeD8YgA/6e77
hB5niE9SL4XTpyhv9x7NFP2xgmQnwrlNDHd32B2LxlsALa61UOph+cFhnT8bI4ZI
v5p1yBD3czOLv/9iD78+vLWtSTTZU/pNV4n8XlF+nReo3bx+XGBMo6cR6TgtDvkX
I2DCwzho0p16WJMTQ+1rDmrfA1CsSeUb1zh7gfPp1TWnduJUpwWlrTICoHcSibj4
/4eV1bwyiFpCqkQwBBSI8b+as8JgqVk1FdoXEKUYXr9GNGY3xsuNvZs0FRX71Jl8
U8LG2WTP2aH2ZN2N2Qiqg/cCxySNucl+cdLUBnJ4AlyobvqjGpQL3UIK60sNJDAe
jt/6avvRKUT06KyFByCiiky9V9QX8QY1a2I8Zyye8jrM4v0m/CC5J6MSjg+4sDGX
wjJd1xosBwJJ06M0Vlmu5tdGc/8PbmJ94SRZQEmlb9lHkC3mUW1qZSWUsRgG9EG8
8S3gywTFuUu2Ky5k65pLGo/Sdrk6DG76JLGLaXocSytPGWZE9VZPcuO95QeIDNLn
gEVoErA9cfDy1rgLRzzvFnQRQBExZb1c+k8JiHczExgMU4g0+cLnVQnW9I4Gn81r
x192fQl4m0FlvzJ/NBnIvQMcIMuJRp5VSPjmTdBkRvs7vW8VNspVPrO5E+LfW7F2
inqb9YW0sb2Sx/mVqAD5x/jOJVJ5dFUDxjLtBjHIpdqEtgSrNtVUGRtBk3PzEEro
LJ5kJkWAnCpGNXGGvTh3gBZM6s5/73DJNiR6wtl6RC5U1SIrQZ4F+1P+HsHkx7L/
UMy5k8+MaYs0I/EKHDfd8IRNpnflBPHC1HSd79Hh+fmpnbb7I4itbX/W/oRUpry6
28gUs1Y82HnDamGB5Itk8tAWGKG1jXBT+dTiMj6lwkRFawzyrZiyX/zRwHe21JWs
+ssiIuE4kB+6ghVx3ZH40zvnxZJMm7a/9RXuyaP2rz5rgGNAbXDz2lp8Kuu5C3wI
ZUop24DYQ+tv7ToDTC7zcBZKyslTpnfz0VSwBSI/0AgXIel84KbaT3pDoW82/k1p
YenT2aMob5KfhcVvXYeNcVz79aZJDuhxpiYo8Sr5BeDnzoujQUwXnWh8yeUvAZfa
cfH0Q/ri37xwqVEJpuYheIn/QCub1hY3l4Q85G3/Zz+lA44eIjiXxKkuXH5+UNvV
o/QFELtl8xg29L8LWJYUTxO4ypS2jEsS13ZBP11smeRluQwlnKSWUkhoXCO9kqvy
52iQpswoapuK6Io+GRKX1cOfHV28DnCyeeO+k7KgeL3ghHzYawTOEEstpNMkwnVP
w52anKF476kjeRdpGp/hdNiP/Tp84bW2qDoRCQIcpSZ8qwryAC6r2bK0jvW6T+kv
rj6uPVy9smXKM1dHkmW2mnU3PvzJ4VvB6a1uTwJwvepFXLEdbE5FrIAFMHp/2JBr
oxj3+Blxcv7rUcWEJWe+4lq0/eoMn+I6LogTa1j+OIR+NqMq5vW2CD0oMiHeP9bf
xct8nFl/NcL81xY5KoVrMVYTtBo3UZ+KA474IZVdJZXcUgtIpPo0AAUz1Ng0aIki
a13ZmCX21W2FlNuO3javQ+ipa3JNFGXy9vMGb81K5Z5E8M3t0WpJmqn1iwq4aR/4
d6CDiqkRK2g6ENDAdHjvPtC0LxiZiIa4gFAGHk1HEzrbpAQ9Wjw+/l9Ucx1p8BQX
9GPxiXle1nQesUyaBuCJcHql1xMNMWNwvCBXe9vL5Y8f+kF0ERRWXLamLGtKlx2c
dRuRhAmijhpcRctC7KDKIjQhHJ9qgfWS270j6JgD2UIU8htg02XOdL9eNlhDHjIp
E0cJ9VKJJrygXLuoN0VoPCc8NsWfWxW6MvT/Wh6PUXnSKc+Z31mu8gcBjcMEOOD6
/WqZ6ZcPeaOrzXOz+oTysyPNoOYB5b8NfGrucCQOAHMAXgqGP2pheM80oarqejax
TZ+uwa0WI88zkYKpYkjjpsu8hV1tbK/1sRtXoZJuC7AFyDWfCnVhAa+PzxR7oNdR
1PHsjQMC4L/+A1ILqiF49gFtOSUDuj6UU3D0xOvA6DhzRfGeYJzqc6vIxjzNIFvP
Ju9Z+sU+SdWIeWlpiBHTUH++s+FDar/lj7Ut1EgeP8HVgpMQPsotjdSf/YyepBDS
SGZwCLuATVmBBaeXjMrk7O7/rToxMRJP7s4Dmwy5YUw7UaFcizH2d0r1TYv1YP66
d0Avv9wHgfvuqvJyrxuj2CfTosNtZ6G+BV3zqMwqY8qg09eoTk2bxffSFXMp+oHk
w1TiFLRu1WZBKORDzSPEpNe24gX1rbcgqQfdZzg8q1d9JXcBkly496XKvPef7aPr
4FupNW8rVSDSMyFBNouOqBAgeCq33C+304w7aV+ospfmE8SnnmVrqa745sTR2t77
mqa1uL407MhcRoYsAl9w4L8ZD8CGklRiiu5Y7loHXhxxCs7N/ZTF0HdiaZMQF3sy
fL9a6HTlsVhngaNLo8ggedX4IfHhEsJ+cj+pVjTQIkDCdJR8CN0dxjE722s82U52
S3DBNa0nvbS+m4+Nh2fKnzdg1MFSZMXIE+Ga1O9IYopbRa8JB2ANTdg+WtH+Nlyl
i3dfO5AIsaL35R+1zIW7xktCFzRpqeKRI8f+Sw+yJ9Sl4c0TYlBr+m7ELZaIxTUl
gpFvfdf2JpRRSCUp2GFvy+swKlcPOX9fNsLrC9A/qqPmyO6xkgIu5TGAt6zUu3/a
7HyMlxt3665urfDTgwBYiBMe419v2WLluxv0Y0wbskOerQ99FwnCFGuqFrqFKKwy
E3gOSO/+TaX7IWtWOvUrhXJe8nIx6qXKUyNmOoyGXyfd+d4icyjHq/Wg9JVsV/1u
zG0IJTytLYHdk1sXrxzlNmD0cQUO2W/bOHvDNrebkd8gTWBLMUHDbLDrc2Go+WGo
NxsBrRAEMAkRhxnEhYDar872b8myqdlTJQMJMibMqvvMpdJdVn68qYJWffAzmc0I
mK47C0s/+BgpIobCerfxkLVPrAeZ19pzOoswaZr68HSD3575DAYm1DHdcloB+6Nn
HHed0pf9udLhem7C5Ate5Rz9mXZ3x+qoASDPEYUjHJyxSvUKTLjKStRSZnZDBska
zqJNVwepAp0QNWY5W23tkHSCWuJeYewmCEgOt/LfIfxxuAvAjElDSClARNtbd0TA
qM6xtVAHqZNeDbtDwOOm/K6uX/AD52y2IUD6Y+wM95IaGgcZz2qsIeTJPAjcNbyO
423+y69uDBa2R4Cy4xZ1mbG8Z7fIkmh2lQAixEDZ5xKibCmteS9OFziUSgzpEWfF
aC27H3BbSAigXgProK8LWs1VNqCovYPouwpr7D+i8vgSp5Ob2Ff4HbBPsxDSdLFs
/kUpph5uqQCKv75JM0CPuK3T8N4y0uyCfgznSlax1M20fEPqWuJxACzNlyJ5UgHz
fjFjI2yt2wPW/oB96GQk5lNjeuSLlWZ6FGdmw9GDH12pvdBae7Cu9bzxaIlhwesL
vvdQlgx8WLucVVTbSqnjGcGRlBdnPQ8Feg9QCWsNYf5r81vuvaEjyeiPKgaxboTj
e/OaNuywqShNqgCV5Zj3f7iLMA/LFN1G9hcRzGr1A5pSo4wp59z76w9aMdD3Gq0Y
KWIypHmGEd857vbwDCMTz2iTl0cx6hSGB6OzgvguLetmDghHQ7BUKgDhyAtJQClF
Y/wAwOeiOo/B436cWaB2Hk7EFrywIkXYRwiEbr21LH/VyXaAkpoDVAc2DZFbnR7X
uIwlOdmmPo+qUONV3wxQlio50VyQxseZz2AJbVp4GFHU9+kxqZFvxTJQ++OAfxx/
nXuQSnxj4l7cgnxS/rRBjHqJlx4zlJtnrkJUKQPdJpY1cbZj87v9ll5PGhCMyGh7
OJrojgNAJ2WQy3zGXd2XApR+sFDVneppebQVoWuLeYi3T0HWA7Ygvjad4I6pr/Mm
0Ga7YKiNKC7GrQvU4amvzay0oO/BPevA1kvAinlZMZxBrz71M+rb68Atvjlhk0YY
gJiRojKRmjEjbhZn7wR8WkpRPxIecys3qpTly6LPciuGyqAwcL2J3AWgedL/uoYA
qmLEZp6+N88f+Ri29EGzOdO9nycMk12vVz6hYZBT39F6KoCsVe2JkrzL7hbRzwc5
GNxNm/7Q7mzk6HWmsJnq0jfaXgSMcJa9jP1bpZJJjL5MMkMjAF9WPaJK2mmCfvL0
/8Ar1kH5q+X2w8xIFKxYzfn0/cbu/pTwN9pqLaKMXrnemBOtky7rZNW3HeHASG9w
09G8y5tQfOY81Op3am9IO6nmmCZYBnVz37+kQ2PUEzVn/iHYOjc7Zk3UPwwgNHB8
VKsQToAE7ABJRTn1MitN4SuIy62QGioNcJpYj+dyMWKtcHLLn6uF0qZQ8bh1CwIn
JzeWRdMHO1RuVs4jT5sH+PD0yNL3rMGOW3PARLLpqZD8kbVpGZ+WFHLfXDdl3JIF
hFwGh6vBE35XDTDZzWdKqVhGnZ7BJEIiplYXTnnMGNU5R7Zj3tgwrvm7aykY3q5H
vk0w7ybI+Q9h8mwXieYeP7WpnKn9vnI5eNoMCgqlSoVYKia/0bhMCr2oAq2lAJ7R
DTqL/aJzilZ4UIXpIDMpax9jI0AmgVueUX7CfkWXLjxXqHW2iDypuYuPIbuK82s6
qeHDlrzlw5gzDJgKnZCTV2xkULGq7I7Q2lRPjx3uIW8blxU+XcLa/SflbO7q2ysa
B/z+hVUum4s/NZsV63vFUGNTSKG+NA4WwjdHqO6eHTkjGR24odevXcHA6xU5XidM
OUM5LEzmoah/dKrZKcMUZK7NWGC113bRRlBuWRY1DCeAFhmmGCJnbKdzZ1zJKViH
VqaLehLvJSy/Mucl9xLOCkNIDJxiURuEQ5Z3G7Pl7khupelwg3zY1sK4/kRZVNVo
umxp4/ByXX0mkHttD7PQ4dW9xSyoRVdwndyr4nXzqIcV2ZUHcHcw6upm1+T0FX6a
nCRPJkUbKMTFGtfy9KB8bM2pRIZCr+GqyRiRUGIaSP9M5pUyFbOEpDRGQTxJGb6G
2mFly4mxKEaJUylQPVQt46qtMNpJjhM3ro6AOMIlRpv+rPVeioZXOa0pwg7ZM6Ur
eNR1ZHM8uvnxOZnorK77YHK7O8AOq+Ph4777Bh8WOIUe3TMDtu6yRXc9p8CxHt5p
ezpEsZf2gdETA+rjhTHOninDgZkehhG2NVxcxqAofFkZCLmdunRGdOlSG7Ibvokk
fq9Cflgs+GDFQUZXY5M6w/tvtEQ6rTpwb8iQzIaLXXIjJu29sxXSLKnyJ2kPAfmz
/2I4mpU0DpvI6iq9w1oo/9MpDrzRlaNn2GfPpjixXiGCWRn2uyBLK0OioOSPbp0J
QcD0TTlUeU/cUmumskP+hf0cED0KlcXF8cqWeqEfMo9UvkP6dopR2TUXLP7Ugcon
Y51F+kLtDEfwWWDMhi7TYrbrxyqirUEWKEGlZzpfk3KTrrWIHK91SGs6CUJIKYHZ
mjXNsOaIQ7tAhE9fPHIimv8GZhXxlQdshH3hlNPzBDs9p0f61DJapmbdn3pj/2dW
k/pWGT9w8bD36lhS1qLA6+e0PLw+3YqQx0MKK5Wp+bAOr7HrP5/9V3DtnuWjuQSc
nNHYsE8FSgBCKGw536tofTDt0G1AlFs2saBC4d4mutdM1IFdo2QAygXjTibtTSzG
oN3DcCf34AQUl4EIFQcMHqiloymqdHtydcbsPV12J+teEZJ5tGHEPAUABwXPeJSC
od+RSVOb2R7trCjAHbVDPoDt8Vlv8qzUHjlcCWbJBTFDr3IaY8N/Ot0jANvpq/WY
FyLB+0dRFXeC9q+0qTIDBPxIj8fOkHk+NXWk8xpSgLBLs2tLIidbY/IrOlPabwJp
5VdaHM5uTy5EyI469VQ1YOSoi3paLAEMfJ7ozFiVU047V6cYSALpcxKoHecNeoE3
wx2ZsINjprLMWjAglNd/6fTK28sDESoEugsoveX5SoM+iZaGTX6l+0etonIySBt3
XCsCuYi4mswp6LyTYaEwGc3q0ZE2hZ8N1apY6rYLFnq+I2Gm1bcc+VprJu3OzDo3
iKcHdb5ooecYWuykFs8V9c5BrhusVNR8y5yJEVVyoJ191e4hG4EGGHKRfebIAQZq
6lhxg7KcVcudfD5QndX9tIvLkUuIL0E+ohumpJ6oJdAOwpoFWqLHZpK7rielbkGE
+kUiSTyBOH6hj8DwqHMn3pu1q9eYm91E0+0ZVzqiCVJK01PY6KE1svidN77d91cr
uk+CfXufYMH8Gtzurj0lYj62jcpWeX6ko33Vw8yDA7knRWmve+EnXGBvEtdcxehW
4+VkkDrQwVkjL/XmiRzZ62cZ7PeHuiuz9Of28LSUOzBpKmWZxdq/5IkY89qydRZm
Z+liS5TXXCIgv/PsgF82sq8uljRRv2ds+0abbV2uVpe0VKEukYFkDLmEyAGCMRyt
JuQrwhd7hoOjHFxeW21jQS4/nMGc5h232UD+tq7E1L3BSaAdAx3ofbIWb8ee3OOl
UogMWF+wjHsiBcag8n78bI2HLDjbQvnM58+8H2ojetJqS3skS8fkiR8w4uPndfSl
6/NjpKhRJTZfqFPHm9nle5FRz2BwtbVM0x0UDQ1RxQcv2RAXUesvTPN759sM+azF
r7jhBtved3uBafRSnySWro1ahHNO5NCU77tLLulc+05xTTYQGsdKDYoERa1aMu59
ieWpWnjQhgkXgcGIOisIWYHpogAC62+Ur5d9V1H6liCfJCZC1yU+spq0p5p+hQEI
vmQh7QwLXBkanKRARfuxUSjOPtV7aLPkzpF5lbMq1inM/iZqJ8FqJXtmjm2EDzcN
uepTmcB2+SBFf65eJ7VUrYDKXxsufbzGAZ2XbMisfUCMIfrYAc4mOym92KXocmMN
V558nIVmpyMNRpgAC57slUI5KTpoROBZ+0t5xJUgXbSR/PyZIObQy7IdfN1roMbh
U7lFzVb1YZMhKQFqoaCZenqsRX1Z7vvWBgIiAGo2CHbyOxCvfQtP9TuPOL+SclJH
HZpW2XfZ8dOth3A/comcytKpYaKVkSSfRpRjksTNeXM3shQsAaarYOuMrOo9J5IF
e7uX6Uch6+1q93F6mie4igwHzYg9Q7Hoo4Ta/Hr5DS5A5dcSCG0igxCv06xHVhsZ
8WPtLtq0oZ3WmgEtutvGia0Suevn5Y0v1+1NlBGOTwUN7+yvnYAWzObFyRLFwBiB
m1idBj8sH39jPMlJUoJfavpThFsYjgJAxQimWvipdH6CYfVd6AMZbtWud/i8hknL
lNitA9UBQk9QtYl95O/1urFE/uRjhGoeAG7UkeitqjkXMmY+WD/NJtuM7r0/xgnS
/7YmoY7jL2loNcSKi5PfmppJ9PuPjshx+FR8Icfp1vqvZi2yUGR7U7cNBBH85AYO
ODjw0Et2UxXqck0ixro4E8WEFKBVUQiyzqKGzzfgettUfKEvlcXaRij0fZL2ePbx
nhUWkrLHNdBZR/XP2fSBrpw/1FOfLxJid6FU2L6bN5iyLj9tqr0ArCz0SgwLXOhJ
I5ujrcXhT2IWLA5O5z7FPmJSeARCoelFxjA74ybtdopy9Odm4ws2n1CmhvnKemlz
9y7XsZBxpPmHYSRgwE7OJbqhkyqDwd8idO1X5R212NpVnSeoxUTJ3Jpt5a3zjFBa
OMYyjCtkiMc/1tWjEsejAUAREy8otWFagHsn12IW7PYIVYEr4/eSQ2cfI3lkfJNr
urZspx4jvfoq4xTzWp+lRfWBJowOThm39RFTiSplodGS1fDR1DUz6GhM0DKhf5OS
Dpae6ChHOJE6TdMURhfPOaDKgl5z+9n7ll0vndrAc34jTSv/bTzMOsND74JI05Ur
Zm+JCJ3jLufpLBRRkCYhJ5mB/GsHUPThoEtewo/iRho82LQGJ5VrIdVt2YSr3kqU
9BRvv25hoCT+FWINyhLOFkQXQZw7PBf5ZNcwpRIgUrWBDkQfzVDeQlMMQ++AVM+G
uFrN+PIeqZ+WOV8U0Yeu45zCklJf6xdbjP0i+iwlV4CIowt9V/NUAB7RTBcuuFSv
sn5dq4Ek38JCZ2lneOWRomaVN/5KXoTYRvNotRGhrjdrM6UoSteBIvH/SJQh9OuW
PuCO+LsUZ9xWjqiKM4wppK8+4rOMdyfND/2OppXLpdTxFg59VtgPhN4LfpMVPr9S
nx5504Jgqxn8e0Ru759i2SyF7c+LOYFSUoj8limB6ZLf+dons0/5a3LLaVkNBF+q
UOwtUhPCs2xgMSz9q1gSH+irb+y0DojwKVMwjQhNcKtKBdGOh5vZpCmzxrZImKWX
ZhWBbt/c9D/m0LNhCHvi9sfgiVuLuV654Iz0TE0AWwLOKOiyGSzQ2iuWks9sWHWq
AqZRrp3sXbYLzKBW9R1LGXbkwnpyedYs4IK6srvrE3DTBuy8nP3sQ2Nbx9/k2Vyt
sF75BZg9A/OWyw/53YQQ8RktPfBiDY5/4e5PfYsftWVS309UWn54Sa1PzaNbf1J5
zQmXQPhTaGo9LnES3Xs4KuJ9R4WbZPFSUzMZ5JVxMPDNMyll87Jt/cfsJhnEu4KE
OjKGe8YvqRgcMElZS7V/RwjGJ5IXPYWe7HEK9jRxafbIa9MZ6j1Jscc28vnN6+FF
WBKWvd7UR7dCUEhv3oZAj6SvH/7ch97/p77MIrTQOwK/bxXAwdb193adXFvoN0ll
eE+cLMjLW214HhuFxhs6hGntTr5L70Z8DayW0933IkO34DHKqC0NXX3f7xwRJFBz
0IPyt7Wl9uQedBOWW/UqD8Uw2IxEQxqllpPd3aiVu0/iSUSXqVSnbZiI2X6xq0AL
1p7157R5b0LCT6qbpKIBarv4N1l4ALpBo5U2mDilFUnFVxmW9EqSqeq5FkR2iLMq
B+mNGojdnTFU78p/ZOU4ISjXHijBmbedCdTfGbEP/FRqesSN/K2zXCZtC/DnuFQV
ysqh0WoOENjKdosLY9ccSGR40qiUIcN9DUYqni44YvLgh+426MO7VqxjJwQKzaoQ
D5fB7sG2Yw+Fl7SIY1+/Yt317hmiPaHFFDcfmolDdA3kBv8T7t8g7nJ/wQUbfkhh
pvnoIOytvUiY7i1Fgr2GqaAr/jvKC48uT6v8HXgmBkrVrMOeEfgpxPmsH+DQbfPy
x1sHY5Kyxn8fUsb6CCasb7/x62gjTKg3SWKxY5Wo9i0J9QvQ6+GS3bZUakqjsJLE
zSl6E9yoiIZPBFEey8cbgu9FqdPUHZ13fwxjxOc3xE7VXuQz5SBF3w09He5KxeHH
KbxU88BLDbph089bDNfHCIKaYCM+srd0UiTyXWlKLgy0e6mc03RT5Vqq5Ypjs8n1
0i/L5uYUQvqTZ+5U+d6JbhbbOGdX/E3oXK2bdi4U1DiA9M1VISdyROI5kDk7wPsH
IBC2HzTAB7SN9gupt+LrZQUydTJp2+p664uPKgVBY80tj5CriMZO7UBlNnyo+he9
lM/di8viDUWCiImOYbR4czTK+1pmHu2nnJz57lzwpdpAs6hQNzcEpxg2JV4lOWTJ
/AlO1IOfHXpPlb8IvlWK8vJu8Tg/HXHSExkMf4+3Km31wvYH3zJM4QBSTPD6Rwl5
cQ01pUEhmldoON0rUKoayQOlqUeL6F95v8PwzRJPEyjTY2Y1sHFnuKZkml0Il+JA
hBZcjrcYv3vT4wKaJpOEhOHKDIipT+r17JE9uc8S4rXYZ3TZ5gvqCRd3E/1tdkET
R5CHuY19AlvLDwfJj+e11VxH17/F6PwMywvbxLOnuIYEbOJrjyzsMC5CK5OvoTOx
WjOBcc4r9tHCh7GUdgZGSfh1iz75hbdsXH+eseINYtsvb0OXx1WoV7v1ijXd1MKa
3kIlhtUa+UPiioAeTeRVh3qnCOM1zSx3hg/hahwuKxd50jKerstDzCeJxdmcyUp3
lf7Yv3B7nQNzjotUdawNex8CYUXmzeW1N7SitqceVO4B3X6j3xxJpw2hOOAWynQO
IIzXdtfqftAqJ3U/6JQmya6X88owrxpuGf+fnyIQK+TdI+YfgV7kWzFixKAG0eah
BCTu26GbWfNEngkCRGEzVyWkUtsKAen+jcI/NpQykmcOhSqtFHZo7S6z/ccUhbgm
o0UCSLVG7dd7SbhTUT/2RT1E+zvs8B9hGXlw8esLUpzT1QEKesuhwrR+Hdwi/bOk
B6OITiW12gYUE28WvQazGev0UcNwAzYhZCkhYZ33Kfg673lhvwpMpkpiti1cs5fU
TBA9aV4WaLSe1Xejg3Q98nKCIAJoZeNxshYNW6JPvOwQWCaQ9DSb25SVu73mqxqo
/dPlNcegkAk0JowYY3AsJIVb0nMCg40QP6O9Rbt/W/VHh7REGav37LcGlZtd2Zmv
TkPRewRVdkNoCX4Y1T1B41FadhslwM+DF+cD7cpVt74XAT2vhRMFe33nk3ptjrFV
Pcnp0af0vqn6aqoHowWiE2jHcqLFfIdCcLSCIj6NJhdn5Eq9h2vJjtLLqn9ZXUPt
YVwG0FOgcP6Urj6DL0IcaiwhPq1PEN/LvajPBBtCX5iWRaUNzWkqEK325PAUCSry
x6I2e85S76lLjIqrRyTE16DA+pyqX00wdfN5D0X6/187bIl0PBuzyUd4FFeahLOj
r3xTBj4GE63uvXk9eC/NC54Bi0982XtsWlmmW3GVdqQiI/AW9oFfKSDQWVsdNZf1
t1mr0COeajW1+4J59DtX70orW3h6sAcO6m94OCwxWdSwwaDOaeFqZ3gk2heX6gBV
L+dsvL1MoGpa15CS4IfjEM64cdhGdle2Eb28gJ30C4jK/801bwjSPiPq4gQht2fa
2D0fbtp5T0kz/zyoiLMnVK0oc3rfd16TZNuJuJGjVygRIDKyI3O1TECi+kXY9ORW
q7CZ2TLPu40+8kNyF3zecmbz9y0jMcIftXpy51GgKlBb0r/7mSfDf87ehA1qQ2XK
3/DJx4tM7JpaBEHpIZBSsC02y3ToPqoFhvGfAYs94cudWKB85X88sgL6+StiOc7z
5fvsCUHECYaa4jc/tRMuk2wG3naU/bh27iYhwev2NcmxXKslrc0BvIEhXvq1IuJN
ow24EG0dv2IkHbgXIWN+nUludenaUKZelsscbzFIEXVI7bugQoKAGgpMcKOTa/y6
BLmLspbqyMuWQKrG+CtDS/2fRN8Y9loZRyxcd54ytuMvRoWmaj4t2SGgH2wcGsUR
L7lP2OTJuCGFqnjMa8i4MeYARFvoZqkkxNb7TMC5c+V5qI7gTn6Rjsh07vEf9osI
8NfELGRjHHmpxsgminmPaCeq6CeFVQc4PViR7lXIokOm0ecem/5B/KZBYSolZjOW
ynXeukjoRzo8mb+Cvy9QtbhcKWT6CbNFAlDg/nLQko/Fkyb4n+/2v4jd+qGD/VxZ
sZ/LxM4NKkG50WYenqfJus+1We83R2rgy9BPwxdviZ1lhQY0Ttbb/gp/fKK1W8be
gia3HkHgIMYD9L434WyhS7jkAS8Q+fEK3++PG3tyVLm18iIUJy+e1HByV5CoBJRC
qSPgUwqlQ5jZ3i1lsOenno97PbauWn6F14iJ7oxbm95K0z+bBaH2EtV2VypZXejK
CVUa43lIsmPG8lIeY6aYYTDo2ysFpad8hyhPsivkUD29IjCyrZne9a8nJJ4dfdgw
IeEuiJaBTQQEMAfp8ETcHSJqfN3BpKAbsco5GNm3+sodChEpPuGGQu7jT5zZuiN2
4kLIFejdyprI82JsJfQFMsxm5ntNTeU+Mx5B9fbaKhSf2b4BR9wkVlABFPtrh3Fb
LMOwFb8/NLSLxhxLYHGoj1AC0OJDKKRCZFOQc/FEci7KAqKitIhJVIjj9GEZlXT0
uhlDlvFvhhAcOz0Ou6TtXjXMmS9i3j+bXk3ozVX4AsIeOaWRuHHGTuGttSTT0q4e
d3VVWxIvyz7bD8jz/GnRB5F55a/d+CePppUHk3TaViHZo/IzlIRQkyEohZ0e0qFI
ApnaNO6/SU+ApdoDhJ+nRGi4eqxRXeCPS0dIe23DUbgcmnFuCkW3lQgNwG/5He2J
xBlgH0LbBhOt4BMdbbfkoOw7l8uT+BT+tFGBACkyTYUe3wZg0PU1D+ZKv8pW1gUa
to6/QbtoLMfDuhlSWxDb/VVafsjcPL09+eoMYYmliBH1trdbDQIidhellGZQRaVX
bFy21/pxaulWK3h1esXy47KNrp6PUVD5Pw0z8ihGa5aXoOsi9D/ecogHZJiTlatj
vU669H00vXoLmswJcW+o51F6PbRPk3P6FT+RalAY86omwRSCgnysXM5BIn5De12+
Y8uvgeDTcQ6u6711FwAyRZ0GMxCdvNQghInxp5HF2Uqm/phpSg6CqLjcxvUuKfz8
77/oKhymckuqGoKyXyNlqLhlUm195H5BgRf0voY4U4bVeyHvOYPg+CvBkMln0xHZ
yDrxfvNlHn9BxX776OHPbFgGO1IQtI5axfYqFAOgqMQ6bUGVHHpdmadnr49LVzGE
6dPM/ZVJmHfhgfikrLZ/HamPjZSMoeupU9Z+4BJzeIxX3mCuDeE0xe5gcm5k5pMP
x9BULUqF68MDO8UrMhCJ5pf6C6IOImTxzAvjGbg6a6kd76cNTjUKGwUoqdy5EvJL
KUGnLnMnjVOaWYo3MzsMsorkODpkllxB0HycVOqb2DmiZluUWQoxlXiUj03PZaBO
nggS5tgmJkpOlKoZ+rugvFFcxsQyGe2MO0MVM9mfK3HGsE/V75B/DAvk+Lku21cu
SQp341pv7ABMbC56y0AZKlv0r65ZxcJttK81KeIlAUwcxEAkihWS4CNWSfEbn2p7
fR7L97fNvTi/fAtDHVWqzptuQ5vs1HQiVFzwqbR+sIH8ysogxEnqvS5+GqYOq3GJ
RpPefMMOEdC6uSFUzh67+CWP0acafM1+vYRMOT28O2VNlT/nVjdcToPmp/YfMgeY
gLcWiehrjx3b6QAEMYGXnpqhfdvKbAdNKGOezfuCYAPYlgyUjNvYVTf895++sA1y
vKp1jjM++Bf08AJDqTIHEE8cQI00xoIpVh8wMacq1ZdDVHsEnsMy+TfApD9nv7T4
yDA29ZmkqaiiyEObD5yJ1UQg+5/43INv5qoewdarxm/HyM8468M69jk4Cq6pwnJS
L0JiqjpINNkCcE1Pty/rRtNyXt2sArxLVMTtDJoX3b3Dp6lcpZfq0ic11PXcJjew
5/HiQ31cUsafMDuNYBM7VhFe+m+LvmtBjqCu1AVvYd/bT21yp4VY3nEPPJdz78HE
68rLCinzuoCoSAS339Q6d9DdDY34a68d5jg7XrMtdOYXtHiwSR3U7LEQ9VNETQSF
Fa1PUvww/R0WYC8IQC1mOOQjNV7AHV3xWstQuHr0EoF3Id7tuBJ3YIIDsNX7JJrj
vr1KkoB+V5QsIYz4heDPerspEf2PvUdF+iF5p42eTpzscczlKjCkvm+awKt/iTcR
PNJESjYdkdbAnhNiI/qrjFgjkIPatmMUlIBDvu1/Xk1qUvxqH7XB+HkOAAZXgYwi
fGwssFwdL7UPXD9Fa0HMnvE4muo4SHtNKA9QhDBzo3eQ+3XJRuLTv3+1Wfi7V11U
+CNZ25falpXKhQ5VcLy0nG65K+piMmUMu6CZjkcAqNBQaVR0FPjQiIgwO2JfMZ0x
ibPz4j0K9HPAkkun+EWll990tO16oL+Hp82DXv6teOOqU0r/lpeuC+HH6g8lzGKZ
eQ9Z1V4N4A+qvH/zA4wBYC42c5Cx0B2TS1F943YupMdeVZVhhs2qNPifmYCI6GF+
X4hax/NCgFlEJR6OJRLktniO0ezRWeetJGT1pkEBsJ377KknL/vNNACznYBLMyKB
opR0ZZssSpP/qTb8TMWed+fXv/2Kt9GqQLa5GJJCpdgr5d6NirpDNSvmp6PPr6uN
S64EEHgS+OC3hEKFA/YO5qMdpvXiMtOMbQZ1kbFIduqNcSZZfD8wZ+Qnjb3KiK4y
XEYQG67A4w4mkucGzKCPhQuMSXAy9C9Tj3gSRCtF/GUVf7z8nZPMCdAzcTnxtShk
YAqjzJGAlF1GIvG86t7YU5sm6R6psmFXgFWS6u3F0A/0DQDwBsT3E/jcDmm8IN+T
YkGIfX2m6p/YOAey2v06XmHI4VqkI2J3rslbmCeMfW+L0unG0aEvM9YAXDm+dMKq
ZjvpTeYEea1bqSsw8VVw0Bsmqd1q/tXrD2+yTn1l6PK91wNjRrhKisIN+vFtPLHk
plN5gsIG1ct8W709WCEmJmQBMjtGdpnoj485xfdmCz1yle+EcaEQlxink7nzZhx1
+DipF2bUdq3+nb+VtvQH6avjXRdurk+Hwg+Hsi90aEd5R1LWlfmLQd+PaDa8sM5A
220ZFgYR5Jq1SO0qoJF11U0GhBPaFEZuODk40ueM+qyLEKhz9N7381JI4VxxRV7c
TDUcCe4BYdfMNvGxcWI96yVBSshBp1UHC6Nj8tgIADgENt2Vw6pbVDZIW+B9Wwil
n3uIHwC77eWJkhd4I6Ja5H/aBQen/D689hUvQIdO8kZ88kXC652UbYUD2vRmmHUQ
lkpdZdT2tFqysHq1J1Q6Sm+tuL/fPPNL8aQe12abTF0s18GPuUeORogrr7OGO/CS
Jo7fDdqerVo4h4h0gW27nhhYXRTLcK+6WVyrEm9lQpcVeVam2OXm0F76vyLY4dKP
O4NsTE6djge7EGdUu+hfeDCkLkdtgJspwLMeqVJxVaPeTbdmGAeJd/K0frpzhJg6
t2NSZGsrUTbx98uPkXx+kJLhD/QvxTxY/IxnjIqHUIhYWp2Xx2azw0tZvgq54JJN
kmYKix/AKrP/hmx3CInejSXkP0U8tPHxF1LoUCXM6DbYiJk+9l6IBy8G72Yne5Hj
yG2BvwU+iww3kwQJHIjTTdAa+j+YfTIMoFD/Cd44FX8qO82jRnLj9ag5WlnAxYAA
QMo5RmaLvkN6s4imWZfbPxhRZOL+1GAX2Hz8DvXIR+W0MMPwWPAynKk+NbLqG6RZ
TnW6+As5cAnwZzmcmJtefWgg7Uavi88ARK1soRsO+ZdJg4og9y/qcdJPv8QzC2Qi
BvXfpFFGpMN4aHtyr6HNDCSy9bnNotPi0kkjkYer+aODOUQfV3YIrwgCiz06CJ2T
OInXI5zUKUVuk8hnr0l3clah6gXpRTKPu4XIcyMy77XtjUQiVKhGTFrfSlZA7YWn
49WGdQgs+51VTIRziNRTO3aOMCLZAIun7rExmh7WkwDK+OsKwmHeRDa8iXcWP/v6
na/CqySu4KQCIB+WoZpV6H7qyEH+fbLwybc7tbhjZIh/zy8pZYZ7EQ4BL7sqsFc8
3YHMbRWuBHtFGcCkINF1QdfGI2myOeDvlWYe+4SzKvQQ3YL3RN5MNsLJwpBM0fqR
/SC2NorEnnTVWHaLA6I2jJjgy13fyxxDbwSZ+egcJINkrAorNlMIOziTN1a7dnK1
AuYrVoB06Xh9deYzSsrTNvWnaQgPy2smlZDjD8J1m/FX3G0+H143oIc/A/LKH13e
yDd5S2pp2t7M3lo3MNDZNgYkDI0N9bNTTSZK8wlPIQw8SSdNWlFQR/JY13PvlbeT
VuwyUZMB//eflxR3XJcsgoFMRRdHn4+1XFEp9H+Stofzu+T1s7ozpHLtQjNoElQ6
2eKI4qmx0UQtbMXA5xpNWxFbwr8pLAMQ2BHElw2BJJ88XgbQwk05H1uUieDpm+vj
YZ4GCDA/X8A8Z4tPD61bxVPm1/2lKBzbMu3+ENcFNU7E1BTDzvwJOpg5+envsIz3
ubt73yZZ/k9YKfB987IEVUUJwAYgDriB0RbWs348kXTnQq9a8BwBJIjrXeqHp4yj
uUIWD+TAG3eweB3eoqKTS8hIkH9QtaM0AO+Y6875depQC0li511tbFCRByLFz4wb
3brPEvES9S/LtEyS03h7OihpKrFIseFR1ZV2syfE91gIsQrCAbEwNOFDShPybpZ6
/IOa+Wx/kx2KeIucLaEET8V+Fd4gR8mrii/aUJcPe+myGqf9hQQWUPB0VYKyteCp
8OlGc/cQst92+is6/nLE/CgOi+5ZJ1BzyOUSlceygfetz7o+lOQGZvEsJgPgGHGg
7EkaRa3LqaQ14GG0Hmsw3kcY4yN4QwZtcBqkuacBSL8SaiwB/oaQtL/wwbTf+K5f
lDfiIjhdQt3TkLoJKkBGTRwCXqy2LRZ7w1iYb6N6N+6+gWf2A5dl4fwLnqPsNwIs
G/Npuem1PdfSA8fPSi3oZ2K+exS5Ai/c/UQQbvYnPg1e37/Ju68PhNG60UsuOcCr
auWBsrNQ/bV5U5xfwE2pPqt6Y8RrGPNk+0SWTDCOUFUx4MmhKAAuPxMsXabTW5HX
KOuGscr+20UgCSljrhSyMY2CI/9pv8BNp8aT1+hH6OLmsfbODSMQQ7Rj43bZWVcD
oqVwvj7ndJPITjEmI77uuO9L51zKmSVVc/UVYcA2I4X1incz9g43oBP6UbWjK7gY
rZ57S9+3C0VkgYaCBfY1GM6WdneQqtJiRSODUtBPv4aGMpC73KanD6ikXwvrSJJP
K9UGT8FjDIyv7j7zbnAfnI/Vmxw8mIMfDP6xXjsgG3CcPc3Px9plV9NWbY822bhs
Q2ZfipZPCAo8c+iZm+wcQU6WqoBQJuHsx2ImusZKsvB8epvOJskPGRpnj104Mpmp
pjSVde8MEzL/6wbryCnAWFU7ZEoZu4lhK4QC1c71h+xm7R2GQi+3ARRp2j5gzwLd
qOs+g3X1ZQ+RRjj7VFlnk0snrw1VpVXsi9Uq1tRLalwYIlxcj2zmWKbWxBWxyNvJ
39RZXWCWQPMU9mWFfOztjhXoiNmnLgBTslaH4NjJ6StRhOvTQiWzq53I/d3+efX8
+QviydB0hjkB/xQeksYRg3+fgc1rutL04K4yayEpGN+dYcHQi/rYJIa+oLE2hIvJ
IcUl+Lue+TCJXrQIoe1agiQdn71hHxEkZNGo5HiTNEQI0o+havdSuV0eEmHnu9/i
eQUwem1FSGrGNgJbHNmMoL0Y0/b6hkonQfzL+HzuyxyshX+hDpMTT5Iej4fi1Ykt
rZ871JtaEB18WgSFoht7HQRjvNX4s+gLzBfp3wp6nvF8Avv0NFi7+nQuqBhQz9i1
PERTVdH6lrJ/9xDndkQcxVKZv4V5sM9rnGpCusNFkV5xiygjq/VbbW6qDyFeSVsO
AG3GE6vUFX5rV/hEYcVaGjG6mrkuGupWeZHhUMHOaSPBysDY5JcaGlbSgy5xz6ZL
4IVTzhDistFl0Qay4iHJkGrOhLunKAwJRq646z9x6AsUBz1WlFd5gDR0/xh7inRD
dj3EjVtpRaxBztRPtCa8C86yDCjwM2w9d36lNLh6S6E=
`pragma protect end_protected
