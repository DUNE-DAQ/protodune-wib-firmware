// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XVPxetA6NZzwJoyoTuDvSlqfdDK9ykNgDfHCHR25CztBYv3cdj/XWDm/wPoFZi7W
WH30g692gId1EreZAmZINZ7WP7bcfb2ky+6+aNNUyLvCXj9YcGeyq7bXhOEqb3FX
K18qVfGutiswaQH4emtraUyl/wXqQ0SIeHYO9UOj1II=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21984)
IqXWun+3NkFKa30y0bJkyge9NR+ekah8myRQ4YlGF9No6pDnejzhABqgSX4y/cX8
5gR+zW4nLlyhUvmvHUVe5u7zj8t2ERJj+bXHLWNJPvQAQnN9nAA0nDRyzp+GSpEj
PCcUjePQAYHfIVfvtIf/89Qpw9Mfiv2fXSw3db9pN2CvKFd+E2/3sqB4+HE3VZEZ
/yVwiJc2U9bZIV9+5pcKh0kr7+6mGwut5e9Oc00WUlyy5kCFz+VbDZwThfOgem8C
AL6FhZRz5Z997BF4yq19DFD28U936vCCfNoT/h5bGUMA5XOUd0D6iycxgpAktvXx
2FK5Znk9t200rNJXZQNmk/FUYtHDdfjtApCAzqvPOsLebCBR/T5B8BI6VKFlpehD
UNUW8Ycn+IuCvv4GKY9PNoTwzePAy93a1AVfQjJ/89gM4MhC7j+FlM0dYcwirYRE
BHsSwO6vvs8JEJolDIIcVGxDDAYYdMZ641FekT0x1qlS/we6eq7QHqTsodX/HO+z
/WRb75nKwarCWuNOrCEPr4OjEco4C4puacwg20CYS5pBEoHwG3zjut6toquUfjnf
BVE1e1lTMynowpBTVU9SCS5VRma9bQF0IsrG8wnquHsPtGcAJU5oib1BG+M1x5bv
MDpnxf+SOj0Y+34O7gotfnsjMS5FItn/VMZgeV7iAdzpHGHhzucXDg/1JCznDq1G
4Rv5xNOQm7oO+MQVs+ZQ+us6EKFLHtWjIRREGTatXMVieBSCSvQ18qtoPLiTc+Wk
SVBAwcOUy0hPDnNixGaIyfp8+cLthxWNYDES0SCxFjMTE0ZHF86Ep6u29OqV6XBP
mUu7OqASQSSglSVORBi9RXwI7wTCcc9GQ9o3Hp4RyFDH3MvB9WtouWzewcC2rrfI
DD6fzbdaCprrQSP2DO5Zm40akh86QleB5tYh634/bBh0fPBIvxwWVAeljPCd6Nmv
VGzefBWjWn7I2/7jHK984FKtDP/QTofBmQagYKmdEJOYqCBxn2RWVEkuvKNkvUi0
r1kXOA5D0I3NIiMm0fEJ5w0imygO2XJJ+FTcvjF08AAUwHu9WnRpxxMjt1dWVIE9
d/2ZtJVXWih2tpEYFrGAMv9FfcmLKfjLAVb7fUlWUebEh0/X+cK5WajxHH/HPISX
yCdqepJ0KR7w8FglTFr7cO20QvvBqYx3/tcl4A9q4vOHUq1358pnidAV2mEvKSyb
I9YM4vlZT9ZNFGYdFZQ6w6BtkFrEHmJrhGPVe5LNRpR9Wb+VoRv08sysCMAON4KJ
+bZLG21cvlmnJetZ3I6svaSTOlsMAK5LRYkF2PmfvVOlP1+ANGFZa0K/eJKAUTm1
+JqpmBAO2fISOMh6yRZuxWz756MrciKqHbITYStV0NpJngB3SX1o0vMI+NH34Oks
nUZFZw0W0zG+JhialPrqU+ml4igTosYmKA8CG3BSBpcwMSmgVM4bEepqBtzac9TQ
CZZHtNguMApz6B1V50bQujADUQdf0ZQ78vHqtWGkP1G81UhCekRLmpSBgz3LlhaV
AWVF7pdkR3SgtqzVvoweDN0hDeI2m0rocQdFyJIROgefhjqtHP5dvBlh61LZt2VJ
cNVZleOfPDU6GdHWDXlktfcjRuYSmU9YY5qFaTJcOC1CqfzfJ0Mh505AKJSh4WMf
YqTzqTJXLjBrr0XuJPZ8JCKWzVF/vDnNtAtz5b1SD+WUhAyi3NPDqY8GBLACrEXQ
4S+A7nir1Q0Aq3IYCKre/RFiCtRY1LyKfH8J0Mu8HHqVSPRLWROMd+Jxh7mfXXUu
fenTo0BlD+2IH3cspxL+CgHCOdU3pWAjFHF3qpGBikukDFnLn7xCqjZLNqQrFKzk
RSwOsRP5FTIZQmMSTAHavZFJ29zG9GjGXnH4ZD/SaKYU0cDNLjvz+U26sDOfFMlQ
3caKYX/TKSdFmGf5V3LHtrfq2lhwSwMnxL/t3D4VZqecgAIuoywL3YMf4eonwMVc
wBPKR45Pfv8bszIaf1tszMxQN50AJeJlh4oOLWU4qX27OqsVAjLyGRUgPDja3jip
FCM4MP5Yguo9keplMAobQuGEz1QOKT0Ztoah3sRuYLE3s7/6lh0dmUqq/Jp0GPRG
GyvYHd2tPSz3hX6kCBqNTWbVqkt3ApWPAFgj6NbEo/dhXLb01ohV6+GLl4QSQj6l
/cgLVJzE1JPFrl+inq5P1fwAVwbXvDV2FDR3beQMO2pZuamUhI68bTqMLWIkrh1s
rMJDem0U0rZ5PqQPbRLIJeEvwTeOvL/KmZxZbg4/Urbb1AgzCy6hN23eV2pjKuZi
tAtvfiokvbAx5iEgLi2UrAtEYbUkNn/3H04tgsx1gBuWTBFGu3GA5ZbI2Wp6+pUe
7eIZeGZHlM9pi6kttqv4lKkZeOg0Ix/UmqFImGu+gN1NUyI3J06BcX0tngLO9tjN
SqKri86dAyZ/xyoiJ3JCKDc+qIMLgWrTSShqN7/LBmf0DGR0emj7edFnvXYxlM2z
g+3SX/iEXtNBPaPGx/KD3zsDV3KrBJuz6lEnXAmiilMyANE6nW5nCzSB1d8OK2ZA
ZTEtX81nJWrGFlW3xz0mZFi/Knf7eNCMSzrNTF4R+v8rGtHxIYa8SREUqKoGRwa5
/dw3XzMj5lhylv/8WSuogt3Bmysj/rGISOhr3UB/JORW2vgKzBUclhEtizl6DSK4
fvUhESAP6QQX/tOQvk8VdLCb0anb9RuXbEnk2oC9/FoQBf7eO6xLrS4pNsAfGpgE
pxp9uWPqKaPRIjfkxZQHKsIK/ufEucV4FepnV7RYJl1arZNmdrSqFcP6462QJ8Hl
q/U8vINhO9bJWpO//gtbxJJTzg0WpiT5TnKN57a7oau8vjLz+0/L6R93qfVW7ctQ
gLPAW3HgU7reQc31VhvtZgUz6LnXYD2JwL/ORPzozxETihumvMGU0o1iLvEUOyNQ
Nt9QNsMAnuMZfvYG+vsnahbBLeunq/iL/U5i9k0dinkXdORv/VpYVn2LsAlL59EL
cM7aIAnutCN7fjbqPTf4HRANmBSHF4yv44+n561xwK+Unq0CHevkSuYLO6MovjUB
guqytQCRJQ5m5SiGm20ycO2PO0wSGg9lOxd6Qy865taruueRph8UdEsj4bZYWlCT
B7muLpCWarS7f+EFdeSlvhQWyZR009lPen+LdAxcsOHU3v3fgCIMRkfMvX9Z7JGG
1w/EtC2s5yGtE+B8GfnVvP/YObXOAY944lqXpmtRQnX+C7/8UQEu/hp1YqbyZDdF
/nY2YpwW6S2nX33OsimMyftkw3/1A1nrtxYNmuFHUfF6PMj5oPk1ZXproWWyEVHs
cHdPqOt/dAQnUhyq7tgREliixfRgeBrMT9byFal1AAhQuvxebvH5xaZ9MJNemiN3
QT48aa7XLf3BPKpTBN7l410dFlm8zV/L/rUKaF6NfOe1k/XAPRvba2chHxTzvChf
692QxX9iUpEInFeOGbupfVkyDE3CB98mFT0XaLdGn/5QavYpJRzoSTM6a/HbEtRC
XsTDWcidnJKbOhM/oB1OAf5OHoO47WGuHqbBHSazI1pm1IcONMPgQkbEbaqjZ3eu
lxQ5zmfWgrsa4Zke26SkoJhLhrJVUNqjrS7VaOiqb0TcQa0xEvbUojDIoJXzZpZG
TDLx8mpZoPbGatLB8xjooEdJTkwXQBc4Sdrepxjry+XZWPpdIjSHVDRSqW3P4/QC
MM/u4OjCvOf7vxbT/kr9d9QormdbUNJsS8y/0FI78OFw0DK7V/u9uoLxLdJKtAVt
5b2HleWHOoR27hcpSO3ogXFwrtqiRlZIVn8xqy5rxOjLA/3lyyYNMXWkj/dZ4mdF
eB1ZNhb4St7v+b+R5JdH+eObXR4hmNGm77tPvplRV5eK24J0kXY1BdGLCkarvMOv
02eXlWVWcPTGjG35+EeAhw3AvSABRCTkHTlXRYVfNXv4eL42+rnkCnZfkQNO+IZf
J2vKfH60vhwmFHFX4/eD034VEHZ7apv2wC8dY85zr5baoNsE3d/gMveEOrhLOot5
Qfyh9U7sngENhx1dunmfjbxasCcqh1Kcv/uH+2GYi61YWz3TqedmzzTwLwawWVhD
DO7hTRDi8AvnO0pZ6tJaNZo+OadZnXbbf3CMrFXFTif5ZfXHe/mShSAFI6uw7cdD
kLB09VrGonYyjQkaJ+zQnsCVisUZqc2/K3Q0h40mWDcyKI+k/Eux6jOTiVdmhwJ8
8FJyaHHltjn/abR5I8YPdbcw381euYT/eWyi2DEI63y8fHgEbnRQsfsb2O03OPeg
sdBb+r5/4BvijCtJz9HPbiJtiz0ArcrYAulEdM0zh9u1q1KxSZpKLwVX+5aRVXJ/
9CBoSKCd3Hv30yRBk0otpvGRYp+Q1AbfOZ/0khugIM3cNuyPSlVKD7pWVm6/3xex
EbSHC3MC6FN0WY7ZzHVy5sXz/nz4wWaB6robXn+R07SLdiAh2cFxBE4ZVdx9vB9l
edYb7K4jvkDrXQvO05FpKJ1DqIvTgsPvf79hAmk4TJNpRjTrNPFZkcrb4LaRa7N4
WiqC2Ry5Ej1f8VwFnHtBVi1pwGoxE41pFrBaCh6dRdQbnZjAWBWfmksGHa0r/TyM
tYCiYwvm3Rkj5m62qSeN10cNfWGW3lD47wfAXmuaPncVvBeltMszi/jATfy06v8u
1s53Yy9drt0apneg3DgajzvcOSwauul+hMtpXK/7wo6N7a2ucpYBD7x5+s6KjaNk
I+wHLcEPECOxJ9RdnHOvfWM3BZpCZKt4f+9KjcmAmaLNeFqsY60y1QgCryoZVL1T
ldNgM9mugqGyrncNcKaJwMEWjZuYWe51ZJx5SrH5WP4l/l2BYR0hWmcjhwAl/r+4
SFRpDtVujw7eHmI6c0iJizYSTtqyFZoXlXYst0AnPNj7akvjoQaZXXmo0koRNim6
jpAZtKCVTO8TdMIgxxmIT/pZl3It6oryQ7FBEV5mpLvgKgXzibfh8KenLl961jXC
HJZcTSSnoWle0INKu0jjeibVbTAegHcURjDEmVvr+LgfKuEV80SAUqFed3jSZTLB
LJsKJhecjgKETtGqHApUCXXbQkyb2G9oSsZHJzcFi5sbdLXMYZV2DG/DAovY8v4y
SXX62GLFMDp3kp605+CzDL9Zx83mHUTb/RofJsOlWhToovJlIarO3FxJ876V7KvD
tPcfDuOEGMzhBO+H0mXjypLZBbfm5xgRnk1C5emhkJWUy9sJXu0ET7iswJltDjmP
DWbW6mAWhBlQE3HClYmFYzyiTmstIiVaSVsIZQotPMHulvK6j9/KyCNGAKVOAf2q
/fZoMyb+OnEJM6d8Gmoumup9asYp0nUB4rFJvv7fdj/dcADKNLnTIC7dHa4d7vEH
kDjM+NM/TgNyCOUxvs9UPKNOMz3rgXKBPE6Yet+gLsHIUcNkeeZucUtDExPRC7c6
0qXe+JBZjUzz9e1agWP2GKZJR29Iwh32H45GbEUtl2ni+LM0C/xudTBuSSgfJjGA
/MAIeNsi99C2oRspgASdgG0ZlPbnpVEq7eotNq1SQl0iNDXgOT2+nVNoo53QzJNd
KLw4tb5ogHDNcgJ9w4Ncr13xV5NA0Skj2539e5xodTbGTmS4gG1K7Coj8TrnBTBR
QhmwTO3AZxBa2U6eO4gSPIUPdKH+kxhkv2QqSID29QWwtMBcUJzY06kSiWdFCe77
YLJMc6MsLSwjDVRkzQvSoCtA8r+RprEymcDFw1Eq/UmeSf0VlIPBv0Rs1gIciQks
+rypwRei3oA1uqJD2KtDhykFQjXfaLPe17ocrmd68dWkRpwbV4I+DS/c5U/AH4cW
za2gZO0hVTr4kK3xW2K3AZWmJyab73baHF7SWHiNzWfxJ7vbAsKVvgPaQ56lWvfG
pivQQZhIWwVhsKH2tQ9Uh7Ga9a1WSI1AkmrLZ2Mj+Fk+k5fr/AQmCzGU1kLfi+Dl
vBce1wq93XZgCUWyy60d+8ruzpmfBYx7dncOCYAmPfBwKlTazrfxcljmYrwiGW2D
VRyFdj6MHYubTZFz6swTAPmv2NzYCPOz/359vgJBdxoHHiRFDbpJoJuwu8MtYb0g
wYaGvl/GJGMdwwXjoCGVHx0u24S0mxuRynuFY8sI8GdyMbXSgAE9KuZQ1DK442Pj
MmSNjeUIdXaA7Gwj2MzX/fWLvn0KHFzU3zVwGFWXgeI8zrAE9HBeSWRBvRumY6Ea
yun87/JAro/P3/07Es+H0K5jcbvIDZ+zt/jWdSrWxaYq0t6EqZOs5HQ5ogWdyC0O
RKDa7R60TasNgrVjykT4ovFT3KI8wvfiHGipXEOJIf/mh0HuRw2pUKlRUTWK5wkp
3U7b4tKwjG99NeDK6XR18wDZZUUe4kgerMAE3diTWu/4aWuZvE+sFI0NkI8Aw614
fTL2Zc6BNFRy+I+ND8KAG9ssxsMGHX2coJDBzu/1Wo+4byltTHUylr6+Je1kUkMR
nXmwQ0QuLnBtXMbpwiPquShnponxO0mEkTlEAOtbmBSxpU6q1mpheKI5CUNb1Cv1
uPw+to43QD7qO1mVkJDV76r+wgdXCG6Ys4Vi5t2T2FYpyFbOhS9nSfxwo9QyRz7y
XhocE9GQibGO7ZQQ5RB/wSYMSTaOdI13QoY1NaKk9v2fBxb5PXq4kCdtQ0rlRqS+
kRnOpdzfuSi/Wyk/ZlKuveYxLJvorA9B6HdqNOjvEdvR6H7Gag81brxXqp9EJCmR
NjHpDY1WrDCfx2Jg7M16c/fviDN3JX4YlohUOA59jaAjXxV0Avsntr6a137goY5k
j6jY6LgseQs09WIR5exT2axnSDw5wucwHufqUH04HQFFnUzEJMwcPfox/QGBCYpU
hip3NpCEPxkV0bWfjxGyUf3Pm41gSfup0SEEuFKrJuE4qeBdRpudkUwVuQch8HFw
AzTFpqUInkd2QHpSvfOo0GBqk7iJHoP9xCouJq/FJRok4pec3y2LovqF+rfdK9+5
uG3LovyN8pWgAQD6bp6diIIuf3yfGx7GBgDzHKL/cEG61tk2dtrMZke0nBrUHpbu
3BegxNtLBzzoS8cWZ3s0lbZwhAuMod5zl9IuXSZLpsTDOajqR4vuu8L4CpVsMO51
zTYfgph5IahImJ0LSC6Vk6UqbiKL/Kc/2JgNhXGcmx6M1XOwhm8JcbFZ/bz5VSFG
u1XUXhK/tS0GMYbOOLmgBWenBDPMZCluAIMft3MFN9ur7Div/0FYAOrrNVv1WglP
FFA8Com/osMEVqYUoCaYk2QC1+8NoiVDie6kviUdzNWILzi97G9Lyb8N/8ocQHrk
M73UY83OiXXFxr8wEWAG2uoJrNSWqVWcKqpdlW3bgN3m/z6VqEN2MlCbzL9K990J
BkxPRItNK/91kLdtQOvsQC9Zr5LJvWvrU4F7czmjZJMUcETfFwVlj3acENe4mR9j
G+HpGhIRifj7FmW9Z8U43LFNUltjob7f7ao0rS8yur7URWz+h8u0GzJ6r/skVznA
k99nNr3C5kVqHJNtpWipZkv56cIyQH4mq8BREwPdLbOB8Ts62RCjKBiK+SSwYo+a
+95PKP5nVYqwrRx1OdNGs/22vu1OErM7SNNfoEnAFxv6j7Od4Q50BfUvpMO064U4
6MM/AEgskGAyt/dRGB87uGtJXfy1L64v4GfmqV48PKmOwNl1+0HngG0gNqDk0YA2
iAo5ZijVvq17G1o1uR3gEG0MWkRrOZ/RYnuZMGjoKgFMt7cfBft+A4Qxb1o4WV5Q
k00fZYadVdvHNU9BhfmMuk2kMIlC8lSBBbt7hla5Qto149roEJZg0tboQiW4KrzF
jkXOW0v7VjHEQhKN5S355WbWumfvkQY+GvVfyYaTB92UjuV0SIx7AGU0MSfa6xIj
XHWCxe+UzCZEQDbvTPSswCp9HTiJXyCsctpjoeiHicUi2AlpJC9vmUPaIH56UnoZ
v0Jw5Zn7GLHygWA2Id83nda3QuhGbmdR0HZDEFP2m0SLC0FR9vBK2gKFyvhfM5UT
uipXDEGqGZ//SILJ1OeEuPh8m+8IbSCxBZemjJJ7yz1AoOOLmUSMSa9PmLA58g5z
4f+QMt1p3Q6B+/kKZlL+AWeYqKJISdX/TCTp3NLWd/XTvcag0pFVQbPhJ1V75Vwh
4vskq/E/GFDt2JvNXX5a1ObIiDNUrcrkJdplQ5JHukfOjdfpg9DO4eCUQywv82X6
H8IpFsj9aPhFERF07u1YgZTMGXbY5OpAE5B9QrpA/9DTv6AtkGHd3Yp6F7/yUrDG
NwYK66xKU+hWN7EVkmqwuJ732PWJ9qxl/SUpSuANJlrQqhQMVSRvmDcXsY20NddC
YsFU0QePynIy7dyNgg6IjI8ihtQuU1CemrHeettM9oq0p4dOAU3zrPI6dMpBfpsE
+x+go8eFgyWIuR7UmbHUVZtGXx1uteFyOEF36F4AQpzfTYwwY1UWSGAqmdAQxfQm
VnSdF6yXbMpD3ooVDyWU8+M0IgDL6Yiyi08e/qe+bMbtZK+Tty/mU5qQ061S+hv7
mnF02l/DQjEH022bbXVL2dqb36fZaabCy3CDRXpyVHVdpAHYEPIYLK2FpCIzNXXg
u0/WWsYHZPaniDYqea97NplCb5C9Kkh0gmJIJ/g2p63OWofAGf3zJ33oSHDxzxFy
FSt3ice5ELvytdxD0JFEKTawnJCxCUVkb0qzo4qGlR/T+lW7P5vQHWvHsMEh3KuA
yYnx5XH0CORT+EngFmPP6HSO86D4YKhrtlBLsNspOZIHybOF7dPmIWfx3dtVfUoR
lTG6tCHosIGgptKXy1Ck9m2kxgrDIERPErTR960PLpvDenzhvarbNeG/vdCk6prR
D3w0dhQb7iGr2Rr7FGoYCcpNnNi2Kogx1DcPXvMz28RJLUHrpci64x+Ey+wevL10
y6GhkTkb1GTikwIr0igzbPrs+RPSX1z4ChUQW5qi7+wt73cSRmUfeXq+PcpvTdoh
57x9bdJOS8FxRaRmgr+TxBemPt/SwUb1hZI2iar1/KxHOD+GOnSKIf4dTkl0T5v+
+5n90G1e23/ghQVdZtm5c3WPCnqF2lefsVwOefFmxteUciE3A0/ej2IBwwh6SKXK
cisAuOTgIVCU8YJCjhnuQkOSqSEKV/p4sJs1WW+36k8XeF8dFXVnJX8QYjFvhZZV
mNHGfEENrZaodsRpoZamGsQm+kPzJRTTqEkbOub8jW9sO/sBR8qaussasUEeBRJN
FQ5kuhnh9AB6L2eN01DNWq9iCJAfIgbjwAOqbETt53fqmaaqPFMpTZcTHHfbP180
8LZZYrIGh6+7dM4NSLAc4DQmR/KNvl0pMDBZm3kZMhzktGyEuTFbo+y/RF20GWeG
PodnZ+RqNnswBseEeO8vG4mVMIf8R0q3m10AogmsjILbpXtHyQ8Yk3JN6euosMyL
d77/xlrfvQ2dQ3Uy6pe7M5g/Ru6vsreuywLxze9KTcFsGueOJlOthipdnCTh3zhT
g9K3whdyswUFK9DQ7494SVChqXmpMAsovmpeFQ2Bx927TMB6Eti0EI3WgCIwG60n
xTinudFW8X3Yrn5+oBFjMHb3UcPPQhD0J3PA/+14Mn+cofaKgW/ag6axX+tiRyDO
pKKPGOiyLa1GMtsoWrGoKjQkKmhDY1AROPcWnVm2i07gmphRTbAYARRBX6h+RFTI
xeyAXYYeW0lAoEzgkzR4gfX/+0mlK1GVvYZvKge+0y1iza0TBbhrSQ+h7VbJz2V5
4CIfNRMdT1BMvOgU290BGoB46LYw0gNNNrTrgH1QqSMJ14Pujb7db+GrMfxiVXVH
QRzPftrmGO69BFBmJbfdgZw4t9L1CnHp94tlEMNYlTTEHJHGOlwyfsb7rgg0EuBK
7N8YBfTyAbWZMkh3qE2UyGDvOkLknU2GFe+4sQ4quOEbXT2omQGsb+pCySnk8qPS
J25GC9MYnpPxosJaY8nCJlpRwFHVFKPiwRlTRl9G8OQUlHMRkt67kSRRiceUKXo4
eC6FeF5EGkqzPEspHXfwpo/wAVOGZ5LiHijmD5dAg7ORxRJus1Q3k/lDrLuInoBW
iIWTn4ApRrw5E2uwc6be7gUx+mFEFGpOLON9ILG2PQXuukg7RaCHoBeoMDYwah0w
rmdMX9OdC3uN+9+WNpv0t/NIa7RumVfrC3vcJgm6ClHXd7m3wjxGJ8blAvDmN1D8
01iDUuY1gFNdYDhsCTLSS3F/6IZitXSycKMd2VlqCKI+0i31wFV3HDxhKQM1m6oo
UJmoODXOd9VOWqGdka/5WxYIGWbEzP1UgVLaudi17Lf+mIZEihwSyFrx6boksezq
6WmN3ueEdgNrVBI+ggFITXT6bWlF0//OznvbPHsMrbucdgfPtHCCIF5Jhx8/6vYC
2vKlPr0P5sgNLM+XBYSei4IyE7xKifpeSaVjsA6COJw/rOzbgPqKCKd0oZsH+vE3
NpZkP+ika6AuzCJnO14d2mhIBL9dFKE9hHugjznYADX7LV5S3sa+YQg0xBGNZVNx
nad6aQSYxeZl+HTa8nUyGleQXPeWjPIjhYpavNCytt4phINMwv0FYoZYbK68YEpZ
yFU0ZgLNGxrduPf5GhZ0ZwwJuPTZtI0BcOnPg7WVVxUEO7tnULnMnsqGNRzlKr6A
lKWBaTDqOJq3JxM1t+U9OY/+7IGSbX3e6S5b/h6wEHaZbu8frA5gZGjhoqDOgkfK
5hF6nmvMi6/97upF9VXpRTHtt6GHc56Gprwh8dOLnfj2L18Bv2V7l5Kgga5u5TvX
esd58dXOuRHU3cVofQC1UmeHZjqs0V/N2fi8FUUe4gKYv5XCMTD4pZTcPRjO/k5F
7sBagMa1tVZNmblTMkSL8GNVULV8rBlk9p8kYl1EU6XPKFZ9bc+K1evLQir89eiH
GDkz+wdZ4yfDkQTWGzEQBkkVq1+hNtaHCmboQCeyR5wN+KhVryD+OS9CwL2ARaf2
6wM/E7ZsTQL1QCys+DlRX72s9NeAwEA2z8GGPuxMOyykn6UiE66XJBjqm5RITeMe
S+MowPJVxRcs9JzKub4hT6PEK1XN3XgAzT3dWVoceiiQtSxsZZr5BA44DLnfHXkm
ccm6Id+5Y92Rj5XOXmFCPZ8td3nivGj+z2Mb+JzbCoMJW0qTZ3I4xmJ0krNoRU68
exgwLKcpyg8OK3sWkujXyz6LpB2TJSGojuGvsptyhJ3xtCBcmioaUeWRC/9Ptty4
5LzetQ7xxahMo9PdiNWLn2r7rNeGR+40vkQPgsvUt0QFzeW/xWXiP75Wnq5QlVDG
qCad7kvgRa/rQsP+wbcFKzjMjPP/MzeLR5Z1iqzkGHt+CyHhUcwc0qiQgSYk7Jub
t5pnATg76HLxrSU6chNyrhq2xqaM94UkwhrG4WOiwHtZ5hTe+248S+9TxksskaBP
2HuSJP4+b5GJRd/hHt1k+WrLYzepFOyR2oaP592n4K7q7ILtv3QVonPQ07r3vn/F
D4pSgfjSBeja/0nNlFRAZJRykS247UgUDntrmOzJd6DLHRV9XrrREMVggTUpxVcN
4wtEb7bDznPWX+GbGZlS2HN5aFRarQ6jumJf51eRrl+gAfAaYogzTnMbiQprThW7
fs4Q034ycfbUXnUS0nsUD4o/FCliMrkXmYtXdBVeevgIOqxNG9IS434d9ltgxJSD
nz2Hj5EXMykzAloy6EummFbkfMMbhn829miXaHeQLb03HdRMsxOsMWmB/PFiEI7t
KF7lOo1LjOcGNWjKyxsLOPjS3kX6CIt+dmp+1cY7SS1u1GsXzVTgmG0dTJpwL8e5
I6wDQOFG3s6QTcX1WecAPre5D8fsCcaLNv7ER4Skcb8kzdR+j2VzMt2WZQjqRhsH
FqK35PmLMy6oPW7XH0zAhM6aX+FpiFSluk+/CvuGXLE2+DVloUvpWMPi6l6ih6Mi
qJC1ar2pj8CQ7OqGLhzOQGF3tvvnjSWUR0SuhY62CtYqAjnFg61EuzmDuX9zMvUG
NxeKzYPGTzeJz9Pf20BYWEsYl+mEyfpqfjwssEWey/zS6y0dejj2F6tANrMzTmZK
XAtUm0qlsKIo4ehKSXfLNhTTj70HLDjgPImxY1hXconDNNYycR1b+U8OKT52LDAk
Dmxfq/79hRuNtf1nwoRnLfsp8dNSZLO0hIikG1srvIm9xs75HyR0hdAtQisicptg
abpzP5pC+sokrQQfAvzA7m7cvKD9kuclgB5MFS1C9/clrMcG29cr2KxiiYsHoEdC
3Tuftcm8JXQh/zcL1p5cY2UP7lwk1tgzDBz7nEvhav+JUSXR7KCpizOYMefSjeow
hjjeYf2CtkIoWLKwBuhOGUsMvBhIbBWMTtffKsz51dB1tNv9ZSD4GCt/GEWkyu5e
TQCeAn4LMJulABzsijxctIqZxGGJ96sCqbg23kYEQvDDBG5jPe9til3w8lU5CCa0
tU967J0MNPw/0hSiYAIS8kbqzC+4rxOxHYZlwSCQ0Vo02QpbKVhxaP/VzT6jdl5C
Fh0jYT2oX7lRqbjt3JoEo6741u5lUWr7EetDvndSXsC9yfwStMi12nN5PQnLDF7e
z4vxBdigGFcAYKFOBVqFYdX/tXRHdBx9B+IsqXuQDmHAH8GKzPzZ/Nqj8iQhZ78H
UF6YDyGOGX6bUEtIfp2z2WZHPj4g7KVSs+8FWL8R5Jg6LwP6O+CIRJ8GcbRxtKVx
i931cjOGB8TAWyInJoyAuzu4BuDTZR6SSTRN3B1wNeCMNNjkh/9gY6R+44oasMFe
q9/qDWvQjUj3Re61FuSeeTOSD30rTkZzq1LhhB4f/GrUyCCQkUF03QlH8jjGBtdW
4mHvl2i4wazQCsqKwaHD7ZZ12i8kdvpF8Nlh6Tk/vf+2UUVKsqABfJjlBRF6zV2z
ah8gSdPdXigut0aJb3oEi//bVZIXWthd5sAXXQ8uYz9/xlaXqQ5gFAqsPpnlSsFU
sehLjFtze38wWYjjEuk+m4i4BDdf4ws8mSNWeVun8Ymi90ZplWERcTIJLMFg3hQ/
0g+JZUr2BI5wOdmaR4ule5CFThPfMgRTwtFfA3JzoR71UJyCCNa4LKqZepJOIcSl
+l3r0e29c9plbeN7fmjHVb0YfpeOWKy4gCC5oYaS4+p0byPsBIKLG2P3iqyYUXBA
6GPK6ZXVYnE3U0yK9GPkX5Ph6N8/WabATZmxRZ8LO75UzR+cc+k9yxfmGNypy14+
rCB6XOETsiLtorK07P6SjBQVPET1n0BQnMT3nstNFJLn1YeJTYyhPeaXBa5OOzKM
eVOfXOeQca6q9E0syu4/6K71oebIbT0iXbzWph1O4rSgnWjFe5bJCYEs2fwI5VGc
oYh6X8WzmbjVZRdCVAiew8knPiU/nd7eOwyWTZGDsss1ylTsZFzWuD2qT/SE9Pfm
xwxnY7S0o+bRcT0oMDPuO2baMXY8nEHQb9l6zWP5p1KeXgUuvlIOcFOd5Yhg6j1j
btF08Ptr1TTsDPRNXRwx+IQ9jBkgQOUTRJxdHIbcfmm7YF42RdXy0mnErqt8YOTg
PyEHBst6LtJC9Ubndl+hBD0BnLTV6Ksmy+0ycBG1LEavnR/9/CfeJxs0RHrmVC4p
eiOxrYTf1yOLypQQSoTgmEb/CNqtN1FSDFGo6+RgcXgDNIX11NB1MN5fNrpvv4AP
EW8F6YuucMpFQtSdgMOa4bBuoRsQQQgNHfVQkbpYXDWRezDzjxPuAlM8E8bFa/TQ
vAaS1Gg2ceAnFQjAL2ONJSUsBhEArwQidOWmo4r8MnbfqWty3N1V5FMHLHLqcmIm
D0ZMn4nYH2PSvjIMI+y7PJyf8l545+Rd1gb9EcidDlsXioDL5PQFntH6nMnFpWOX
ZqIiN3e1VHRJHBMz6WuMZzrND4udahf3ATwjjtTuWyZl/eTMOD2K4TbNvLqhIejk
a4rsJBz/xiirIv0YDcSuCUJHfoekoXoeqczBBrugYJIWvAi+Ly/NDVUbV1WkCjsg
lQY7Fh3z+r17sy+RVjRANeXQdHD+WMHwCoOrvxs1/7gXcmvQ2GpQWODtIll+4Sf0
Co4YP3Hta1WMFEEXfUh1dp7UBX2gzuxxcC72Zh3tuPywByC5affAOVu4o76xVrQh
+eu8gT39UU/3iWMfshwLlA1+KduhsCbZYbOrvc73M9f6Yz9Iiy4Q24e68w/KTY04
4GziUtUozxbb4l1FMTFMfGMqPsJlTbtJpVx/13yoWucpwLEQdJjBKzYzD7Q6tJZ/
LXxkTeziv98p6LA962Ud6N9OFxYcpMAbWmExSHVQCpPzDyv45YfaSlYjdD82d4eI
7EBxUQEmgseIrrJnzIe1SVV+YOKVwyX66UU71QZXw/ITnSyhX9kxX8U8nC7Icru0
VV2wLwC9aPWL2hM9/w1m3KwByL9YuRRthdqLsv7mMpwVHVe+V/kGL7TEIn3Mtzrj
W1vuULrneP89ERxLxTtFBsI8P/DN+fhjl+kU9jIp7qp9eXQw2drznuzJl1iAUfCq
O0rjUlEYoAFZlSvd4/nlzQjqzj53Es68CUgk68GxENqiejvyWSiSMwN1Dn4uUunK
rJvZqWflEPlXwLFMLnsX0/aZsjmFNqSzfWcWuySQEYFR1qY4AAuUF5jQwtK4GtOo
ww9JgvGVuf4sHJ7lwlAE0Q7BiI7HPTbPK8yrBmnVftS6qLbOWyoRY/LKksnoLd8b
7JoCXOZhsLEXYGQeo7AJZ973gShHe5SMUQx7Q3EtLQML1m29RfMKzziHabzhPAkr
RaqcKtyz+HH4RVGqKPYeaRakpiCnMVQAfgF0ZRjsijkSVRNLTAHdvrkAlm9TW2ZP
eGnfYiq1f+jd1o4BSamqBbWy1uENsoSR+JP6cMlr9q4gGZZ0Qd834iEV6et30jwu
ysArk0xe5h7f3uRLikpuabLRbNmYMSCQfH/nhQhpOP7pz9uNKfnf8nG8+wB/xD5s
CE7Bu7ka+IZn9Yv8zt5Z+OZlnhmeyBtEC6Byw2dTAHkCRWef3zWTejPaxSlQ3EOx
0/Vpd4y9BUar84sce09eh3zRAHgn3MGVecHpmaDGpUr/oHWmDT5mD7bzoWOZVjVz
AIsBhAG8VwV+TRrvO35xqS3mQ3ofapz6iEHRx4eLyo9r/aDLMGSKZlOnTKHqPF82
Xhotm8Ccb5N9Ksv0c7ktHTAK8Ha0K5LnSVEj6DKgqtP7aNH/NV4j7pSSsOzHFc3y
sP2YTktzB4GC2ca9AbEbn1PgJvtH4tXQMzLhANIEej/fdcvAExDfimwVoWDXxitA
0I4rBiBxv+GRJVdnvGl107tdbEbYmrEXdS8W4ebAOJ/E1g4txLXJNv40uHomOdPy
KhtLlM26GnWEtL4BmWD5UTzVKCgf0NakNcSxHa9vDKdSczMoxUxqKZkzwxJtCk3m
074hmks7UI3mYwmpOeXfWlvySvTohuYC1jrapvrAt78+xwJjXHaw5WhHsH5Cx14Q
vSS4xLsgAQf944V/lCEJTrs92LXGfEBh+7Q81EjPTvpAEg2vLpSNq+EVHE6qId8T
YrHYXwk6hLCZ8rb/ar7UNQHd54KV+mgW9od9FfhaAn6Yv5AGaBwodvQyy7BuvSJU
hV0hBw2i/PmsBoQT+YjdELaVEBRrsOKgRF9CdHOj4ZAQ2icQpfRQW70Qkp/oI2yv
ZnEDBytG34ixsBtt4auZn4L19H8Pdl7cKarGjkxwQ4qUri81m3bsJTR+kRQEZyfv
G3RkFGFqNuAH+xU++DV4OqF5D5rU/v9CXQHti4WM12n1L6vpWqPbflvBpuP64zl5
YnyY1LLIC/keuUbG1rLd8WRgJudKIc6d4x/y5AS7xx2ZzMZUQ+IljMSzsL9hRCxd
WdtdlceS3NBIc61059CVzrVDKI0PBlVli8WM/VxC9pgjj0sIprTVzraRPzJ+oLXh
r6ZCg7o8NHW+guAFwLzQAN2dybIL+OuoXeEKHNaZIiS0vBXri1lmnhpIEkp6IWBW
9DnjX1vzcMzUuEnU6gZiVdPQEH/vxEhiJSB7bNutlHkJaZPG3WO/MHQ9Tng4tSQn
3LNs3fvS5CwyE265yK7fslUHXzh2Due3ZfPSSUKO0IJ8U+J9/HqvkeGiWJUz/6Sq
mXftrLi8RId89t6JPRFcZFz82d+DvO5IDPoyqYkiRDZ7D8HxvQKoAZY1yxOV6H60
ceM8jiIVE9ScDlB+JdwVwcz3D4RPuYS5uvvpi9WV29kjicHhZ6/fFceaSselmOSC
Kbxh/kpddaIwWzGXHJ7Am+EzYt8uJZ5uxbdhoaW8+YfFiZkGWtp52kOsLTT97m8K
Jj+PZlICwW8PdAx4si8nxihR3uRoF9VRgFEVUWjeWzE+rLqlN0o+4KdKdWLSXH/N
N9flBGU6gAU9tcG50G9NSGNOQHajMm3ppWHMOA5fMKSZ7mYOYnaZYK8PSNA8YRln
hfPXxWk9Q9tt8n79gl/WLyn8cyeXaj3qmm/gT8kDzUwMk6u1jtfmFlFWbrm49JW3
j96P5Wje8Nq/uI0C4EinEDWDBpO5SJ76DmJyL71Dyl9bt974DBg5VA9ZkrUMzPbu
hKbelgp9RPJtgV+Qoo5gW4DO8bPjKBUK34DeLdg+301EprVEgQ1agxeeobpdRAto
lu+4hDhOOvkHoZCcLpktD+apx5CuNBGeBINDIhtr3N6bH3n85KSDQjFPajfodZI6
wTf8xZ8zrp2R+qwcRGBh8jjLGgSAtfn7TFRO4182Z10zPx+wferLzuIdTywvdSc7
5QzL+tPRKnndjcEeUt6OqvhI4TVLRZi4qXrAMYaLh0gFUS1kpY2nYNbCj9mbxTP+
WTzoas4OU9rUH5hpUlFkIs7TlG+mPFFEL+sabSpU21NjUS83uVO39vGpIurPlz0y
GES2AOywPA5ixdx3s3f1+t58mvbaCW8bxQzHRfyPP5GVGJsMDcCUQw7hjW2AKItV
GVKyXiXNT4KREXFXJ4M/1nbCXDk9plc1xg3vVuQGaZ9kdYbcpFPMDrmGbayl3NmD
iepoiuHEHS3Pf7jcA/M/1MbRdclnj1v1BDc+n5cTZPLIPiHzazouQ1BO6jx2ZAgp
8+n4FJpJ+ga8a8U38NML0eM56oVZYyI+gQ+Oa3xbHDkSW+WmHdj8VCL4AuWgkbu2
aSX80mfLqEnpax6MCsfrEjXgqKe5vt58PAJAhXHm+kPYWqReqTU0/5ppsJL+dSGS
hHr5DcRTeu3vHUY/rTJGGoXhgD47zYkwt0B/AWfVYmsXcsv8Zr7yOrT9MLU0j3EM
wLp8qqZmUNAJv+/vlgsIrcrQu4w7C3u/YMXSXbkmnHkcZR6dqGxU5HKcktv4pE+K
guGtX5JInlwY6ABcNXO62oAIt3EwnrBOxAfKzQw9RqzhzgUDkKcjLzAqWlNCGupS
r4HqmRjssgC5o2/izo6M2iYdmZLa+45DYuuG/MorGZh8qFl9su2t5CyiRf24pCMU
/oRAmYPApayWJoc9zzkVdA3vETpJ3aXutqAjkubPtG0DPgO3sRTBlervxt6XyOQI
CgvrYkkK8zuUrdbR5dZyrDBq6Xiu6AwN24v0Dk3oEnN9oCayI5m08tWT1jRK5cAe
r3gOgY/5HtdR1i9f0Riva/Db+mh0oDJ2DexmqsQT7vFcZcoioy3gan0K1zvJHzLr
zoiI2RGFnjCfsfOsS/EgdRepSB7OxQSDR6K5ZGZ16qaiGR8AgD6sOQrHec0ppBze
s7bwL7xGoNSlUl+Dk6TnwPITLYpD7ZMMSotDkI9qt2+ZCdHBHtTIi+I2A3+AI2Xv
mUE6VoNrt5IsS80OXMDlWFU+6a5jdy5MqHkAv/hCoRxbxguVhHQvYk7ravsVwyyX
b+xhfApmcH2kSu2lnprE8agDUqZWxueEDfRnu3OiO86qY0Tbohl9Fnz8YulcnIMt
ykE6XcDBqOy+eZXEYVdYrAcZq/TIr46Gc1lEQl1VHAyrkZk6T4fG07mf4MN0Ux1c
JPlORvpO1h9JU5xlhB2cbc4iNA8fk1AuG7nh73xFxABIPZAxTBvEJCGIXMYhp/9p
yOyM2Hk2It/86MQU2txEW+TIDGTvKHPjDAdHP6oWWQGT3QU5PDUOQ6XHTRd6KcrU
wSbrwNK6HWDmV7/nWUB/ggRUrCp8XtI8lBns3tEfZt1QJ9hhZpdmvs/TP6mfw0Ew
JfFSlkcSukPpBuXN8rr3404hD0wLNQtKrcmFCWRY0qD+38bFn6+5gKxyzF7A4JAA
fSSmG0oHbPrCbLXQYqLuRYf5nOqXK2uX6Hj8W4DtDK9xa5FcdlNnfM2LPHz4ZvwM
b0Rpi277KsK+ALvgPvYyqc7fWraAo/NNsMZ5PURowjJor49d+1HgT0IK+5niiWpx
0U4HbGzXlLJ2LTcWLXxWkQZe8DgeBhq3nlQeo/jwpFcKHLKlkrjVx56vXnmyl/Kh
bFAM3eeLLtnVMY/phaFrSTZ1M+l/TDV/zPlkADQGTu+z73vY1XGQmRD91Ht8aSAg
NHFtwG2gVbnZ5p0wrDO8qd7z3tvvAXjeS7nWv4BLta+01ycdLDzi1Bxetq5GKLlW
UCY6zctIAsVRpHWqyJ3dQmDI3WxnTF/QFP2+iHiLFYgDp9UObzwY9EYye2zlOUl6
RUyjJtXCch/GhbHu+nQbODFVu+0dCItl3Q7y2vIPbPZmWDGwocQxDtD09IiE6yzx
hUNXHfN8I0TOmK7VG7t5s1EvZU8QAyOdaus3FOgrO0+Oaw2ke8lvxLgjkk1ALeCD
LTH/c6faCWWkk2hiEPE2GJTCaeNcZdk9U1HqtotZJtsARXXil1AMtX5QhVnT2sEZ
vU3gO72HLaMOdk5qY0jcZQjm8mpt/6flt7Z54bBodOdn8B/1XQS1nRDk0GE0yRr2
XcV+uhAuG9H13Ob5zzm30TjJqvcaCiu64Rd7tcOdoX84iuJHck84VyZWooz63xh+
apI1cisD48LTVoRp8lXwaB433JRhmY9g6k8eWdqx1sLU81Z/X+DW0nmvnXaZLIZ3
MOAKlig4Od12SHnuPuIDTBRqWeGsJsvGgz/k+vvA0HavbhRVz4q5s4LB04ra1/U8
pzwWWvY1HIzH9vEzg+x6hx1nF3wsfge7dStpLmnWQI81zn6jrcHKoH5GJSTO5gTR
PJz6vv+q4K2EUortpFBWGSOkJEd46Umk6/0gowKDkguI97RaFJSuAW+ttxJX7YyT
Pvc7E+cCUlW09k7LTPqk5586JnSc5wgM7b6er/K7vWwIXBN/WJo8GmeezCbKLSzL
xNLWYgsNm63xiLKiQ8iE7qkHaQvIBdEHlUQ2S9rQV+ocnlBAx1Gnv5UBIlC9zEef
pADWrFD6gDp5lFGn2Zhf5xber8rIhH4T4ieDe1Q25brWlA+dD1QHagUhm7D1wCZX
cUya/+M/53aWTvy0bv5gXbNYEtUqtG+hY8npsQ2hmQQxsbEGhFFTD2TzzOjmwtP0
pYljN2Bb25TvQzFJMUvbzeBZ4lQG+50QtVadAdB7cfllmRW7kJbK67NFb3WFDK+B
6dPNWbggH44L9n8KX0vD0GBEskyQziYRqYHyno3fGSOGEisu6o/bCoDMgu/XgKyy
UYsj0LNCqvlVUnCVYmcuQrndrLr5lG4NrpE9irOhCllc2MpewceBjxmzhnd2Br8i
8txTTj500dUgKxpHDYNZNdLoCkfTRidmeb7qNg2PAd0A2lKnleEYpFR6rN+puB4P
E/T/T19qzjAuQsL3aBp28qUJ0dYj50VsSN3LcCQeKQ1WLLQZKSKAHAt83ls4nEnE
5rDMLExuGTIXU57d0wey1JPD6QIXraFaLz7fylNTmGJNopkY+DPOMceTAre8o3Ei
l6S0xhWBfQNGr97qoDOb5LCFqdm+/XCYCdgP5m631TlYDficVOuiQ/vJpRQZZqe4
qwD1x+7Dktqzys/yqT9Fr1410QnuxYakyvPaYQG7dVhy/VFPVvUguuzrft6RUL/R
opbZabxOYuqbbfVXkwbgFHqIqDjPObV0pWLWDYiCP3opGcY8oUMtMPrJSlsMgeBx
JT8NXzsg7/lwYX2XyK07B71Z6aEJPsJ1hinmyXqgfRFuhb8SA2Pwpb2t0lmFSqIE
G8TpxE19obowc/bqQ1e6TQbS7MdEoQe5I5P90M4ekHgmXHdlj/JfnBj1XLwHO9QN
QLWktXh//AeU+qLWp6nogkzFZEtD+8nQkzgBOxRNoXDh/fg6ynysrqBld4lS4d6i
ix3WB5F74iwMbpRjJv6+zUvfb9xCyZG4Nnk0Uk0YTuAWGyW9Yvr+mYqU+Z4ZhtCM
S8+j0Rwuty7TJuT+r9nJFcrIOrb9gCwvHwI/LbUMkbJwGM/I5onJ8581zrbbyl/a
MFNC7+3RZ3SiK3u4EKr+2wjH62xObqMoQJmO05G5X1b8R8BrZSKyLzvqu3oivjvg
C+pfTLzOrubwOam8TQn6nwiisfV582CiUW/1ZyZi/Y+FYTf/iDSLVDNyjPCYsGg+
VPc0zU4zKoUc9EKSWDlD8KRYbbxH8p6JtTvruqG2G2rdWfWtqTwxXGGbWDNasJb1
i0pdegsI+LIpM0ZGCGzdkJRCsZAAmo1FZ7BHuqwCU1Y1I5i33bHAMNVxPsao+Pf9
0wnR2URi4QVurIhKhLBV23JE2lYXPri2K4/wrOOiJ1KyT6BTQGsYnV6/VhJ9TSol
5EU6cKW6Rno+ubW5jz+/ioUfWbSqr0QLuY4Q8A+9BQsQnTslGTpvX6BuR/FpioWo
PUqbm00ACZjS1794Evgu4DelOqm9ilexDcLFGi4xONr2pAaLAjJRKrRyJv3oxNua
9ssm+ua6Lnif40vDb9D7hVR3Y6rpSTGqBeAPvoLmrCSGugVedUtFnSP/hTgoacXq
qoBq9BlAzvf2CbXwxsLd2lO7f5WJr52NmdR4bOVYPSvgtvNQais7OPghx4ln4G5h
VkMaPfVQDZXIqWw8MSjb5rB8EkZfnR7moDQ1tZVA2o34raR8gvKYEQT3TMUrs2Ma
khZ2O36x1BJruxPF1ZQcflproP+QwY9kxyatcaQ3y0ToOUk3WW6q5W8VxEZ2IW/+
qnq0nRAJEdk0gPQmE01iZjAxZkoO1/AygO526wH+9BrwUjRzgctRMxW0wN/c7CuS
35FdJqJEmo1r10LiMNyr+FKA2drKlfuOcK7novQwRCdd3DYFbpGCFUl7ehzU/hdq
gXlSuyDkoDgvGoWuXn8x0Xyv11psWLFN0tE1YMyDt5nVDj2AidScrV1+kFBTvUey
H5uCJWVAA3AKl8s2nY7HNrkTCthxqZbI81pUjVxNL0WTdeZiy2pOR3+DvSmKt5p0
KUlzFhfN6fSt8USmq0CQVaHDIQVAuFV35NVj8/yLuoH424azwEG3NEkSJLUfYpeR
6Ayr3O6eT2Zik8lURft83K5D3ivrTv1BfrNMBonK2vF1pr9sAmQjjL0//0VM2N9/
hwCaBhFIzMPyhaytbUHNaLaCUx0ZRyziFoFgh3IGtc0vRHee1gfG16GGXPE3dH9g
YwNWWfI0phjfp2Sek1l84gnCjfsSz/mGjT5sT3YUA5QmRg7CgOn7RjMvw4BRqibl
MkKXhlDeTDZ3LMJSBb2fdZDWB3Ttne+yRa+k7GGtxCvcUbmp+q2Yv/x8ayTBxdUj
AO0wIBsuvvtGB+wAgN+f85tlq14Cbxxw8C2zZAyqpSO7ChL0SReGda1NyoD8wm/y
bmCGG9FH9xxhDUSv2B9CoanFnhFmemMe4BM/nnSgPfWaA56rEgdUgQVfOn3bYjBF
0FSRb1Uq0m1AMm3fCsWpi/iJwU9wT/hpm2piYjClv5+GJpLtwTuaNh5ACHDhZAkW
lP3JUkSlC6l3S+z/vlW8BXgq7SP+NeEsdKJBCbIef4xpWZR4mzelZ37J3Ahl399l
8E+2R58ZE8mB/YioxyQHpaMRL20h7897UYr6TchSHgsD01f0dthB/tK+wFm6GhXt
/ylYN6oUaptQ6dZUm+vNMPhk8XNKqWBc0CLOrDodUkA9WD3Rr+ZiYMAlvZtUm1vv
QmEZIM+GPkIKFQOpy99G02btOy876aTop1leGcdc2xdKub6j02bFtFonAZphvcPm
dib/vrFsf0R5KgVe4ZgZKkcNebzU6fNLIDW2yMaKQe+nQ7LR1fpZcgpaVLbvPgrX
K0tMMaYVT7+iylIyDvWrFOUFQ/7A7pKtlfH/DSdnBtUnt8NgZF1GtnWZNy9i3nks
cTXSC+HQ4YN3tXq2mAxGwWELx+g1VWPh42m5Hvhr5RPuVUHTlLGMHZKxNn2q7t69
aWPWA7OYZcUMmHyLKSbUh9NplqL+D4NXw9TKHZFaLlfB1Z6Fd7C7ZDvEUemWjJsz
QhBLTNf5PKh4EhsG+kFVxYcJ912+YcTeUM00Ak4tAhAfhMKlTk1BIBfodylLEYk/
9Lp8oUxXnq2g5A7rE8jsu2PLNv32MzWfX0V1STIzIt5cxLVWQ/WSKeAi0GqOTB64
OGSkiPd5lZj4Krke9YszCypBxF2JleAsCO69XH7+fLRVpdQBvV54evfbyvlF5m70
7ThbXfj943bn6AVrkpqzzYaFUwhNQrYqH1MPupCGM6KEY95MV9tte92iRL0/lLl1
qs7wWvJcU5W6UC/iBXDKFxyoqqSRWOICrVYdtfqEW0oNy9zdF8zEwEJA7A2kDJ7c
4Uip5vL+E3b4a30c7n9XrB1IXDjRfIJ1zpTYaCpUr2b4kI4OZFOq8z8fIEavEV/d
yh9HEplN3fKMbe/r0XcLB5ZrP63QRFul07KWEta7geJK/FYSr/uCZVR2yzicQ6yg
E6B/AgnsXmwIHFeHzskeJHKkkop4KR4217ir/f14EDRjY894VHuYhZBVx6tVYOVl
7Y7ta7YM9XU5dNgy8T43VpcXiWkhm4KIatfvZ+HZV8GiUqY+Re/DJ/tt8VWf2Mbc
ct7rNecie4TFiJkB9gK/82FVQSIX7+dJUUfzlIoVpQzQRQxN/3GnrC8uZy57v/N2
figwrSytXGKWh/pfMSIG2l4h+KDjaYitojBHG8HcQJX+ql7cLZVPcDlsPZ+Zcg2q
L+iO5hO0LDRhWB7jhofopeCWitBvI2+9e33Fff1gy8O5lBrazKrYrDaCLMU1ghJ/
l9uAPlsrx7zd06MGRbWuSH+bgNaCpmx51P4wemF14pEq6v4Bb8ZEk9As8mU1L6Ha
mP1j7Y8+Nwu8hmxF99RzTqAHdRIQHnj5qRtj1gV0/s2myIhi17gyI+gFskeQuQ6z
TZYI6GGXdDJapKAjnwS+I/T2B9qtdXqcOKkR2tNmE+0xx1cCGgXHgZdUM4h/XoJu
Jf8abOOssbqD2Jqg6e2hJVK0FFOBOD9WIfqiFVLG67X6zwDeLKtLIGXOA6tgjpsa
T8EjEetfL/moBT2WbC6m60W0tK4CP20x4HvHNZQlwPBsJ6vFgrqWuTSYsBk6PKqV
0MegsMDrr8cCv8xFAIhnru4Gh4kGWWUH8ypp+ADKMPE3oz1lU0E268k+CbLkzLCE
4HRjIEJ3njmk3cVpQpMMvSzlBlPeqZzlJcGdrT/wRopeEA5W/Gfj97CSI2VLKAqP
SReJZpC7vVFR8IBW8rvfM6pl05zUnkCFYKdXUZYSzKJcrS4OgPXgjF/j4hL6C4rl
bv5k4iE1l1l6xUlhM2sGBUUiGRlPHzlwOXQJhr8Xr0qzjYGmNAe0Qb32UC86KtZM
A+a2RRjGmFxiiA/Ydv/Lc33CbMoF6ECRebice18h4bDKebJufk14Kny9WRbbMu8f
XO29UVW8ducmVxfy6AE29o4rENErjIAPRqPLQ4WkTNscTEgMLfhI8vfOSn9UMuwE
+57aJJ0bnQISE0ZIApBbtzi3LMPSi/bMhfNIq/5gWo3aAD/Deeg8c6Z4jI5RkRls
hwagNKWTM8C2ByDWkENxqO45tG0WzVwLF9w0VoMrXKg/lr2+PJOFNE26LQDG64N0
H6WWAGZFluSRNSIeAOp2Rmq1bk9eB9atTpYGrcrdIUbM4xAjvSvY39bgwXOCjLL+
nS+fYF+HbnyzHdgytTI1gZje56evADd0pAv3Dj6sQxBkKX7RRdArS5CG8BqtY5qC
iw0XT1ZeClurIWUnKmfFO2p/Q8K25uwuVWuj4U51zfpaUsmNYRoR4oUde/f3G3h3
bYBdJDMn1PxG6zdryMps/x9tRyTSuAGjEfQyJd2UpfJnzDeLe5tSHNVZCiqTU2mf
oFfx6YEZFelIhMu9iUw8XoK6Y8U6x0gmWxWwAfwRAOIUVy0A4LC8p895qpPIJiyN
Kpx7GdQdOyH9GyDu3Gz7b310XU0F6bXmoKhgbYAL4YJK52R+ZtcA/JLwWhdL0FMr
THvSrWn84BqyAKoU61L9dxucL76REuNPDNoaMvEJQ4K5a+W9U2dpDRJgR7K2e/gE
7t9O+LSVg6YCpfnnVJpsy9/CE4yLqSnBWXisLGU3QwWhg1ynwzlZstJdBxQzAFEu
Ih/c1Ff74Q2mfYebPRSkc0shMt2kuiBf4gzhSwmxHPpHd5cz9rZSN2FPSH83w9PC
pDLuPFzKSzOc92X3wmy+rlgUCUUd5+2WxmGdae3xJYaZ6ysfIGVUD366tUvIpvp7
mQ1xPAwft4FQYsEwG3R7d+nszoC3NNUeDueQBMvIHEpiR3buLU93vA1LyFSxCJ9B
IZfds16Zwf+YNZpcZDdqNWW4u8hDwi0jOe6quIwKBP5SfzsYAQVPk4dET2oJog+B
Snacd0C6oQkRm1qFpxNRaSbVqfl+teK2Zg1ePwT7wUmDKcsWYFb+AmvATk50Pcr/
GGy0SDwgl31qYVL+dAROeqLOi2CZaT5jvGDjDDZdeR9lkH20yrVBWF6jL8SEo4II
MnJC/zb2/UHNP1EHp0aAYC2QNJi3TGhRmh07wKwGzHrh1na9emIrftqY3MHJBmXc
XwQEtODshlqLG/AflZWo4zJ6AU3OUGmx9jSA547+cxdRFM0RWrJYneIHHMUC5QKX
pzd/seyXRc5kyTvvH814jwgG/eXlUgSwW0V3/CBmuWWBUsfLGHEqzxdtqz0wEBkD
SAoWp/FICzDNutnzI2FJJ2BnRjHwYa1faepGmgnSbz2dHiLveIsxuH9CMLdkcT+2
pi6nDX+w6fnhWWS5IbwWuQsvq9eHIXgfIxGJuEH+7XeJiDw5jDzZ8WtQmYI7Ixfh
kSg9IT96S80moHPhBbpd8Kf5SWJN7ph+YU43v+V/XHm7EPxMlsS4kL8rYuN1kgOx
FLnrqJ/YsANrE3jhYuQaH/UixqXvX1flrpa6GSiYFwWWcgKivzz4Nyb9u9/WUAmf
1Hpf9P2X25qSMjaarbUVWU7P5UvqxMEOaWIP+Y6jPlShPd+drDD56btmqOM0MXrJ
PNvCisIlAlyGsrHfumCxU/KZ9MItSVbI+vpuTokQ9lYhqIsLRAzyWxPwHxC1t1Vn
0ZoaatYQiJPBDLHoAMpI2KBV95VC2s6HYN33VIuUI5MRPXAtar3ne/Vzpgm9prY2
jDY8P8r2Hux//iHfm54FGtmzubyxr0SHikImKAhGdtHKhJyPejZdgN4koSRnv9lN
uVO9YkSWIzvOxDhkE0PUjJS1jnNndBEWQcWjLaXpfWf5bt5jTBi3a04+CHB5XarQ
+JN2lITw5KozMX4kZ+qEih32gGGPchA4bUTsAVkyxAqanxRRlYcIqCX0xlEKk3lc
5FSLglNwhzhaTvU8mjbWuINkkLJ5yHP/BOZ1h/oIQVV0IvvjIC5XSk0fzGmyhM4m
Sf4FyrDBXqZ0owf2/k6xg2kTIcXFHxN1am/W1v+Ef7RTrmvLl77Ojr1+ls0Wl4XF
ftD7cAD2v2YEbpMbG6tL807ESeUxB0OdxPNRRXokBg1qc5SKXkjDMaOg4D+eT0Jj
kfky/MjUs06OZOROoE5XwLnUilN6pjY3SnlkDGFVdj8wvH+YSrDUIowdfc3MxRIL
Mig7zIuerAQaLgRZoZ4HLVzbmmoOy9iamzehn77lFH30pJpRuffUk+Si+EsDTp8I
jvLHts9bI8Kb/d5Ve+GdyxPsXqUvAuIGc44m04I6r8YdjazbBsa8Nzead0Xi8m7c
3Yym2V/RwQAOH/ectMABrfDv3CEn3UUpgKIIzHWltHjcsGlea6FZ/0qul7fzZcmR
JYgeABtY8TucN/jErcheRQ6sUjgqTAC2ct7iH3LysZk0Ef5tWoApkscmkMT1uM62
CfYEI4yQwhcJw/2scCwCM6HOfp1q9jHnXrxIrh1bCGzYA5O+2DHP2OMluuROni+8
ePz4vgtJGLgSyvBGlduH5ned3qrhLwVznb9Oj3jlTwVbgjjVPussKKxrn1DXlofb
yu4/1By/PUOEWDWnXxAaFE7XVFFe2JZnh+IUSgfOZ4duuUxx8ANaV+CmBagV5P5j
TVo0awt3PHFQDz2KxIqhyrWzQxYj4njksva2ip4feSjwRBUwkOvke3SGIaOWOdh8
7IF4Wq/+FeClAWSyjLO/uQ+DnC4+iO0j08LaspsfO54nImqiLqQOD48LpYrSXp+c
2GpjEsidGAljQxkTuFe3QTqFAKRFvlpeEjn6C1j8dWLSA4s5+qSGr7OrNajS5hMV
Or58ULdZG9wfgJ+rwvLLJCIqxZF6R/aXsMwlN7q0fT4TMaS7TQzoNn2o5fuFpwXI
fEH5gwAfe1Bc6BohwHu56Pvlh61uxX/6aAqnhkhOmQVIhT9r/8ua5gP/DVROg529
+wabdCJsbCwej69v6FuAe5RSkUWPaq+16GpcvPbjDSed/KUcl6GevdfSX9F1jYA7
hrr1IeIUtFBWV6W1k9iQ84W7xB5bE8Ej8JVIoCGGp8nw7MTTGm9HzpowgN+e3kSH
jW/NtxPiHAjM7Dt7oIVCgEUKFg+Zi5TdOxm29hIlonHUzkKb9sZx2BNM9I62a/Ig
z9PUbXvSktFamLPpLK3BAmMIV/yNtSbFkBKzuZjooF5iGlTmZI29XTl4x4oInN0T
Uu9KWdc+e9gS7vclxXW8Z6+ZNdTNOwmrtcy9yHMSzvmkRHS7rCb6cLFPR1y1PYnV
DNQUjzw0KCQ6Xe98DaQAG6w0n3Ck6e7wFzV/oEViPJM0h8ch9NEqhCNP8p8oDcgY
3E0FXoB5c0clXu/ln3vP0kSIt2DloAAEjJbDVqkENOMd0m+U8oMgIaMJk5I+vcQj
h5WlZmZ+D+Cu7/+njmW1mkDVLY58gmLnjdhvjw8aIJlK8596d+G9lTEYyHHVXLpl
H4fK86TzMMNDgxvb988BDvFfSmJ5A/6dVYd56Yt55ayZYblFKP1hH0Zs0uejng/A
xwgjOv9c9kETvFp6H8ZBIups12YkYFnQr1jrAPp+EEGyL4WVZZ7Q9t+ka6Y/QSMw
sA1qG9j5oEPNKy8s1qZHFi149cw6aian9oiAmJiXJZpb12kz9tQNje96GZwUS/Hj
rbbUfXOaRm4cBU2pnLeZOaQ/h35fQHYLaXCXPUcD69xdOIajiLx1PP01rZT8y1yc
5e9Xs1VeV9ljxoiHrJzP3rOftQ0IV5v5QoXpTAyZ4uySRNFPOsz141mpNstnIeCX
ImEGF8jt4H4aV1lmMznJWNMORCVl1bbU9kGDugXMmZcll6E05B4lSijz4wNwC8WX
W5wRCV/lq0Wr0WWYLhYwUB00W+mCD2gF0hnl6hbxd9JEaOnlGw8OSveTou/CdQHB
Sl8ZeZgsEqOTHg3C6r5ltKSOxmW5nipCzHHFHMEBy4Z2z7UExspX2hs8lzg50nDV
PHcZmuuoTTGRJgtXa0xikMuTh5iEUVmRh8JgcHeV/S7yuVfeTZUOhmE/Rgj+E99P
pyIZ+HTYxrD3VuklJSvzuZ9qByg73g8OdqWfiNwv/cN/M0h82JH5TiTg9HJFhN1J
yz8iOIPzaq35umJrbHyHZEv8HDykYN3bHWkUsk5SHYWjh67PR+XcokO2JULi4Lqm
NRiUUPASJ5suGwoY8abNfS35Czruyf0mHg4ahQtPrQCw73r3CyYVeyccLG5O8+1T
83Z615ieLZuutz8DIoR6y+rHmmUoNN+T8I2eLeQ//6QtGc/c55Mgza0W+sKwEXrG
OPU9zqrKwB1tMyJESw4iLFiTCX45cle51pP8oF+Y5IFi32HCc8K3F+sUO063c7eU
dCna+boWlPVezXzAxo1RHFtOktKsfBpk50RPleQkVMHrQcdcbubsq41DhjugBsma
+fSAzdxwSBtwEzMwKfQAihdIUXQdRR89ASKxrBifcBRhLE8qS87vdULdB+/jN01o
AvtOHp9M+3paiPywZAUi5KFAjwebamLyCxxbjzED6rMZt00rZ3lsMH5lKzbD+NvI
mBuo8EPUyLmG5lrh2oy3GlDzNrtEvdmHkz/0vWHqD/fG2/TDqvTtN12lNHiSYauQ
u4lJ2ceyaAnSxo7qpMRgtmyuC56CQhWkfBjKbfx/4mzhvB9KFiQwILLk2f0aBkw9
S4Ycnv3eqpTi6DkL1CA7D1dfcrwowOHkTuDzQL0rdRe5DzS8G8uKxQ47t6yiJvp/
7rsLgc/5HA9OsFmaZVNJMelEofTpqNN6p0lYqG93LVTd5vzsgLNNV7FbggDUEdPE
mD6NSILgG8aErH/oqEQqlIROrplg+SzoOJ0uHYYiHsTCUTcQ+2B9jItKA/OdRMZB
2vBvkEHLOKxkhfwtuSHESFYyiX9FC2HmSXzyLPQbOi9zOkDsfdPx4tXsC8XsKYQG
cYWidGMwER3YY/y3vhKNWS0lcXBBmpj5YBfcblDT2MT5TYqP4wLJww5mUY9xbYNn
nn284g1LHnOM4Kp5LID0ihAoDOLT/xli8qH4JUtgU771vAyIvN/Pd6bYAE57fgLC
GO0iEJO7PYsnws8nobQ37yw8xBA7IJGqh1wYO3IJez7pjMdRZXHadskfpDAwaCUs
Hmwk71KKdkE/IESgiRYJ8WG1EQcqEF4Y4JvIs0hGclfLnnYVI8cKjnLFv/beBrH5
w0RujdT8jeBICWXi21EwEl1hiUd2/PHmG46gFr2E993xUC3gryTjwCGTIZDCmAiw
80VH02mOO8zSwrWYIY1t0Fq/vWQwecBOPFCzaXH0EDeKvctJvHKxps5qfom34DyO
v/wYai+fuaBUEHh44cdEgsyf/EM79CCESP+rVgjE1EQDp1YMXcSMviH80yXYrINr
dZpPSLG6JT9+enJuLtruRS7sxeMNlFL4Y8Mk3nD/kgmesV9UiCcBLv9w0dlwwG9r
AYfAhFBt1hk35MRquQrFBmBszdmEVYv6wZQSSm7NFjLRUewp0iceZnxI8EODP/zw
x0Y2E1MmtHgDUzYkVumUmQhV0jQWAGOpMfS/i6YaWs+Mf+nL2jqM0V3fIx0yvulb
sOoCaRxIUpWKyvvWexLQiS5Adqy0xTfOAFEB7t+N278qef0Z2spQ9Aw3ztzeJpd+
`pragma protect end_protected
