// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gXdQHk9YkNSsI+I3nhVmnRrHJlppL44FM8DZ5NS7Xq6Adwan5p+xcrTB7GIvDbab
yI9TkH7eDWXmnW549Xb2aVqHpvAOKaqQm/feL8esX9P/KXC9ys37edgAcQJftbv9
FKCMzvV1lh6yFZ3oMinwU9GwvPpyQdZ6wA8zxZ0uVv4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12016)
NyZuZxMskpt4r01QyMUjcFFS/UMQrZxcaFgZ/RwzFFPkM39pPIqXZ3ckH9zcMhox
iNX1aPN5FCC2oJ2qc5LrBKbh/+BI172VyBRVR93e+NwXLpDbfTZjOPd8aF5F6wcC
D+Pc0pghSpeEfOmihzTEStB4yswJp9szur+X9dGZsnNia33G4CvAJHgADggSSNMO
Rw+tYAfH5nYSbZfctbs9TK0v+CstlWwD9pcFPX6JvE39+kIlYDuqIiBptwRNTC1+
paA8+XCai8F5D2V15ZU1TZD/HvbCMQW52BiLQJUNu0tKmLeLQbQpR4B0zjzSwQV0
GoCg6qOLsBOGKnC3lU9gYQIFQXCEFdUD4kXm74vU6mtljo6pOQXuGGEYjXNb7Gwi
aoJlljLKcJA23eBMUVCKKwoQBp2d0F+jPxdlwji3IiqGLoO2wqyEEdDcQSOUrvb2
07U4TYcA3byTv2hrRyO4G2v2oz7MrJ7LD7vVg60Gr3VdgyNDWILVnGg9wAjklBri
H2T4DBhNmMJthm4axDriUZon4UlNssUuMTgc0uOZ+4+A8457b8IJNxPBpMoaiYVO
rdfxta0c4M/uERAFkJDPs3kDgVXtJj5G+ehbR80y/OHofE+ATjhiE+HEtz8AMjqP
3WEShAYUdCqbnus/r13QedVUzdes6yr/kNlNb4G+6U7ZpLGjyoqf01KdJ2VKE9cC
qMq3UsC03HSmrfZK0/23e4RgHjN8SttjvN5WMNZWZY0AySjCN+X33c/KJhU6czbR
5Mh5JlYvGwQs5+8N4HzruMruK2SVSz9kLgSWIa7NCoJbxj4BHMk0bbQVqkMMjIGt
F6M8zVaX1h/lNFjlpNCCOpjSz/aFYEknWgACinch8pkNgDH5xjq3RnC4aR/wviuI
Vztkdj9Jw3QmzePQ0AEZ+TNcEBId5p8dI1r/RwqwxSKjtLIROL4qQJnc9qI518bR
MN8z1F3U3sMd3qg5OcXFw4aI9KTVhhfJxGyKp74JCI0+CK8nlof0mpVIYOBfUbWT
6sHCJVUw4ysPPHESK5TJKn7DvRuk/ucQos7afF1VfMxDzSa0xFF6uOlx6RlLCsNb
1Q1ksrM79YBSrU5Yke3HYm3+yAST8IaDUBU7Pe+hqi+AOfcWQjsLysz1ITRfl+kO
MhBgqOi3i2ZlToy0gpQmbO1mgjnGL3xAd+CMx4hxb5EnMpNPrUE21w2KwcO+IUx/
ihSCupUF5o4AWoT+6CxNTrL5EUdd5n3WbY24E0427wB5OBT4Wq82dw+dL+0a3t66
rRGudVtsN6r2mfpTq4A/edHpj3j3i++kk2YK4icM3OS48PnUJDSG1Z7NX+TYJMG3
Crj0ZNVJ0rnZQDVErhB4m5Sp9O5ANxwqL3nzML76xJbDWqBFqlpPGPXDP6xXhsuF
NZdPhbw41Cj4KaIrGDF17e0b61m+F0j8OBI1yAxOJhRliptcZowqUPpgvWrQ73By
4DXyMOzmDAJjVznXiq3P0St5PBiOY7DsbW8B6qrflWxcvGJKJX1FRAY8oQLrSK9O
ZrgxRox4//qTIMmbOhJV0JP0AxDrlM5ru7mlG/kbgSAQCM7+irF9zDpJQI3/euvV
lkRMtaUKKj9cOaaMNN+lGQ/OXhhtJf3agE0k0yE65/PYqsFLl29DMC6/tA8JMz1Y
8ktpVg7h5keE1h6TG6BNailxRMHqahcI7C1tgnnxQEXpPQfwIA0fujaNnpbilhwe
ZmRDfb1rV9exV6ewFQjlA5NdF4ep3fMfOlUOTNilzoTWDwqI9h2WeFy9M+jjohN3
sTb9//Rbw2LYMnzzRs6RhnyW7HFWTGs60lYSJrHT/NsQ/smMwdJGLpOsU9UTtegd
ngtQ88zlym01B1sd/+uMMtv32GwJJkGJvPAio0WWE0t36ibbvo6zWoRO4XQmzZqA
VS+iofbAF3pf0u3LKoxaTggGlCLmDFFJZAw1yRR5ZQC5lsARHCaEGAhrT4wbHcxl
13bA2cj7gv79C9V6lR18+lon+pI45Dj8hFJAUzQFIdZfw00wEXzxPh+Rw70ne0Y1
dwypFRCdWsOouSGbiWeEyvKu158qwMtAFIFSeYhSwPhTFzYjf2M9xJrinUcL2QsM
X/ajHpasXpR+0cZTU5bwn/hleax/3aPMimW0EQiqI4tO4zMtP4bjB73Dy+0nNjcs
3xI+ptxyN8E0sEdB9wVMQ87l4nL0AIOEVBOiTTVrvRHPib++Y7JFPiRLZJaWwQjT
X8Da+m7+L9N0b7PlFrsD1XXW0FsG3k1SY+YchOx2ODkBaOlsjzUbMfgQuyRZKn2F
1pWilUOBFhXCdTRGh0UtY/GpKts3ylhtZxi7/9tAEqq5JZwl3HhK4AcfwcCYd02U
8VBTU8Djsok2EvkzcDHk8AyKg/iyFuLxNhE1NeSq4KWkilm7CBSYStAsIHXa3cou
HrWVs6S5err+McUkOAFaj7vT2vnyd0Bltxrco4lwY16crYw/puKUD/mFgSdGQDD7
6l03pi7/EXD7tJkARNIXezqVT7ta1JWzed5TUbC/JWv13uJQx/cOKnBov+zKDHVc
S6XzNjWr/Prye5+/rfsAENJVEePaFh7zeh1BREb1/VmxIYfIb0e8QCv8mYob3gv2
/eD0wb7orowtK3wgASRyQcmo7qdJqT6Wo6x1WJOF6+LZSk14Gdej7xpu/KPL8FsA
Sbl4zXx/tJ/XZuL2u4FQURI3wAaPQnxW7UwFdmFw2N27xpBnvLiGs4rQFGwu8F7x
WkJ7thQksp6ilVVaKarL0RvzR8CP/NF3mxRcv51wvl5ZbVs8MGi+jieghzejuwhk
IRlK03+2Nzi+05mRw12Zox1u32rn8JZ29dQ2FkB2EvYZfGsvNTaXadzbgqguwwcM
3/YWvZvzLOQUgdhsCEp2b/DexRofC7UBTFliI9TJU1reK1jJMKaDE0t9HYSPTSlN
b5h2yffNEzVfCmnWyDr9negQEZtkVSTtjtur5hG2KzkFyJTsljXH7YhM29TCX7gk
qyDRlOJgZ6PnipCuKAXUFJt1Z+Z1e+Il0V7khGEh06ESO75HzGZijKsqVHAYGbY1
Fn6QUelMyYSs23pkEWebtlG2wXg7rgyUUslepUCLJ50QzN6lsHKSunYsvTo78AnL
1m+2Liel/bDxu4uQo7XwSXdnZqSzZAivMk+Qf57VlLbxj4VjjCwDOxYtZ6AIM3jc
QyeRRTlzdF1ssRMh10pW/8dAwDGjWY61hJOR//li64E5Wh5P9kG0WPYJ8nxOXCMY
BNjA6IpKN1S5qwnMDGSXsc8c4ACt+M7G5eUrCLoIFyr4CutwUEFDZsLmbp+t3GSW
0CQP7KTcQQTlN0BTn/pm+bT27IX/z3wTmPpOwMKmwBahJJM7zFLCyyIgpwYoGS8P
78gLn84hAgYEFtBBsWE94klYPuKvOC7/i9RCbZGiTbRKaMtOu7VKyjUDC76oY8oX
RcnGczQ0auNAy+hDfOe5IHhcGzNvJEMaUHe/QsPcQ6eoeYNYDpTqdX6I/9qS/AAZ
gKQBiw9+AcCET4PXr0/nR7HQujuzMKrLCec2eYi8oZb1EhJ1xiV6VX9tdBTqISRU
XjQL2uwBFFSmxf4Q/8GrWwHvahb1Hxj0AMbboxzLv0UNsS1Vdewzm9Kx96JAP7wT
HvmfeXdNucTfzi2/mr6yJsc1txnz2rrJs68MAhE6DlgQtRYkvufDFe1zyMUYPDQP
xndNw7/nfXDVpJ89xbUTHvaYU8dicYSaLAuKBy/SRJcCS/t2mfPJcb5xoVEJtZnd
f2dZ0VRvUPWcvBdErfhSJyxRMYsYD0qm72+1WQbjCPrpu5uGarQZG9Ah3Wv88fRm
+n2zRBouaQU4MBindBDuCjtNfHx5PBc+D7qRze+XkBN4TrM3qkE4vncxikUFdtBO
D+QaG0FlUt9/Om3gKAvtTcp5z1PFP3v4RGhhqE2B1YWzjtHKEssTqC6+VSaEXvF4
7AiJcPPadObbriVNlYo1qOoenWZCVWl9Fru4WOAJIYwms/aH5FA0oRQz+7dH6yPn
nGBsRSHAxjekxukhtFf8ejAaRHjaUYdQnhvUQ1URZRxwdmrDcM68j8ccui3qURUr
lr9ZvUfJYjYXHtvQLdqb5iSLCADjTlPlj2t0ZsKkk84kCAkJe4CPRbWZwDoKnlWz
0LpJVWzzp8kT2HTIVBYQUuaPV37q8L5skODQTu2PupzzFuy/HluFLvbkcIgyPJ28
6+rY6hlS6+oXwDbHD/LJdLncAd/7g0BjlSlPCQf8y9ED7JsC70QnHrFykL4ooZaF
ad8SM7rE2ncmSvSXfYyOS69JdpJ6MKzKlyYZ/ou6XnpCsBNVw5l2oOg2EhJLe5cd
BQHpwEZIdrEUmJpb7gcckrlKxcsroCOXkD6ZBNzZNk49YoLz5JZBU/HxHOGJwB+9
hPWRj8Su8R46N/6qlfe0uZ0wEeKaOXVc/ty3o9KghSzt1zSAn/EqWL3EWQSNd68H
lA5MyqSqLgEdLdLaSp+cULdAloU3NIFm3+b90wfBKj9Jy8qjOIOkuANxkEhlIZdb
VoH3Pi7sh/7fgZYXTYJnBf+ZHCKdQvQTfdQyLx0aeTJbKolfDOKBA7FxcHOhVDRZ
R5GkAzoDRlLamxv1rZxcawh66okOrqlEsM7RTus/SXJm2PlB/VOO/ryxDuct3sDB
cbOiwQH+hQS5ij4DNfU9neDpxVxIzjelm38N1iejroZRcOxy9HjbZSgEsnmbTILG
2KRuRs9LGlEkIcO2Bpj8+9jn4AcRbOaswUyg67tZ6e8U1v2JE3qkvv5zcI0mw6Mr
tF5t+4ydzszxJIFLGdoGosvdWohlWMnOwpq+e5UISC6dzDd/UAcXftwFZk1968wc
WUUqAfbfOduq5ZVUs69TcLUeY88D0VURaY3v+lJ7qrGwYk4WB5DEN+BFqtNvCX92
agukH1NjxqKpZQFywtbm7cRcUvJowMlL/eRjIykaxmrNDR6m2prRhVQP+yhSJQPK
AUs/awLtqgB+iuqxyWTk0H+v8Gq9bO7sFgsWBrlUMU4TYeEQfBA3xZybaJNb0iKm
EuLU0hjsuAp+C+I1hiwZ8cakYDqu5yQhUYKNGCTf9TnHsfWm2Xyh4KUyoQeEyccE
LG+fboI3XVY/MF0mkMQPa7oRZTvru/y/yYjV/T9myJxdbrVeBCCNtqqIjGNdjlfV
7duvY0OAuYqH+Y0eKmnt01xoevg8tqDi7J16uOCYJTw/MPqE3TgvA0+sEEOyClJ0
zh/hytL+P0ZQPgj++vZMEBbJJm6bumSUJxCHs+tA9DZvgBrAhIhWc1jxxzaPifC4
f/GCdm9nLUIgIJ8iSJS+l4ws05OMRZ6p0nrhXQ9lEu7WTB3b78M8YSrU8mX/v2l0
nkdS1pbUwYo+J9Db6OoTtX4gl8t8eDcKfVar/1AZnYiukZ3ON0TAQBVUCweoGC0Z
scRKhMMoNzIDqEETC91rsOrhvFE8KGpgq+aIl/jRuud4numtEinls6SURW+C6Y85
5qJCYM63qI/L/bep5tC7aDw88eIhXjNabRUSaAHkuPqO3bSYUQbFUA0XFxXBKVmC
zTpye/QVWFojJAwkyyoRX5Nl8sUKcydv2XYVauCquR3CD/Z6OLj0Mhm4IIR5Xqxk
EBpzvuwbxCe0OtoTgV7mzHPgbfu4eoUDnUgCWpuCM6iVUi7+URd3TJCD/mQ6Kr7k
eAJdB++ftafbPh8RpRRtPlo8wRW/0N81zKyfFx80GK0nB90v1qLHagTssNg+VQ98
yt0OJ3nOgBiglDtFUk25sYFMY3ansvHW1fCloNJogJmVE5rVBcNre/Tmt3fb4vNA
a8Qk+5N7c7aILwKME2MJQSUztMMNjKSWjYgv0HHycy2hr1ODCZvbOk9xNZUjArCh
D7w7kD/d3fBtqCAlNjYEfUJfK3ADQG0O0eCZWhdLNZwGiJhmGo8gG4R0uT4gZvJC
QeUkwPCm3ZPQugCR3jlJDItPI2v4mLeukXWvPWLcHZwkxW5xlhIV8f4/Ud3BG28A
fZeCysksORRTSF5JUBFBwG03C75rApxvM/qkV4ErQamIShJxFRAbLufs6V3eKGGn
RKmCn4OX4B4+WERyQ5evYb74ywdlEAQtMUFkoUAISwJ+5TqUcfIufyMK0oWXx4I6
3Q7MYH07eXCJNj1bLHvo2J1ulfQ8x2yZ58KiZdX264bNVrKA3+ltIdl0rdTd7D8w
5CjIoqDoDlCj9Lh/J8mzSVx18AxzPEeuR5N+jkQBtUREXqQnC2Ku+Sk0Yue2Tktx
6ZpK9U6IKxWUHnK7C2LVD+wdr9306ORMjQjeArcSH7prt/d56Ut9kuljACp3UW0t
e2l2D9ePjhD9pAZEMQp2fz530/B8SlIKP6BK99pBtJBhskIz+SJkiy05WSs8nfzp
PBbjkpGk81TGKjEDclwcPAtYA2a9VWvPnFvUxqbG0h+G2cISKYHAUBR/RhXaXD9x
8yjtRVyP1SkhNfOVNz0FSRFhDNQBriW2pp9duQxfJ0kheqGPrsJhe323PVy0RgNb
xjSXLtJ7xPu9ERtm863hQzesvHPJqGx0jlpCtcFXpCt+OcXC3TCu1bSeinUCjMlT
r3PnZweH4kF3K+scHAJl+qiqffjIck0HukkpvTnSffajiMUeQPIly0ZPhgHxGLOo
COhSuxkpBpJvaQXOYxcUMgBddsj2mUwqWCrtz8n+Jc11OxtoLn3aylZvzxWxctnz
nrBKyncxfsqkf46cRCGyTzQhIpuaXkC5oBmHIqsNOecmUatGAOH+uvYrI9u59ca8
zWBgLxRt7q+XfOo9x6AHWCLQcYGVxsUAHOAsZEFgFVjlBsLRB5BeotLQKzHEzHos
Kd18c73KHH6/loK9/zlAxmIgi9lfB6rxf95KPWhrvT5dRA7rO2cew/qD7mh1pukR
kcioKNeG4fe+J524oycF/owUHJCHl+50C8wqXfxs5OKOw4etjWZX8biyZ0j892+V
Vd9i9HC5cMDVtdXx1DpCPzR/FSAvoclLxOCOn7xMlo+uB34j6K/P5a3EFsaSvVAn
3dcA3tAlz5FlqBpSHOVinLr/kpDRwwcaTRPxRifLKLkf/pkzIdpWsEJwYBYwQXhC
CwVv4Ijsgsu2ajVYGA4yHWpH1wA7D6LByoDGvzl9bAGhjKk/fJvrXqNWaWt1u4eY
188zVWgw7AXBX/z/JmQ8E3WSn2p7N+2xkWutY1r/qu5ijLg/mMiMn8ptoUajd3dh
Fnw6IPhpJ4phs1/w2HcN9/2/RTAS72caY/gWloDlxVyiFAKf2U6ikYqThInW6cap
30+pR+PrMuCaMFCp2I55fbcJVk7Xw9bU35Vy45JElU5zbV+cRh1sCB2TpSMGUcH9
VSy8Docfm2/v8J8N5olylRFkSeEkJh5c/2AYOKDVE1BLKz8+fFqU/s4IAaTo2OT7
ptaeOrZ7SmwQoWACS/TY7tKy+NGei2iYo/KpSCxYdvP63pe8QEL4SmhMpRJ7f7a9
6a+6DPtcaqgxvYAqUI16m5l6tDO9OZw73jJw9WZL00JKZFeyZIDGwllXnCQoVmHH
5LiKubEp0wUDQcoRShnGl+pXoZHw/oih+ZW31sLCSmEFscvIbSyM0lcu3B6Vf+6Q
VtlsvLwuR/xNvPefWxkLesF04j2qoKWP4/B3HVlxwev+5mTbxIkuBk/Au80D2dxC
m4utdnmDtrF5jnt6bDtZ1/D31cVv/DooQzikwXxM/wVK9MOPjTwZr2reigudCRWz
+sv1Z1S5sel+31HaEuEkxvPw/oXabIdJzqCjODDj9ptSzTF+osqp0a96xJRvgyDC
o0NU+viaxlq+BqWXhahbHnqS1DSnwkgFOtOUB5AGyfRP26CqAJrsYVgBsIfN+CTd
qdmgIfSEjEHfcS479qcvAFcUl2Y0AUCGC76km06xDvAcdzAUE28eCffTerLHxTWc
pyPwbU84jppXnd8qW1+3car0psUZXNRRBXTDrkl9h6XeguWbFdSUBP2TSEDbIIOO
uLk9Ia+qmVXXO8kYmeK/oXMMNSxekj3pnQKtHVZ2BUSU5464/1B7EQZ3nuiS6e7F
DVDouxowdIT8hOxHCucMl2y/MhxyMKSd4zuPStxPL3UbLNTKtZJq4MyxwzgGG/sv
jIOTELOhboeku1HsbfeA1kSh0YXbQLOeCSDWqzxpJZchOkWDWDcOfOUeZ8Uwdu0G
15Vw1aoGvQPquyQe1QpOb8R3S0bXlj/DwJ9McZNVD8F15EoG7pdSbmIQACPj8LE0
N5uoL6y4zm1Bn7dndSQ4ARbo06icTO4FXdKxcq5q/taP/4ffb9gyWjvsHfA3gvU4
cT3eOfCWSLYctA3XqYZIVSRWCwez8ZgUSKZBC1XkhwIb95MrC5jXUHWsjX9uTjRE
42QwufiZFciNulCgij0Qw0NECWRgD/5unbjZzDtXpoetJiwZ2cTmJpTXi2lJaPhd
64w6Nuky8PlGg5aGw+Y3mDJ3ib3rEX0Rmb3GOx7k4wIVmpVIFLHWASIw+eSFnJj5
Mbulj5mtAoiQc3zhe06ffORCeg4NE8lHRDCpc8ZryRY1FUjfZVNYWfJr2Egck1WG
PTvpzAHx9tYPwnZjd5/9g78+NeV3hVKX6K50VyN7BpnwuPcuMD6L+NzBhN7SwI0g
77TnGWgSHegoMICAYUVvPHgIF6ekAVTt2Za9hsR7AnfHYaJXDK0u+bTzGNrKpKvj
JPc3xP4jOvVxYVc+YZB2wKb85L7yajY7nNXlwQiIf6AVaPFpbt/tJG3aEr0/EOWM
bK6cNNgg3jiLLYZC5C2FYjNO8qFVuFaLnNL3WsGUGJlWDhzMMm2Uww1Ls2YuQWLp
qinWcl+C9QVSpOi3qdscuzi7fCyf2Ykeun/x870zalgjFYCEo8MEkTdH5OtWclOL
NuMM0DO/rqpWilSBXlBIinYfHavL2CpM9EBiUQQOpk6l6YeS9nP6WJup8ICceUKU
HRzjloAmpd0bZuyJg0LikP/DIu+XooelBpOXYqzjMhB6+5qydTxgAp+Ieso1L/SP
/fdp4xtPscv5DVCSUfcVyAGtwXpZurpJ5tYdGKn9cw5lO/pF1TMvKpvrSX5Se+hO
QkE2zYMEftcThSXJ22IN4H9Kfz/LRBvV8rLWBLbwwjL8YpPf3VKprPpdr+Df8Jww
F8MLarhFZ6w3e6lH+gTUUJrcyifAZLpmUYSl2Mrp0n5a5Ej3KbHI6gUNZ7kb6+sc
4Vu7RJAneaEduaSpupumZxwxPPe7ykCzm4+OudDDuHNk34qIz21B8Ft5ZfpcbvFl
47P0Hk/N/CZ82t1ZI0yXp6dCfgKXRKQngdzlwK0gpDOPWcrFabkdzCY3GYbLsyrs
n+tKP51Lcp80AG1w+yK9+YwqW7DNrmlFGvwMCSyhRZCfI06+y54ml2csVIix8t8x
AUM+iws7lw6OVcmrakS5XuKUO8Zg+2LWCIzlXizSFZ1HgLTH9BG4wP+fmths8x+4
KXZ+JQKULk5K+nLNgOf7LjptKORpFaD1WyCH5O4Omya57V3OEGAHb+VL5zCBgj7G
Z9iHqNCt4YOuZOOcjbYp8a5fXiU+NJBSyYk73O673gHsaijs06a8l3uTP++9FBIb
X6Y6U3WHOfyVBpuL2vjOp36I3X/Q9Cbq+reEKIODgrw4Q0l4GhOjFy1VN5TTZWFa
h0QWr/rGQw93i/oIlk/XoKGlXKtbrgBXBfXiGwcQ/NjDCQbTTYO4GLT5QKi+hFlh
e3pjWThNNSsTLJT852rIJxrR41eg1oUNtQEx3b++E9VVneySi1ctkWZKC9q1kurh
WdI/G3AiqrC7iuXmFgDZKdIZ4p3KK2TuWTLtdX2BxTyXlMENom3uzOjmxyWIQkL+
IXta0H7+eW1z4Q/HMgRqBnoJA745nshfwygUDxwbjxirGh9AFbp4uKiimHj+eT/6
earstTjYpwGtJpBvwI3IUUxSfRGzjD7wZHlwOmhkEp44Ue7Ks490YexieIbxs5rD
aZ2P2gr2ccFcAVYpGEc3WPqVSU80rr/rhMOxWOHHhSG6TWgWtVM33v+bm01iBASw
4UDuI3tRhx7D8r6LhYc/wvVGrpwQsxMKBaB9O490IiKFgn7ho8Q52cwFbzq23T1A
oid3B0JUkgq9V8Z56VxosckzHeXufyETs6X+/xDoNnZbAA5HGLvN+3siQWOPrJ0d
/2w5089klGNVDiKDhEwOTjAgaLvmdA69MPwC/pTuG7XmjfkkH/qCa2sqHVxBTnOR
p6G8tJlIJ8EuZ0eME2pyO3hyFV/ZFVwZl/HDfw6QCOuQbljRLTuy4PhgrjNfXsvY
/K5GIxzsUjGzZuGwNiqejlsGKYdkDsLoazR+AQjonqNpKG0DJ4i6/KAw4G77K+ks
c2poWpBV5AQuEf03SbV3PPeykUqSPrUOhLsFtvjlYYOdT88WKV1e/UVYcqkc7NMP
BVmS9I3sjtG83oqZ9X05kzhChsABkRgdLqKSvrStNpbQUFWkTzbJhoEtKyH9DihQ
c9nudB9F55IremKR5k23wfzAWz4hYIm9QtnYsfjE4AvEebIqt4uLns7e9fAOsmED
nl3fnecMoRHBY6X8jQF+YXBDdlbf7UbDUBu8GXmRBJNVGt5uMw30Tc4qOccXzQ/C
BHMm9B6ki1zpIP7RIbBjI+zLozzZ7LNamQW+pJJiUdBkyvnKuMo6tHdQe3xESwUN
C0z8I+6U2tN2/8aUEvu5cYq2kEpQuVx/eUKhgqRDy0ixYzUkaJAFUCHqrz7vpY4J
bT+FtB9VZ8R4VyhuteNvu0jKNWgcLcQYEh5Pd/qaW52dhlBUEM3WhfGfynJD0KUw
ucqsvCj++LLxPM6sqAusm/zBvsB8gGxSSeeB6wIP1TOrAG2NSrQ5DzRhRUY7GT/A
kVpKpO5k+lSJn1cQXOf3xEyLP2AkdVMBZpa8q8m7+QXx7L6CGN8v972wCu/QR0mP
6mX8k83ogBh+eScta2NSWx2R2rq/HV5758tzJulciYPWR6SChg0lWS9weIP7Usmz
H8dc0uy8+89f+4R1QxC9HuM+aWnRyd1zCmjcRmp04fu5Xw6NFStb2ZnBnEkboBQZ
vJYikIgzBU7Hk83DHM1/zNkS9f8n7eHimQ/5+/4UlCs1yxQCu6C0fU0fKLq6jMJ4
sqzUXHKNywTBg4A/xjT/aloJLdND1Sg5lvVccu177TnZ6dCs9oSsMzeqJO+zwh+a
alSfUsMtHzTLDMvIe1wC2dPE5+xdEagMAyWSBxkfqTaWQAACbW/ko6v/QD9AsPcU
hduhU9uRNW3Mmu0JrwZxp0yLZb1imhqN+VAEDw4Ankcw28edcnSDLj9vqXHqYBKX
Ht1G9J0P38thoPcpY7LYMdtQYj52AMNu297x82OiuVLeL+rGCHOGsJN7ydoiUJQq
eU0ILER/AdCna7MyDhasfe4UnjI6BkbL/NgFR/+fhl9e3WqF9CYbli7VGns5LkQF
Hh/7fvASTWCpsQhWX8CRMuCVgtPa4+Q6aDKLtK1sio1gflJGWenkT7l3JwwmxOvC
xaxoQplTsjTybQ1ywwuqpJiPzjaqh+vKvFeFIeUTys3k6qEwvQUNPVEU3GmFso8K
l53fZSQDyOA2N4FebDjvTbxQ4700Ym/T9BFQ5XAqv65+f1FIQQUO+9nhAETDdjsB
VphvJA6X3m/JCr77INc5yBkkfBjeX38Pzq/6kgdq96+eRbb1Vu/YchtU1c9U+r0v
G1Tz8HSqFT73MgXdMq+PgLjtVScrJ6LAUBGka423GO4ocTMPS1LQGuv62+cvEEG3
cQ86ZtNnFZE3ZsXac/2r5Z3SNZYZhzNxRlgN8vWtcNg6O+K1YGzocqQhZB74/JBt
p6ktqBs9XNM8u1UHD7NSXoLdRr63clnaNp8wA6v3vWhfZ+XIxbcfDfeQZ8ZBMWGo
+gzJxZ8vNlzS+UoXpE1BY96ObjGnRQp93deQaHlB3qe3LHLcPdGj0x4NLGRojLF2
tL8tfE5qAI/UI3lekIy+Fg5gnYoLp+ozqHWNUJUkofx26zJvdcZ+WK2z0FJbqRNP
frX+yreKgaugaSxKB7NaU7u/LT2Boal2ec45tSph1Drdjy/e55jzBjvz5/ORvSzb
yRYyzF+DVRhQxsARPpB/GWY/RiSo3dbeJ0cC8/jml6oJfVy+lx+ptEAJI5F0cucs
slAULWv/hJa6+FQ1/cpozfrtDycVj9BwasivXJT1ADFv/ew90vO0On3yVe05NivH
LjYnSUlzji23HdAe+5R6J8XJinellq3o8jYiubIf4bkulDR5mr2a5W32ugvbsWXQ
bjuvQOArMjpHWdFbR7gY/tKbUrzlsm8JiE/j8GVpZsz8mbyZbtWg54rerOUYyOUX
oD4KKWrvl8wkP85DMUJNomc9XdOnoKM372VFePR7z+ZNI7NCgm0LUtfh4HroQFZV
/Zq9+1pxRU++iaPl4dehpvDuV44PnYkeGVt4GiqRjUT0U04cAlhiGCXy8FN1OqAj
lx5OUFChi3lEgB33rL2ylPyo8pVQ+QGzjz9/4kY2pSyXU/I8LHRinC9uWR6xwqyC
R0ajaBIZbF3ZPEkU/dFAcXdrETg650ScnPbkPJPwLbmA4y9rjv8sGQ09sCCZ3xbp
4fQtgkfEXlhDYUVmMWLBGv3JDMuxN4pkzsWu0+/BflJg9RQy9QY0RMNuvr3ZTWVS
8JpOi37j0b1MXWgRL2AHYYD27uKTg7ZBQSAzwWpXj1AGUMJ+yshkjD2L9rP2c9yY
e2V+9yfvR6Mm6EEw9CHk4lGta52QZNL2CIe6Wu+VDXJPNpqGg1pLOjA2UXxkXZ2g
fbD+dIIrnLz4vzapKs6i7xluN3QWAnxm286b6YX+RZ+u2mzaC2gQ5MmZ8CAOzmm4
AlnU2Fc21MqZBAq4jTt6RC+S2+TJQwfdiiq60v4MU4Pf4FqErcYquTnk3OBGaIIm
2yAeQhUinDCsrfbcad0mtm9XFxl+xuBTT8ulqSe7vxoOcGYzZuqnOlf8jtxDFEd1
+UyZsQAt+/Obri7IiIDOJfdbyODXt9XwsqotJDfft2dzweuNTpq18nIT/+ZyHF5Y
HXM+JJ0trLMqIiYd5EfGYRSn1jfha6F+NlGmuERv17naDh1t8AaRxdk3s3Awg7an
c3BpjBosB2Ra9JMgPBmJj7eiZJacWxFdsVOAkWT7AyC6e/PmnClDSAevI8ZgDZAT
/40ojkzj969SrdxRma8K2hLKruzGHRAn4E/Q+0SdDNDO0F31QP7hPDmgf15yGch7
1CHQxYYAXewdilTywxKTpDucAoEAdRiNthQDZ0O+TDWE0is4EEsuf9xUqZNKsnsL
/Dt5ojMrsxn1kwpR9Ha4cyY+dwAjrXqEUI6I8yGOE5wa/GGDLJ43ixTe3x+W2YIb
wGVD8rSmS9jKBzzgMhtOXCnWrMbcix5ECDSgw3he3easkBM4fx2GtZjs5Mvh1xko
pKp8fSIlSw+yWg9an77QArZQVkb27shtifljHsRCac3CdC+GMxMDkL9eRLu0W6tp
JxUi2fuTBbrSVwmb2ior/44Pc/qj1CNM+sOGpuT030klbEzyGElEGHjUd1sHThnU
FpN5dHfVgffEwrzDex53aI1MPA5Zk0+G6mgzUt/3g7s3t6Bm0ObnBbslOOZXggEY
aGcmmQilwiU7syz0JrAyBkjOMU6THa1jPxgU7DBLJSEdEa6QrYtHD+u18QxtBoKs
LuCaVDebMsxH59OXLdfIAK5VGMIl+tBSJWsfIJrhhCGy9i3Cbs8zfoD4DyXeeqb7
kybbwEW5RJprrHKmkyaMSLtrNDXCcrUlxq1GiQcw+XR/ayBEofNt59k2FzLDsH3x
uW7zGAZNj2LHSunw7ZPWrQOppnL+f2jACDyxQ+ulmzH5Bbi+F7HbuOPRTRjNPZOo
U5kMeSeIFj2pBzxj2BcKAAWOU5Y/ABotfwLkkKswtjYq+aJiLWh/wSRxkWusqpkl
pnbNXGwr7NgnN16hMHUAsIU46E3OnTugGQDfdP8ZfZnrLvP7d0fM+nCSGiyFP509
5zusNvI3XaXnjRwqJ6T5Sobr+2ZQsXO3NVWaPobrhjZxfTfAugzngR0Is3sWNwsx
QBE9U8OQnGvwIv+930yljUdW3if/HkJfFJpkohXBCD51+D8biLXyZdBLbY5fbKIx
J8T3Bcy7N2W1EQjHimBE2B1IAJNpo5Jp+cYAsfWFYamJhZLk3Iy8URzE2ZEMePAe
3ldKRa2XdPdtBQqVuA5PQFpekeHPdraRKALL5Ugovkl7nb9o3MaK1mbpRf/2qnb8
ELhwxPg67LlYSR6CyC4cc0BjDozdhxNV2a9clXuCsB2GiGmsN+KJB3cH/GrrbT15
qkhLALLFZRxaYElGx5c6uMX84w6SVxBQXY+8eLbY363WORWmp2qQRjbyzksJl5hr
SMRv6r0Av/OJIabqwneLs5a8ulRrTz/5xsOWoqHxMmzzMpqGtd0uBxysyLEoBTQL
LO+STPhjWVX971+jRdnBxROTeU68BPPuoM+Bfh4VjWqXXR2Z3mor/A/E2yksEuTv
GZz3ywhSYImi6sRcrraB8lVyEoCYjiJw1DzJu9ht5Ub3iSwVgImQBpGiKS2Gehpo
QN+ZuJnYiw1G10/t52YdK8XYSVFMBbAvwjAT3tWpksNsnkE9Zx/iDaz6Z9vgCRMn
zyRrmb7CGENCYzmzJYcRLuHbNU4g5xedUh9XguoKTD30/O+w4vvUBWdE8xIPNAVt
BQHHiyKCgejyxkjn8ANAV7zMzuRzKU4pZR9J3qGS8sJv+8AB7RRDPy2FHpbB9MEF
pGnhJwzSS/TIrjNFq2fKxngG5FbdYGuoBqSyJEF6WDZoXEByVkj8YjL1HcCIe7Oy
UO855CwLKZmjX3TwV+1jHtygrh5hz6JWj6MRzQf2Mw2YcwJ3R0wUwPuVuirB6F+o
9WII9D/l2whSxAJtAjtDM7sI0XA/aeLa2w0ns/aqb9a5PMJ7HDXjux+vc5btiHIC
Cr+0hJvSovEIQQKND+XRUbOuMQjFtG/FajKx7jscuctp0x045mWsJfV12HSuzQqv
9qIMWWumsbGmgB74q7xK5h+SYIHmmUt2VfI5IXYU4ewpcZNsU07cxj72T9vYUMDx
suN22mRW6kLZ7blO51EAO1fjxXrsDFXISNC8m1S5p8ElZEQx/Hf1fc2Ws9i0vNhq
xVPeLs4hBzFzb9pHAxP4qCR+aJ6ovlHNfxVib7COQPcxy5aRi4rlZcbFozEmnFbX
T1Q3PZLfWFLMDwyOJY6Wja6cvpb7RuGMDABjmAKQIkLw7nZnPSwNM1UOHaaNtjHt
b7hfiCSTOnT1QbEJD+2QVYoHV/dHNUovMy28r/qJOt4eAvbDL12Ttookb288BNd5
TwdRPzPBF50RPQVI5foeRdFjIO5Z9P2mkdVpwgJwmDI96kI5aijZPzUlXJI4T16w
V9JxYXX6Rzv4y3w3RiR4lSy8sNDrclLS1OL8/7UZ/+pNerPIV3CJrky2nZZYN5Sc
76H6vIYHFl9VXz4pG9DyRLGFxReY7A60jJceLwIVGrsoBUbVDeEb2Qojknjl+eRQ
VlvAI+4Vj5ymTemPO6LsfBvTqzBa9Boxc2ZgqTYGzYWhWCqhOMgjFU1ZH7JGoKZ8
Jz2FH4Z3kF7jsbsyHs8O4RY5qVRwYmh3pfWUDEGxqZUJZ9MbnZWO2JGFnQsBQF70
SdA/JYWPNNvFBPZI90nNFX2BEz7sV0pQFqvoRDpkXYrPCARWweI3q6yK84xBXEO1
+tHIMtBXUuOsRGUjhqUGeqVYgz9Dwt4W8K57wKR7YjnSYkrHmaIfE6L7EVMUMcpn
jS1ODf1PeqidbDDzXr29um7wp+zO+Rkf4Hk5Z5dAfSj8o4RQgQFNbCgQ8dvw5DOu
nFMccs8EPQ45yPo+Ki2L7tcMm//UV7+GtEPCS40EjXYBkq4EvKQJOtXOvF7E0xgb
MQ4qluSiKHSBw7PyHz7/F7R89XNO8ob4F2a0LWPIH1R+1j7xZ0rXCkeoPdFZ2Hh/
X+PqkFMHkpfZoFTMSq/zAA==
`pragma protect end_protected
