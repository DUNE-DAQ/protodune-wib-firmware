// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H^%=@R(JG72^5#OYAGY B^7?Z*94E\T6/TVN/=0WMP<PH/I,0"F4BC   
HDH4%H+KZNK/_0H>CW\^+S.%S,$NO P/$)?R5/^2JIRR\H_1 Z^#:5@  
HW[4?;/G74W6YC F%&2C91&O;@I6;*!4F*'3K0S>7J^ IUD$JT3BA"@  
H@%'Q%$B-;*=H=R_V)\L#QPY=IE%C@)"0NZ=[_C&8L'$U;-E-%N\S:   
HLM97O>Z?C*]@G<M%%=ENM?5RIGF7T+W=S&#N*P9O81JCIK(V6/G\-P  
`pragma protect encoding=(enctype="uuencode",bytes=5216        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@M.=WR6")]C7>PVHV?K.39/C0 A\5$OAL+^-V*/ +](8 
@)'WT'(LO9#X:4A8592@!ZEFL]G[P%;"4#MLEMX-T9"< 
@02&T!H#!,P_8B6@[[GC3/DQ]5T=BB; 8_2+>B'D1C1H 
@,)1'D?^PAT\1MOAC#_X""[/!R%Q^>Z=<#Z T<X5137< 
@(^<$D E6?7L<M\%V#8$@$KG+5$<,Y+:FFI*@@6VX7B\ 
@ <.WW]L-4(B0T0MA*O11&YQGN2ZPT+@*G0S\7WIZS\@ 
@[8TS32L29G-IQ!'+Q]RE(":H F$R/<?!S2S.ZZ]K28X 
@.\SJ*FW5\TY P4Y'R1=_3^KR"OT* !R99=G#H=Z.(C$ 
@KU.OI/OWG]Q6T1X *BWVD#CP),\. 1-W^,@ C"[(J1( 
@4@Z?Q(.-@]WSK4BU.EL-U@8()KQ,^:'0ONANX],R/XD 
@A<S#>+SEGB5\7K0)I^Q6P+&;5Z3($!S!=ZHVS6M0$6, 
@A?/S2$E-D2('Y9[7Z<R"^8IC=+73))KHY$G>S*#$]"D 
@* )A8/Q+EPY)P%+&BTV6AQ0@G>5+N(*0XRQA3-&_IYX 
@O]UQ#:R1P(JK[ 3 E-'?3$ ^4-F/)\QL0;_F$32M-A$ 
@*_L\/W\C7P-3?<;?VZL;-5$"+9B:<'=9NJUQ'H[N/FH 
@S%WFA29L%R[C8%WB-G^0B<^\%+%(R5"C90!(DG+CG]P 
@ 9:XK".">*N\^R%OE ['G5(1R:H/4BX/L*6X*VA[Y ( 
@0'#2@+1PQ(1:=3:EB9VM: 5F<5VE-].04N2CC&P1/AH 
@K Q.:Y1;';Q7SCG]"@<722A%B=D^K$\<_XJ0)Z$5B*H 
@A0)A2O&W"Z<+G@WX4S]8TD9MA3(9?M'<)^[1OJ./2YP 
@_$?5*K<#2D2O=DT-MF6>T"N8AQ3R&T#F1_*F@\8I,Y$ 
@YG'^4K4&H>[0$W)2_-+GX/F[U]7(]!X,=^HVA4A52\L 
@PTDP'F;EU-S:%KR<9>[E-K%H$="\LC;;K-NH)EW&%B4 
@3?6M'B7%QXC<:1MHY:0.?ZR=B+"?N#7"GP,FM1=GN*\ 
@]IXH5)>(OD7FP:2E-B=0!5C6&2E;TP5RJ<1^-O1K]6L 
@$+<MI1,LG]8?J3D+I ,L&$.NO6<XR,SP'F-JD*.&4>, 
@[#=06H$G[]U]5B9!F]3EY2'6^%YMN._U*B2PHNM*'>8 
@I)Y#?5Q7,/9[,B^ ^5H\]DAT5%[_I;[(#CN2+<_V,84 
@PTS6N/6Y,%,JDGZ?MHO;1DP R9Z9=UV5U1S\1*!',VH 
@(7\K@QO26J2K1_%]0??PFR4#C5^J$3SI9=25H M7R^  
@Z*U)V#^L@Q\PDX3F:4%E!5=PC505Z3-M _TB'[I>O(T 
@*9P:V;4IU*=*3/Y7-\_U*$->O4"S7L%\MY36TVP?AN< 
@.]MF>K/GCZI2"&J3M"?<3;0&.(43"R)0V28WK.5^938 
@][W^^O#;V6%E;;K>/2@VT*1\.Y^SGA<&9"Z9'%H^D_0 
@,B@]H"TM=E9<!9? J:(>S4-"#,, %<: /9R99F3-U=T 
@%2J)^8.CXH4T"0 ?K1+!8WO>O&B#Q%GU)'=N7E;]^O  
@J['>*=Q])1<AOET:Z4$J620!_N7G$A5?B$'OJH'!W"( 
@*[JE!HVJG<F7Y[DGPB62P/-C4>HX!O"$AGY$L"\;=>L 
@8-)*D?Z92!X&7^#@:_QEG%2/_7-Q#,I%=FG&^$T%^ @ 
@'')>AR!(_N!D59<@ZB7F+R^;3*2QOCRF5O!ILYDF!&0 
@$1C#E?N%78&3XL"9J.G72J[*T;<$L:E YBM#,FC@@J( 
@%%0UY=BFGL<4G7="+3#Z6Z,OYY\;,8J!Z?G12P$#)R8 
@<XRNE3TM%O8NWR_0E(KKE%4S(#?=:)M1+X4C? 0^P)D 
@,JU !@H-#R%2S\U4X-25?>]$=[*>MKA17W:NCW$^=U\ 
@L.E#RE#T6+3Q,_;0!Y7]^JKRWJ*,C$TB'(C/@%YV3/\ 
@;"6G#!5XH"X7.CUPE1SU9(9G_TV?E%:O+PC#5]ZPA8$ 
@D%)%R'>)XYYN3+ET73B@O2CP:2T.&^PN1!"LWP<LA0H 
@;7]MHIA_4D01>5I;5+4?'3M #=]#]XP * .N6Q1']=T 
@WL%NF<N$-WZ2U6 I%J(D-*C)6?:=7?@ "NF[';7I&WX 
@E4GS.??-]_/B)!&$A ?*P5<KG^D3E!(7!*\H,;I+J(8 
@ ]1MA[MRTP[2)!&H$]FA=HPY@4V*.".Z[DUF*"9*1TP 
@$9/!N,HY'4!8GZENGM=_ZSWZU62$_DJ]"P\8REG\M*$ 
@&BRMSL4T#F;B#YQI$F+/NR%VKN+#:/'5TE,$:Z((!?@ 
@.;M*-\+D*7J\:EYN>>RCKVD]C?@!<17\$^5&X1_;T?D 
@33I-7T((E]59:!U/)I$C=>/^3-F@X>OZ(-B&)S[QOFD 
@S%L[:\$-A[UR?(GXC6DOSI<(G!FLY)36\%X1,RV+WNP 
@(,*]%D<</=N!$W$)N7CK#=64=^;J?O<3'I9-Y8&,#4, 
@)ZY+D3#24-BFD/O.MX),V!Z8)9%*=YNIHV1%<]H> ]L 
@4P>H2*5$*&"W+SC+:#-6OL-18.73WV52N0J^0O7HPN8 
@+C0D]F)$PY&_%^:'(/"CP?@O!QR_4"$O[B]$ZO;?]70 
@<CA]FLKA)=7CR^CPQ/.M[;&!H"=E;1?5NZRV!;(4?/8 
@^V *!&3/1PLX%7)[@,OB:I*6%Q71HN8R QY:+?NR> 4 
@9AF?VP-\>VFHK^+-/Q3/3^@J7IZHQ<D @'H.OU,"Q]L 
@']E2$_EIUOW*9-2^(79.I]WU67,;1;,L7C!SPB'H"D< 
@L8O8R:A*#(%7TB>Y#^AM?T/T"&+2@4(H<3!:A79#OY0 
@(A[64V]R1M[AW,_VR,<2$EL?/<T3NJJ2M?#_85G'0'$ 
@DQ<YC?2Q+8$EUR>_$\=BJ @9#?=T'I94RN)*'?\2<"\ 
@#YN=?CQY(P^>*!#1+R>[. M<,6-:B[E/%HJ61H"9'\$ 
@$K LT/,J,SVNL0P<8DJ(\)4NZGH/D076$KIRXH1W7:T 
@D_.S%&UG; L@@*BQ9Q +E)^B1^N6EQU!,;'<;SLES#L 
@QGM[:L6P.Z'?X5_<U\3%K!1?:>S"!AUL0<$D)OB(E]\ 
@S8ND^YQ@^=E !FC7V\./DG1TQL'8=*/" (N.YL#=MF  
@ .  $@C;4]VI6F75ZS.;E_NZN+>NHS^IDBZB(U$')V@ 
@6V7IMM^S3(Y7H1!R%7EBRZ9S)+FD/(OWR-O=%*MMUD  
@H.>F]D+D"TMSZ0]%R>]G!GYB>&5DN0C5M42G(PM)++< 
@Q.)1[$V%P?\/2^F<!Q+N5MJ3.O"]B5_ P0UR"FJI#0P 
@W%7]/RK3J\5+"2#(TZ:6D@.JP_>(^G1.OR<]-YW<K&D 
@22NR4Y5KZ!7.+1)+7\[7M!'X6(_X3=2-W^=/J/'#!0, 
@SE8MX<F!(])$V)SV?^6:NM@]!Y)\@7-8KD]BX]AL82  
@J5UJ2,S'<%#MN;D7H_G:\GJ]+L_@*^*"T'1E$^[H%38 
@78KY%RZZFP&X-XTE>;RE&$RNGC,9"0*6A^NW<QDDKZX 
@1T9]LK"0BWS]4O]AKX4\MEM?L^X70QN6WS/?X=B[0%, 
@:/EV9=6VLW]8KE22" XY:D[3[)%C29P3,YZ]AU8.3S$ 
@?4?IJ%<=_FO2$T^NC0*1TC6]PFF?A92CX26Z1RDJ*=@ 
@C3\%[XX<8Y36'HYXAB_=TS1]C"974_@X ^1RZ9!^5OX 
@04^YP('^??M!;0F"Z&/^4L+H:_\&2'LE"U?ZMQ=V,]X 
@^0=[_MQ V7;TI89L>:H>KB*?<LHYR,H7G7LY5_@BX , 
@P%+7B6DU--S0V9$PXB.QX;25X.MY(J)4X6IY.UIWBN, 
@+#RDM2%D?#2%B;]HZI3U:[#\>Q7+)94+6=<3\M ");D 
@F>I"_A<K/D9_7_:."B9 M-?<_D/G[+[@J7,LA4H?V7\ 
@70UJ!-1OPY>Y+351PCYSCFR.(S##?J08WO6./R7B;04 
@ ?U$?3,(_M5CIT+%TUU._FQ1CP,N[I=KZYH(F3B!>WD 
@H[:"!<4VJ#LBF]0)I#&O1Z>^XK:>R*6E2VR5K""0U:4 
@(EM7@@(BWAMS3B*C#+,*<5.7].PJJ,2V/>,0XMMU"%4 
@U]-!+6&RE!B%_\)1 U32'[Q71T%W#)#7(OJA2) N<C  
@8]>B7;W_(5>B);\"3W1S"+XG2YB)?R^.!=L$2-N/TCL 
@/8US&=OJSO5;(#3SER%2M7Z>GMR:-9%^P+(GE?,\9@< 
@K$4Q^TP:^6@3?5D#.'%I/,:'B#()V_5*PU7$#2NE:]X 
@#I$L*G=I74G0Z+,3*1D3SL>WJ@^9WL+J([?3X.7)@>, 
@=M!.V-ENIG[!4VP"-XM[,E_YDI\72X2@R(=$ISRI4HP 
@M-=D5:Z/(.MD_/Y@9M-2.<+;@DO_$HFL9@X4X,5 F#H 
@Q@ !HOE D2FZ'O/&-7%CI@M^$VHT+IRU#Z*;7%<)LW\ 
@5N$D<9QO*C4P^I@04>?[(S/3G8^/=U%A;-__J!:0]FL 
@*@'NW,'0@';JFX1* BGCNP6 KQD<AW>H[=%>78Z"Q4L 
@VP1X?E>RPLLXAK$]]S0I*F_7^2_63.%D-$#L55>V)X( 
@<D!%*/I]?9UEMGA7FKHXB(Z33[1,^NKN/7)VYCS:8PX 
@W[W.KB]4[LS6?;?'^<8,?Z,-S'$VQP,)($ZA0/'@VAD 
@F>^44@CT6YRY5F'K4DU9/=0B%MN6W_Y!QI)<:2&!9&$ 
@>T%.09P[>B[VQ<"A)YQ[*YDS\.V?Q18X^D <6M$;/(@ 
@#[D?0.P[WPL:5D/&ZTY8Z9;1DSYF:5;9C#-W2=:W#U\ 
@GHI1NF$*/N10C1Z*HU*2 ,A V+BW)+'(=OPTR0:&J5( 
@<&S.OR] \V44'1J9&_.QSM][H]>N6#(O#A-Y8&W'FY4 
@\K7YC$*/W$!+6IU-.?BW6#MH,=82;=W4'\JY[Y<8XF  
@#YQ_X2)A?TGE'MV5<K_#,3\[CA% 7] >K,7;NQ&NE6, 
@_E+%( 7I=JN),S-1.Y8VTHN<Z O5>TCT7NHL#I+8EG  
@4V%'1;\B,_MUM0__!QV_-!@T7?E8:93J+UF;F/@6K^@ 
@%:D9%"M!EFTG\7\0R'T&B#R1RZVTD%]. WUF]< ]$.P 
@![GUO=!@B+Z.E91R]1^E.>N*J:[.$H--"Q:\PK'(F%< 
@];N;6G'U;U,445S."RM,N]>Y1#S0U)2FL:O:R1C!8GH 
@DVC')M=M#D4/Q.PHWF)?+7>I'D;1&?Q9DR6']@<MRAT 
@*$Q'6#1Q)+OF6>#K6>-FY(C7R28I)+L!)SW)SE^*#1< 
@)M<4-%!?8"+_$Y -G<CSV#7"RY?[C8.19[Y_R/$)V!T 
@!:MF-5I9'SP<**OSN4K.O*6-7F@89?,TZN^IH-08NX< 
@/J\3\2/2+51D<J04;+@DRSK5[K,6[WB:IL^):;A)6K, 
@=Z,B-SY(]!G+-#)LANAC980QGVH/]+,NSE),YH%W3DT 
@NQKIW_UQ65+(BP$6F+J);#IJ62_&T_=.Y2?G,JK+CG( 
@-D$/(C_!&3<C7Y>KD6Q@::Z91-' .@!+L:(-$DZ/D+P 
@DB?Q_G0=E8PZ:&T%4XUCA.-/OWC:LW*@0(7PQE,\B+< 
@UQGCL_BDW.UIL65C.LAL7-B#X.NTC TX7U4J];3TAE< 
@8 1P?UP%%0'!$!O'I$KYA'A.SLD*TF2UY<O\1Q[P=/8 
@/S4(0:.[M8IGT?]S]P^BY'TC>_XJ&WRJYOC<%33^*U< 
@H;8U& H-*JF!SD*$,P<%VFO<X@]1>.QC;3319K!Y(YX 
@Q)7[1EC@/J_S\N'I=&I)LSJ*<8?*\_A^=*PU.*>V1=, 
@AXL'K_=DQ<$]70/2;'O2!N$,)ZXOU07Q6$SR,]\_PM< 
@W7%R^$;#QWTB-LYASX^&M.Q ^=+!?F<#6/Y2D6=!J:4 
@TG[T+LOF)/M@7\RFA1OJ]8'<E[;7[ZQ+NNOHX##OH<@ 
@RX0 Z;9 8/_QH>\#H?,K0Z[M" Z6;?YVZ@K]!*FK8(< 
@:J.-K#\BW#PJ!_W-E)N1$MYS40#<*JXXN+*"6/CJ6/@ 
@9!L^494XKO AA.VB$/DA8V;)'/E($VF&)=BT/5C> F8 
@;.%3FY:SZ$7PAA^KR<?T/,#ANH>8I@4H#B@GGS (G $ 
@]8"Y 8<IO%95'(-83_G?3[P4H)CYQY-XSR7F4+/ *\, 
@R[3E2O6FOS1WZ8S[ZJ"[-8BW7_XJ,-4!H"&8X7,4E8< 
@?Y32WK?0+=H8]G73/9<H>3]8NC@XJC-SC4 ^ZX$O@HL 
@ML@D",'%XNQ(\QLYS;"\B^$"<Y2H?EMY!R*%;0%A5Y( 
@J6&N^Z7SU?*:LN(B<S?V]Q()@6BM4&C!I_?S#[U*FH< 
@*TH_G:;#R*Z9U@\K_5XO,<$J=W%R(1-O?XK+UYA6?XX 
@!Y[_$&*E;QD2!!==!.Y=9RYG<"Q*'8 EZ^56R/89#EX 
@-3=W0:;A64^#&;_T]#>>TNX@-(Y. %F' R =3 ">HQT 
@Q2+P)[!0759UF+(A0/8!7\WX/3SV45EF IL=]68&2$\ 
@=&E7K=88H$&_0Z#>G:R5%"[Q'(4HM@N&*U;[.Z1$UP0 
@K!GYW9.7CUPQ"P?LHZ3B;=?]1[D#7%8PIA5$PQ?(*2( 
@@QH" $MSMO:9%J1URC.YX9F0/?D;2&AO1>,X1'?J 3D 
@!G&=ZXB#SX$<)LCU!V 3,1O$5S38BC8FDOUN&_2%%60 
@+-_!3Q$<E#=5TQ;=<';6DT/RAYUTA2F@,<[)E-R'%@D 
@# G4VM'L/[$J7MQ2@#8"86]UP/FD,S(^JW$VZEV)*YH 
@,Z-G'@ EKHW!EF\2)S[R2=Z">9'+(D&Q5B\#_3-82:X 
@;3E?A:-&K].GH],,^L ,A3WL536+01 TNQ6*Q.8\DB4 
@EA<1I:1QN7\93H"%[(Y(JZ>\9M>SJ^-X! 7\HY1$Q4L 
@)$&I*2*8],J.EIA#^(W"0G,"+5AQ'>@RD+%5%;QR4T( 
@90PMMKV4><I#98XTQB#%,6<\U5YE5)9]NN]>SBS#YE$ 
@^972W[B#=,$I@!2KAC,]XKJTA"CL@.NP\3SX;>9ES\@ 
@<R.[ ?1) EW8&$8?PE&.6')H,E0L>?8.3$X3A2QSW7@ 
0!OP6L@J2S)H5.%3YU=DE(0  
0,[.@C9#:D$KR/?LG6.\2A@  
`pragma protect end_protected
