// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BnYz9RU3z5ZzbluGFeMuLFwkJfkQQjjNInH7tgx0AcyMnpeH3JW7XprgwYAUaXMk
wxVebYsKfsq0nDs7IXSa700GP3waRqyypwbBY3yr3sEgb1SA/rrLlN6FvVj0oCWM
UyIroTeClI2pDmnhxBUccAxJFAyxIlab+MgRTa2a4/4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5504)
OjnxfSFbUPICtj6S11Go5MI/tpKi/PxnF58J4n8GgnHodkJYMdVdCK7FPXoSEFLT
ZuQGz8LHJM8cAm5Uo4YgVcnQWw+Up0RiwRBPijG8RXK3xDgC5iPEQAoFqOytuqss
xLXp7vhv7d3KD2Kt5+lB3ol9DvBwownp5yzfxtSBVPdydiMrTmIqhfxIKVeKhbZa
obLpgch5y+LZelPgwZUa0NYbAyGR/VXbREoD6LbhqlgBhcHnVpQYOy2/fOBdYmn3
EmL5HAGusd4ZxUPsa0YwITtw1owxrX1DnmC7QUyOSNYhc6SPDoOvu6qm86xNGZrr
0q8uAzoef9lqPSL7vslZcHrbjghq+HjcvIOhE72O6k7iAj2394hbEHsKcjugUQKH
9P09JxCoAc7cp9onM8c5XPf5/nMVQSUntbT9y6c2b2Tro+YWzPuT329v+ftOTLUd
wUZ9UC36oszqZkJxJICYzY90r60SZeXmUMlyY+U2srFxd5DQO0EjNeeskQceaiXN
mQMeGK7U1SH/muzQBTuIan/8mRmTk1N4a4KJoF2E00jkZgPgHmGOcdt8uZuAA4XR
Ix/E9gVvCzab3XZnoANT0QNZx1qFzQSLipTGd8/UiSRrINj7Jk+FSv3eLpNr6Cb1
RpJ+5WL2GwlCjLxGf+7fFismI7oZ0xJ1pc2NZgvue8uyJIghefBM53Oeo86RZMaq
BYSiH7CW2ydJcAAbSD2qI9QqiQPKfeyKPy9Q8f3nhCUK6QwPQ6h+DekwJhugtR5a
PRjst8ix0CUeFN2zBX4zBnwtOvcXNIo/k51YIoa73lJdtBr2CZYgO2GQLk9GiEt4
Y4dhzUhqj50Q+YQxjtygt/H37mH7npM6os4Zdkhbw2IkqIJcz4S5GMUwDSxiugH7
6RqDKmNzbwlwmT0HyMUg/giPqR318OzTVfYBV6LQaQgpyJmrVTF1JsrsUSbD80KH
oaCXhyCD2ugm0ANcCxe9GMeszAspVCJb43PEwDtRGdwvyGUiSJyVcY+1Weh/+Mru
eb1Qdy1F1HSGWv26Px9ns6WhCf1DCB+pLOfC5zgPfBHe+Vqe2IeTn+J5ERu3JI6N
LEx3heql4X0zkJkyAq/SQC3k70V2JsKKX4QiEAhflb38o5n09vTsaMM4RiTRSWVi
vYjz0p+c4x1hvzFNsIbZGbHKpvDGU4ogt4ZBh9fpNrX/TeWozheyYEweJQlvmzn9
E2KkvA2l8OVUIF1ZqBDM1ryDVP5xb6QYnpyTsOIzaOiQNFLCmWQYXbaVlOGV3Wks
UzWauxN6d71054F5cHEwqrafJlLCTkLWGyftyHCqDHCJg8XCYMHoiMnoP43st8ue
e8wpO7njCBcuE4opJYTwoS1ZIDa2bPqxZ8OxLromqvL5zkzWRjQMWzV3lCDtSGQM
2DxgUtKS6zWxYZEtn/ZJVL78Ky77yH1yHN2h1ljCrPak3ewTWzc/vONaD1gZXCd9
C6bWhAmxOIE7bTmzMRbboHLmx0AafKtxr1QfjbNzp3xbX5YP0ZeGpcS9Xr0l3iSN
IIExI3SpS34FkPzA6FaZlzffNFLP8ndjKQqTjZiXBfskeJDA4cg4LJSHWkjTjoog
quDQQLaKOzbdbDGJaWZh8RgWiIwdzRS/5RHHhwFOdgaDgT3fcsPKgM8qfpB6Lcy9
/T7ZsGzAZzBYr+9kmBW3Kw5le4qorG+jktGAT/VnHelVGb95xE5S1P0NR9LdWMnQ
rcKlbxYWhLbFuQi/MRFW0lf04fT0rehOI/+6ktAHIDwdDRWnChVLTiwEffmpI5Cg
BYlEIIgmIhWBgJjr/2sC4DWEAuqj5x6VaPXLyS9SQg4HF9WbQ+fMYzvWiptkr7dQ
P2BKoWV+MaA3IiCeziIIdaYZkJ+MzoppdZTK0TKl9D9em/XdOXCJBRo/TdQRweXM
GiN7E36rBUbkYCsdtJ+qqQFscyo4QxTskwjfaFK4bPW6rot6ZsQHL8eH5KAxxdId
fMoF+IToWk8/w9iO1g5kBD95WlUHgYk86KRxRcmK7sRfwgiBZHBBy3QiUrdAeHDx
mPYTN0B3yn6l/A3yWkEWtBuql/PrIUCXD9oJoYizWWoJHhUQndBAWVIgVBUoZYnD
YpA2CV4S1pt9PAuM3W+p1WLdIEAdVH1ZB5hVKT6hYhPsr4KFfhpuivQV+qveVRH4
vNF2oJ12JdVv25P+QeGIeXEGLa//KM/MfmX6L6dScx9EK3D9Glg7LfG9lB2ocz/i
UvN5EV4chxPDUStbsa6a5eDhpb7IqhofkhEuu7x4NamTZxoI7y07+btAOVHlrEiD
gz845FzvZtMosO6zinknYr95Tl056ZrAqMBmrFRu0NnH3hq/TjIozLJxjUOpbxud
YLtsq3nZPUAtygXmXRurpr+SuFr5L1on6W2JHuPtZS3GzQjRZ3ok0my1tQYBahco
cydqGLAe8tQon+zAGqQhafHaIHcWKteGhuPc2/8VoYZ3tphZqDLXeWxjgc75zzgz
rsJsrGIsaZkhhW5HNKdf7bp89fJRx1sPrjLmitf9izGPbR0Pjr2LxYVG9UegxP8M
6mafQnVKt1JYBiq1qaZEAm5ZcsD0QI77DUO0MSA9qM/8DuhaJq8LC1TByd5H9MiA
Q0+NjyBtVn6nrhliBErmWBNFvmS0HSbMenoooS690KhSAcxsMtZtNB81XF0Expij
USbVtlMKs2Co/8J4sFGwBiGdMqpodrjIzhADUv3B+9gfAWOMVreaZoScCv/Jk5t7
HM6im365Q57jUv+u4JsivpP7Gxn6+0s3rxe169hIBPzqtOEoeAEyn7PMydWVowMM
MU4VC6Mlj5xFzvCsy0s03HObMxHciYhCJ7YI9XeVgqYRB8/KlIpmFb01EoWk5DDp
8INqCcLLfYsxLx8gGC+Io548c9tJJBy7jNhDXM+TysdlObbI9M7b43l+kOq+B0dN
PQx/sAPI1f1o1ojTzZIegmWXBYRxJscoGK2Xk0EE9p+vqHC7TUvtzL9wmCYdOf98
XlETFA6IvDgcTeqqh2jeDxjY/LuOmd24d4Hc4T0k/9uDoS51XGA8kmyObaMBy9vi
3FElp9aBuMLO3WAVR9c5pmbVRVR3+RkfIUAQRh+tg/n+a524QnraucT1h1x3wsU3
paXUoWE1my0FH016cmoqjuuR/vWIjRFHoFvqDkYT+vsM2rq5w9vInp8iQcE9FlZX
O3pXvj3sNAIQlJsDUsVqMbohjI+IkQKqooFSCWj72phOFU6UMyn8xnMa/LavcVKI
4xWzsdZ/XHfkAWnejkV1g3VY+Z5FJZGT8NZS8Gqcp644BEzhRB49yBi96JH8/1as
G+/ONihwc2lnWxtrXRj5pKTy/uioa6u5NojyCR8GE2TWp7LI+BYepiid+xJMCZgC
oFlIBIdSbEu3tv+9oWDwj/0PTTu5GMT8o0UOieSv6uWnpOWgJEoy+FwxriFme1G4
Y4Pzw2ZJiUF+9qBuie6/tCu1dxT/5Prj+FKoku5z5JpI0TeRnVrXpj7XLBxNN5Zf
0xuE1qkdoCrBG2b4M8dZObLDU8quu0M5n+olDYbnFlkk6yMbxgghtk2p2wp3OhTw
vrXT2ntG69CR0MFPFVfiKk7sN9vaceeq//a4Vf/EoNaw+LNPMkcpX3CysGPgQs1Q
imXoBmsl4BSzDmN7NzhcrbrP6rBBngxBrixqPwlWJ4FVm6x2MRSq3D2nGGrypdfT
ZNNpqgtZUL4PmO2tHpMiyk+XAhOWXtAE6kkZ5F4Xauaqafd4sQyvS4TUw8oB5Ph3
j4M6dkOj+N+8bJ+YjkiG7p/e4tz+P01SsRFIVB3j+wyVt4JgPj2oC27AM04IqUwv
xH7GRUsxFIWiEj0JerqZS2joR0mYbpQf/Xmwhv6wfiSiqX2QSIPP1leVIthmcuuc
R2Hf1IKR5riF2pn6xvPfP7W44IW9MSso9EG6HkRRHNbrs8n8/px/DwqGKkR50hVK
q9UCvaXLoS8ht1t/8YXI3jMfOELiJyn8afNb0Y0hrCSbpZNN3lBRIm72jkdHKtUr
5OaMXXL6e1mBmDz7nuXKSHDYr3nayqOuPMmejOaGthSO6X4yC+14GVjjQzLfVNUq
Ar2MBzdWZMhzfH7LJ5RqL64li4kDSXqMGD97Um4bm2cA6AODzAwWEU5IOanuAJn1
xAX+WvLZWIxdJyV74D/kp3BPTkNlGL5lEtyt53t/El5tBTRP+cO1gvQDh/De7Zf2
DjJbSvudbFpmr/2NNx1p1LSXW4tJn4QZ7edpkPncJ4/ONAA16e+G1V/ZwsI/OUsT
fqnJwUsKAFWf30XVN8yrjZmBj1TTdcbEhXMSC0kDHnpDrcIuqJ22MynodQowx3y6
yIOT3ZiuXe03fR5bbqlEdAGYgF+pz6fAHuRo9rmALsIewAqDCjNiZF6Hz7vfontz
Cob6CAfcazkFfyD4Hizsd/2/jKjB1nCbURVa5+oipbLMxOXRH6BHXbDBjWpr/JNG
LIHgXMo7uuvY7C/Dfy8eeL4YeejQE7gRVQ4uiD83WjzyGR2XwVu5UnZgsdQXptJQ
8M8hw+EWXNBNj1nBkk7/Dfk0sp9VBRyo9sJStLBM9LnW4k2uy9RLRjyE1Gvys9cl
o83Snxkyrdlx5DwvCLZyd1/ZZvIwLYy49ujOzgymn8VXU0S3AhMldfSOuul2pDy+
E0H6PgDWbz8O70pIL6HnOdySYpdS1XD/WFkgwC1JWYnZyzprXp7OwmnbMLwc5CC1
gZ2jaaj9qzEx+8jcdtjoTf6O+aM+Eg1Ma37yDaKFi5yqAztDmiiE7U+bvQB2mFgQ
4Hd7NtxPNIbXx3JqNXl74gZS9/UuTX687gvR+DdLBPn51oPeYQ23JTKmtZL9FHq7
aeRj+JZ+53Ah1y9WW6M59fQXcnF806uXC5gYIaSCG6H7L5QIoA50fLGZZwkMHxeb
gREbaWWCtNOCZISllWdCVmwuxKEdf9yHjqjyxyLt2rI2+kaL6iiR1F/18LxIf+N/
NVNfesJZnmx+1R2vzrew+JlyoAt5OUKcyOBxJDCv6b7FmIgoYAhdOi25i88beITG
OvPTbWho4hbCCvOAuwoWZOlsbrn0x3pABJ9iv1xemsyjaQhcaP5UpMgMqkD3y7VF
c5m8V7z+bsx7C8KSh/jGA8xRv6WK11ld39osvFyVgu9pkvZoV+ShV15jx+xQ+beB
82NpAeZpJ1X/cwP0F8aJETaBEGoB54h/vw4ES8dBeqnvJvemWY4QuMGISrKS+hvE
Ii4WjNx+/wiWXc35OwzjXLgJdzeYnBs8D/s4I5sBq9Xda1hh7BUCo19M9bCwa3rX
xkHfevsZinqhXuu+4wTQ9ifrDD8l/csAWdxT7pJeOF8FdfXHMvnYSPU94QdO1w4k
JBkUs0SOJnhRCpkcqhqikpAvF0yH8FFMjWqpO2oGpMGlZpaQy/BQqlhWsl86zQzs
IQf4Ki/GHext8avSe++Ehcnix/7OMCbkZ23tdS/sNjd1E/Ntfz5yZq5EYEMqjXJw
Yjic8OmuDeJ0Zd+nTvFOC5T1TyyXd0G0mhADJJKrh/v51RRdHDzys6vJWt6eFNvi
sGo1tQdEO5UhZv39H+4kHVhTVi2l8o/ZVR0a5tIvYzdt7JQBAfDtAoXLU90qCcFs
svcOJrWIrckWDQRpWO/bSGhRQanE1+FThGIpp4Jth2r4rEvaMY38dZmjxL3CiRf/
jbGdkXo4Ntyz3rdklsw8YX+k00ITSI9usXDW+1SqiwqGzPD4Q4Isyj/T//AuPilY
w1lPrIGxvm7SCuow8pSMMOhU65VscHCaRKvLrwRMLWXFlsLRiCvkw0MZq27xkz23
OvvL8o5wI9I0mm3Wg7+kVNLLSeKJ0f1yCfN+gYSghPaplnAb44GFDT+IPqfBqXNx
2Lj7BJWge8bKq5hKGTUPBHXSbp9/H35EwK58tc5N7XLiaBxGWFiEn5q2Vi6Qpe1K
g0UU/Yv+zjkoekOVSYLO1Eas57rtbDm1dgaF0epMhpBJLmAwluStMoKJndG8nSDk
3u37ugT7wVHLnnAYkwp9Oy+/e9mmrt7Smp1rP/T81lrHbAGRCIEnDwpJtv9XC8YN
Vl09WR4XMyJ88QRq0lZV3OCcSyLBpqmrThhFkfAxzAOqj+SxEhEFHujxvB1fb+Wt
o65d7I/xgQUL8/jCk8G7trYukBko5kmXMj9I44s7S2EZWGwajpoVG2xmZVP+3Hnk
TpzB+RcvsZ0q1+Jt/T1JsLa0LbEIlRGjAIGJ5H/zoLK1sTaaGdVlu2RSIyBGEzVg
enYh3QS+ouhvUbTEkItyGaA3q/Lu+t35krZumNcg5O6De43vYrlqskmDEWFO4BJR
GEJ+EA1/0RLRTUtVu20f7qwRhL0GS+z+GRLuzb4PzDFxUvLtnSoqdIE+Emy9jLjD
TIGP9zOcAEgzptwU8hw9SwuvvCiZShJMYlQWstLoRG6WAg59UKEb6vX+dy2TnPM9
xoGITmYaQIOL/Ljdd2bAdytt3eBI4xLMTj9SPdrH9kCUOuWwIzbG2nGaxxpkfqqn
gGr/1I4oAdXPUFgtHmdep05TlcHxJcBCl9kntw7sXqsGSxb1jxCuDPQgj3h+PO4y
1WTYs14i8Agzhmhg2CNswLcxCXQyBHIeQXbTfe9XAljogFVpQOdHMopXJF39pSjB
E+WIs8TWNHwjOqss4bvXuJWizvv+jbn2f+6fUjJx/fYMwjWTfx039D/4qIpqCdtT
XBjgU4mRZCWEr3he9usMQUmuRKmeR/SQ32SOJhbZTVVPKgeityNxl6RoG0Y0AW4Z
9TwOitCo61BrkhnqhwjSt05cavR2s74ew00IDK4TK6CLilKL5R5OeTbpEwlcRsNL
wE2I4Gy0fK2ThJCdZ1yNEvAstbXpGLWQSsUaym85B8r37KNksDdWTGgSko5kd4AB
uzSKbCvDWHY0wfSGW5WHKjDfuPF2StM3gCMldNhLhOW66+o3oWHHiA45fKaMZ9tU
FH+ww4awdILvQsf9NFfASoXIOuqw7grGX3G3kNoK6ofOKHlCx2oopBfCeR81gwgu
FQTu8ipNp5JgEdUDxYLWV/fE7pO+bgGicD3HqvnaYSaWbDEpgwquGgFtDX6zFryw
bE+eD0PwOpRpuM4AhgWk8i1lNir1wSuKSeeDOXlQAYoDe8CxX6EfqcroEaHfOmjD
ukpvowKZgGKx5AUvHcB11B4ZviNMbDM3VN4OgyzYNe4Vi67sbO4w2rmJP4ic+2Py
QYTLIw+bK7L32cm/TVeZFDHUw6NM4VxpUNUhJ9okdQ+qMOaEnHi7FVL49KCa7/cn
QjnXLXsxmoasRnJXuisjvTIa3MDuIhwNBXjrcmlIRe8=
`pragma protect end_protected
