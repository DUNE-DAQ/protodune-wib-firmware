// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aIBCSxetYUXwEaSiVkQJVemC4To8kdp4fdPlgzs/aKMWpqaCLN7u9T38l3+/UkW3
z95mmZByy9PgAUw4AJSPcwiDXsYExD1voZVPmF5ndGcw373TgFVR97mrHkEg6HHW
hF5cFKETERnjN0FbAv/NJsC8y6hBEya83v3AYlpsIH4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27600)
8JI3O0avcJe142pSNMSKG488nus5DF3RicL/LoBPIUPuDV1STdA/qrG8qbgKyzmy
Pw2n24aJCB4PwJdLrYfXVlU5DyTFPAhX17x1ewS6f1Idi1QdztwD79mkwP89X72c
LYl0MrlJyfuPnO031C390ld3fhVpG7TnD96HSY24QtP8oizXxKf1boaDs07a4hNC
o9LIFjx59ojRpKgcR1BBzAKy3XndOq8eWwhroJGiMPNF2LjhgZj6ggH/6/uVMrUo
XuMukQxA9J41HzJX+RpNWpCYhFNDK0qzhug4eeRMLrqv5fOcg1SIjDuYoJTDOa/z
OHRStzS16La7soJV1pcxnD1+ZSXOcY9GY+ibdO90kxjbeH9GF+yfY6stHJppL+pJ
jFLm18yYQSbUS5adgDL2KWCdInkT1wsTbsZqocMLUSz6m7TauHpTQy1x3rLhTqDd
Q5i1d391pfVNVHPzpk0YJ+Q8OVj4Xaiq+xhK9hrNsTMB8RR1/tv/Xw7W1DPp67o9
Awc80WYkF2fIw60F71osTxc48nvad5TWVW0xvSJsrPops0ZpUKWNS4LXRFeAM3o1
08EkZT+zSd6uflGNzzaI/+iiFVLcvZzIUfBS0Z4kloJwP5XEaudcGYSIKENdKJ7G
o3fgxtg9xhr5dqZs3j/WvTqGzF0eFureEXJQofE4bnL8F5cHWB9WozGk9CIKsiTQ
FkL3uPFXJbI8u9q9zZaxVWcmFINjfxWoO1j26bMtIcwNQCxfiP2x45+sMyWVgE2I
1f7TP3vUxJGrxfb3/Wf/555rq3TM8Ru228Iu3KNB4rlAO56jHal6L+J4dI/IP4Ze
Pa0DkcCLD4sTUeUwtd89OFvR0+/52MXbegNBpr07+KX8cKcKaHIpr8mNMV4paW22
2jc8M09AsjSzUDy+hZuPFeirq2Nbz6fSPXQz3GIhHUeQ0h6NhoCuiboy64KasEYm
CeDxTlrVvPPzwrnTxhv5PoCZq5FDJcryNMc/b1p+jbAfBGnCJ20XVWwmN63W966F
29WEFvZ+i1msvEzpRqNIoaAnYkxEnrqL3FPUy7mdADSAw4RvJoSWIWHvrqvUYk8i
ylNHbIge+aYUigo1KdIMSbqo75VcHJzbTfhA9FC/1/JSQxC4pNkx0kr9vO/2WzVz
/OHIroNibCSkG1yFe7Z6iIi9/4Kc3ImMiWr3+H8rk3bgVPUjTJKUA6prSV/0TDu8
hXLecCaFoGJsFzs/KvxSyJ0tRnfTgeRxaq7iohhMdM7YbNJejBdRxmgSUboiIrzR
fE1OUSylLYxDJhQ4lH9hILpIkxo199rLECY84AKrt2WA4Vz1aKcIkMV1M8fXTBRi
2f+9h2eU0DOiKwreeBH69D+PD5QF8k8iKLtfLMhY5UNy6V/I4fzGlHPutzn0r2d1
TmLyqt1XrQqBq1LSjYCHWxsYcQGV9Wh3hlFzLMEpkPzBwsO4Sf83r6qTLpF533BN
OGWWvjQ9KZ8g6JI4uf/hXAELicXrgJ+L+C0DUB8ryfW28KndzoqScULsNt5Hz+MD
wy8mI6D+vU/PmOLVqrKZUUmLRe1QaIEAZfUBiyWfOB4jEDvcVH61wGBC1ebvGu6x
PZwqBVHgTaOfI1s9C9TVXBaZZwsMyn1yoh7Z1VWmhiPFImQWyC9xECaZhhQdp0KV
/mWA2XbNZw+oSqW6UU3yEXdGY8HZ49sXKEcoNhT3SU+3QsgHEQklegMSTVgh+Za3
8G7sh/4A/c9y3Awd65dwVxawzL6niLh8eRTb6LLOCKdQqxiwzcmbNEjCWY90nKSz
wkjmZMepdQ1Mtd1vLh9tXR1pKNRE53hMQcTb0q8KgUWaeRzFkz1QHY7YAz8cVLLI
nq5h8srXkcUO6otxL4nUY0lvQMDE1XHoDjNm/9Zk5xnEXFhNt1Ovx7rLj/0CZtgm
n2wZhaTBJVjP2I5tqH792a1HfGIxIcWO4j3WABZTQACQx0grCfYjSBfmgGZqOfrs
l5A/+SoAuEjrL1iz2PNzVIc5CiVUQIhq2sN8cFTEKubL0My2ZMB0bDoiwKe+3aZ4
nPZN/Rg5VjlSoSaZ42pfpwHRJY+aXHEMc9NLbVMs7yHdn4lqgAPWZt96TJOwtlvp
SrirOjL3ewOl4+3wiS/O5bUe0ifgonB1jcgg3XhsawGKF13yInHRGYoFhlpf4GRC
6C/S7FJVdn1x4q0j7y0ZEWdyrQPmVRkib8YceaHl3iw9TNPnfP6XE+6Tq8xI2ZbX
U/FW3cd+3zI0bmA6JUazoPK1vsatfyfeE8BzyB3/UMk0KdMJXiW0nDmYsluYCck2
ogkh0bvjSXvVJqH2H7czlgP2Prcy4Zno6BQi7BmqTpabzGcuNKyXCNfqmOWwxxeD
KdUasagmr+UbOACxIxL/Rbf+IEYPPwVz38tbyWn0H4BOGP2BEVvrfjklyzO7h1KK
UiFsp2Fu9Q9K/wa4b6FZ2aVDKQk8yVefUL4deuo6bI0GWt1TfectbOV12aEhQuLZ
+MVBphThvZBM1bzkImr0oUmDdauZI0kqIjrXY8TLTh0l0w/8APm4K+UehRzo6zN4
4msx31T6i2tNQxrPYN4JGEXbt4LJmdtKQLC8GUm9Xgton5xFQCPeSvmxMWYT7Xhr
p1ax0oLGiYJGZOTDV7edcmCawHJ99Hco9XKQzeDieSwgDxKKIdeZugzY2RiGRaHM
4W3YMxU0F0F7jtMpJzEk6SZSnpXqQjTi7xTmPFCv538uSrO4MVTGiSn+h1pBYX8W
zJeo7xsFzaqpshuxfXcryvZhH8WS5qTYrCOwKbUkJAHJh9tUpO+Sw3CtCWvpQZf4
k+djGg9X9wTgs6EX7t78yU3tZ3sLbY60wdJeJx49j9AMchf+UtF0gJjrMm74YrDe
TBAd6vjaCok+6Ss6dK4V1eANKnpK4vlTcCr6S2zhrZSJdLISyyFvNZV9CVvMKBNo
4+IbgouMMPN1P9JD1MWGso+FYtVkYf80rc5kumq32+Vj+5TTSMmyO+6/Lxlt5efQ
4RN/66qoVWAvVNwSnWJmZ0wui2Mo+1UtS250zQCLk+nP0ERhNy8lk17VqWewWFMo
UGbrvxChVcPxKKmvO209FHKj0tv5sPGnnzqTnOshx4xn6OxbBVYL2uuMcTbk3yB7
DaxS9Nfg+TdBn1mhXx9KYsykh+JSIbjHK6MHf6JfPxTlKq0dV6VpyNVUvt2ydQBq
RLvN25Vj1u8wbCoiSrmAhPTvR7rRRwLJyp9+qqIhmvqyIzXxw7890jbPMWAGwRA1
T7ktm/MagXmyqhzKLGpfq7VqQ8jgAk6YVaIhBg7MHUTwZVTx4pJh2ToEi/xlGCmM
H0t6eL73Ts9+zXiaNIP0+nV7FrGSRb44139s/TXFgjNOupCh3MuHW6s8Qipg2fOd
pNtjTck1tw6d2u1eAbfcFTzNIzhUF8yj8fc4XLYYRv1m1CEc7CRU50xgES7dslYu
TPiscSxfq+j/eavqmgbai05FbCwwWryLe05Z8xvxK8R2iQgvLv3k8w2E/zXwxQD0
XO/ZymPaiCcMaRKOCGujU1NR5efJ5hzh8/Df3ERK6pzJt4OK4Qx2tv8ehSgP1wgD
NVo73NL2JcgiQu5Xrox7toEtYPPeEtHwIHNbUsq95+sW6jcefrvlEDS+yXV4Wdtp
j69soE/ObSWjeN+9mj25hrdmtb7lWh5Twj/u9KUqv5RZ4d+zcUwU1rYH+svdCMuA
2MgUxLuNd9cUfIf7DxRSAXDLkwDz8toR2R1UshO0lVVdKrAWzMOLftZzR3S8u2Nm
nV63jC1kew7GmLmH3cgpt+bVU12TJFNV+FeizFMB86qfN3YlHF5ynE3Glrj1KuBB
PfcLHQUc9ejNu8a6kjFoLcgG0WieWX/ItqcLASesy/8U1C4DaLLKv9zQneqmmqS9
TQMc/9RPacGsckpt582OLmhPtGaHgm9zGBRlLzQCg6RWUPWq7DSJpBWdFpH1zrAO
HyIqN9ARoHzgzSv9vl97hpNyHNg1NRRbbTny+R51qgKmZI5/zbbazt1rVaROnQLm
4E59mmkm8tg+sdA5ZOCJmLGkgXJW4v0kbPyS5rG1qk0nbRAc9U0ApMk/aRBJagHa
ojsHTyhlO4EyqrTk8V++YM3/3lnvCd7XFmBUvsGMg6noRkYpIGvZp1HzxMA6zV4i
rmXDG/eQKZDo5qF6RQ2RG4zt+c+M2EMgywWQI/+G0FiYuvs6LjSzjFoXtrgLVFMQ
DEL4ZDVMlrVMpD+zc2TxRe/MkxZWJ9YY7DojxYWdhbo7etswGfoESmQYfNarstYi
Qoo0PHkMnDBjhBCEVi5qZkh29AFfYkY0sY2KALC6yDldlb8PrFM0FRC54U17GLzV
pnXiLcSUabF2vgfPqwq6Kxw+4rJ3/JaLdQ5t1Qes0xhwZ51T+aXSwdKGNlXGAPNA
kH3MrrrHzBc32lXysyDmsByB+iVZ1qi9oB2ihECmM8ddaQXnawlI4H5JPcbO7573
ruHn9QCh3ehYtipo13uBMZ7QybF+p+DGm8YLZFcUH9dJ5/H9Ry+hWIO9+a3Xaxsh
z3hLEMWRAqiSSMpPg6bqNpI11wzWPH/J8breLn1Xom1S/MX6m8llZsn8bqlEM9LO
Rk/t0Zo+Iti9M12BKxVY/dpJx/tCyHvb1/6aPuubU6DK82XeavENuhEUQx6311ZS
MuwfhlQbYwKPmCj2EbbsmLV5Js/RAPHO6yvbQvLgtGO2N+U/ssARm5YqI9Bp42nt
O4+q4K6uN6slEsTdZwYvcWPwYX3QTVA5MCA2SRiGWH3+xZ3xAOqZwjE7UqOEQVpy
3a0d/Zq3y37c3tpzjtRmc5U9qK84AGRlwV4RCo9HPagKMTpEEX32RJ55jczkgKwR
+6nqHrLcgaOCvI8xEwOMIVvoNWkW9yZBGIgVdxfm26V0F7wBvRJpqEPp8auJRv12
Yf0RjeLtWTU64F0o6LRbuOfNvbREOegycL/bEMMcCIIW4KaDCtfSF/yZw2h5a/d9
xZpz7/a54teWXWDdD96F4RGG7ohmo8xg3+rdGIBYAYKJCyfhPmnZrCOHQvc+4r64
BO3njgvZ0VstLVfN9PVF7UNPIunpYULNf6HfOJWwPLbgUUFuDvHMqrx5F3VqUwrk
9Cc01W71oES386PuE+Qe0+vjAW6Ep4V3qbTsIcvGsNlxdeI1v0vEPavXLUebwFAi
vu6P6fQS3tT7eR/o0vY/69syXeCZ5lNu7W3oOwF2lKDxMZ1W32KrkHxllLzfqzYV
y0IuejWQWJYsyb4dn9lES1l8oqJltAnBkHRsMjdhpo1rj17tL/UuYN5eMEUir4n3
4AWZuv8VXe7Gvaoraab3uKYTsJLgtUy3+HLOCVhvFPQiOIZ4TWVFH+OXcbjDRN3s
21Vt07i2sLne3/FsFONmYN3C8A68t4J9ng89fnwi927YEpUe8zsgjVCEQ5EcSraA
VqJMXUYFUa+EExVUUoBuQ/CJcKz1lKVbRZcSywKQ2FyHk/WW1cNZBeHI8MNaj+Aw
KK+RCq4XOiIFwevMoU3kPbG7fJw1aQldH5svVejqSz4+YiVbWxI8RmDoeGM09MI/
BIoV93QoxSYRJ/il3PksNzSzZ0AFQY8aCgHoiutApV77n7T98Mq0D+hED0/zSIpd
doFN8XrxrtuyLc6dIGrarXqI7l022CbpaPKoiJVFBa+jQHoMv247fNiLbm9dE6La
RwzHtDhBdyQpn/YAV5RzP3wHHTnfoCYvqcjd8flKn5B89xpE9ShoSg5Ye5KeVnpV
QQBTrDXE+ulAkkgT6Xniq8sg6JEEGX3rRq0w31HHikVXoh0Gw8GCboTuEwZwo8oI
b4w2+5ig8uISYIO9U/UJRweBZB07QqG6zpqYWHyWIws5Ea6rK+2CuOQgFQYjQRl4
M44XZ+Z1yRF+wScAhV7enCx5b8g/W6kCkHLzKcRelmfnyNf2CkXG+Bw4DYyWPR3+
GKghiiLXCHrmWSC8MS9ZxcpuMWsOyXH9DqQr+Cahhy7v6CABmhCWGCHxPdCZ+0DJ
RB25jSY1Sh7N1BY2IwfienGxb8yRTAzDS4ZQ6//WHCeGcJpAddb/TvxWv2XquDp7
jT5bP+AqToY0bFXh804lQ+L43/teQOa4ucYSRySHjXgvWALa6ZT8YV8N+8IeU+wo
BKawe1KcPU2pjCfKvSGtKrPS26f8STzuKWaAT1qWqJKeLxBgF+Hl8X3xO1S8zR30
tuM0VYDnf9+y6Hx2f1qMV4qSO5IZL11AiQix42aoCyagJ9N82qYtBKGDF3z8qxQ2
ePdpKA1+XXMEwoeCXXtTy3erYLWHNtPSinh8N9a8jh4s2wwXwcJWwiGTqpC3y2ha
qBo/pyWz9Bpyb3UIfTKivLyBhVueF+dJbN2VNn1REONCaZa0MrT/yNBjXNF3I6PY
xiXvkO7Q3izNAh+weBjqdvjWjqQWq6xhnnlT/g0jiHfHhXSVe4WkJSN4ODzTzjRP
yZVo4D7PG9mM6n79gceN1aPcGxB5XReC1L137e5bl/GUuKla7p6EZJX8uNoTmKOo
EZbNWdamd/ZB4O8KODCUiP8KM0YFmVAbKvz+5MkocRelzdLqt1khYDCTjpqeSbmL
fx3123K14JU7NqIWiyU281WE4aM+dvuU379Ng8QPklenvCFRiOnevxj1CwGFS83x
VcRNTWgWnY2GfqxEjbyPcPPS9MtDDn5exEVrH6R1i1SlszMIDc3I7/72mpHBzdER
oSqAYAhGQ4oivPvxhgaZLzTca2BIfDGAyy2yqutv2kUPJjv1jVyHdb4fVVTHqwwC
lt3mCKixp0qOG8CPg4AwNfXAxXhkmx/zSUjsu2GbiT5eWgnqLqGBf9kU5nLGqkvA
2+rdH0fyEq3YEzkr+4qAlZKyU2wvAJQz6RUyEOaU/rJjZ9MHgvhQjNof9DKqMY3B
F0clBK0b2BEdCUQ7DgrqEhpUwSiU3kekDAFOMtcGekG2ngQrEOP8GQ1tn8Qyq+mB
3BNFr/JF+lLt9g8+wGUROPzy4f/h08SkNvFzFU51hJQqbOs7ViN5pcHwjLV+FeQ9
ajEUvVIfG3Y1m0MnA5yL+SgSvP0xmB2+ciNF7qfHYhJlP3ODod9S/NxR4J9Gu0k7
aMKDEYwexLaURqv1Zz2lD0G0gXHFVFoagQCtEMSJbHJyLrmDaYHO75V2FVNPkGSX
ljjfP8tB07VIOBZeiJuPVMyShi12sqKfBTLWy9xwisQSgSGO3sfpuI8iKuSF81Rm
m0sGZqdeV3C3qiJHxssH2mUsD0KblgQ6OBhHLHZg6DYmPYsi+FRDDK14ZTZo9Q9Q
8raKEcTVNHmqYB9SWzdKc+7TLVlJGL7aUMY40LSCYMNX27M4K8BWADQce5hmmqGc
Gtg6aLgvOJUVllhE/P9X261hwj3EtUwqQbp+DPVaoUThSLH5uR64wXyesBA6Us1H
XUm8oFBbM7PUcMfqMDRG+uvJaQNlX6ov2L32Dic9Oe2SX/PXEpIQ+XneKR+GERPA
XCjbUfCV5hQiIX2MNZclTFG/2fCd8QmB/po/LgcjhUGqDYtomWOeHirZznICycca
ksqYPFN5xfI77fZ6NcZw5+QL4Zx1HFlfMvkw/dQx5ZqcrIPKe+8lvh+dmtaV0Aiz
ADriT4WUP3UygxGwGXMFp/ptOo8gf+JYVjFGcqRVJcglYENVghy/KqtZnx3JB/mu
VZhqge4bkCGuHO60I3U7buzXkmhUqBJMRF9JW1SdaJE80EbJxaFtXWb+ojokhmoR
y0JcjLLKY8YAnimmOLTAl0g67ZOhkCPFR7XOkgvBwcR5Y05JF5qM61uln2Em7ipV
zMtOvNa1CHSvxZYkkdbAJBsoXwRe/YDdZU+HzJS4tbpZx5QYooMNEZ2waT0PS4Eq
F+zq59Ft1g6w/sBvzzjCpheWKPE4qqTSxg2+3OqGTPwd5QGbmWBy+ybbtfDfzgTW
mFoh3n+9DkuAwhfRnyn5tvWtRIsD+6GhtQqaH6tD+JTbg9UEnniUpfSxl/gJcJk/
kieSPJfQzn8Syktic5ze7L6085Wl2B07PxRg+z0PhpgN8RS7dktI+H1+BwboKfkc
788nlnfpWsglXan0NIFFirbnUi7Lp3wEkXU2CRehBy1wyTJPtYrb6aW8eW7Gr4c1
VUB1MXFga7EOJvLQyKfxhOef76ym0CefP6TgB/ay12TgwuJWhvIxAjuxm328MFOd
wjbRt8a/Sk/RvzS68BKNwyTdlgpFGTL8JHXtIOJjiQvFz31FWjANUmTFFQBVCvuA
+lHMD8rH6Botnqhfn4D8OavYPbNMU0VseluQGyrLKZfcFr6jgTcpYoqNo1f1GPHH
3wd5jcQr80PQK6thLmvzS8XPYf9cbqyuo3HwiHSgpaVZVGHXcIU0wLMiSEy5517+
grwO2gZjipEIWreXj7qEZ6gV6ho7EJCP1MpLFmmKvw7LveOuBjyII2i0FKnXutk3
BDTkbGDi2i4tOUvPssqqSnbjq66eQfICpBCwpUT86cT9T4TGg9udRxADjCteMb9Z
FncxWw3PbIjVABoeqgSgWS+cCgVOXOhEI21gFh0dVfvf+GMEOhV/ZW0izJ2LEF1t
RCh5CAv4uVIhousKphcNNONuvQp0S/JKS88Rkpd9AKMwSWHzfSkn2KG2Ef90YM66
fhiZ0oSPHllAtvsnwRQ/0JfL6CgYQ9FtP5ayNDAL3dANSWUyKQtBM3ii0ok6hm4p
B1N2mK0aTALvTtgmnpb0MDOSIRZ/5tSNSDgU7KPpe1e2aKyrJJqcASRH43g4Z71p
/tPjOIpkEbdy8FiX9GUGxi3YEcshUKPv/cGvVrF7fcJ2erZLsnz+YGubOOq3RpFb
dVeX6sAUJuF/7huY7h7jhhc2R8+dAS06ZFVBqNNZaRX9dORRv7SeUCTLSJSDTsQ+
3Y4o85UYdswMQBrARGigytHbt1dgIEIx17zSebvitVdGyjwEEWD1ZVYP8X3kRzDp
6rgQQ6/t6FMwRS77VPtYHcJPGsFM9RhHJuk/m78R6dQNe8JbccX15Qu+XgtWvMdx
4AP+iKW1JrB4UVWx3Jmaj/dC2b19YdyF0qrcI2gE9xUlPAr1Po4roX4qkAHK10cb
wd90UmGulerh+KHr+4Ayu4uS3wQoV7ujt0u8dmKyX6mQ+rdEfekyR6wKZU3M2ekw
xTYnua5leW0oU+HWwM8wEZhSIfTCAiRDZ2vKFWy4cgOeUqLtpIyv4YlVDGxXULq9
BAVcFGBbHck9mNnTYGKMijVRKlUwgjBPr9/TYSpu/+z0at/nJSWHPLWUS6+GikWa
/JG/cdQL9cZHM32ppXXNZoV9w+LfbCT7STO49buoEgKt965WjydMkmO8bbZDwitz
/LrrgVGt+A1fCx4muIeXjKDVo+lWjfFYK7EuwjPOgJPC05Z24Y8i+EwiSO9SsUQc
/3asaN3xl4HnWKk6/xMEcstI3RqIOtRjm6AET7bhqO4z48xPJCfMkvbZJCvfyMie
PvGo8F65Bmlen1fTnGPxhlTXJYWoWeipB0bDPYGu88Z9ISszId+PVugzqn4ZQ+vG
cN+dwcwNgj327BUJcpMv9U9goPe5RE0zhBXeGWnTz1ARw8549p4GLQXr1ZEOOuRi
y4yb8Lof9hwJHQnpK9+i3Pr4hCnk7Dzgss6OJy9yTlbR5BG6TKsLLpRAFsrrMxeL
ywo7sa5c2ejMoCOIj4zu0EcuPLItbFUzS3N62BTANHHo2DV3wRoXQXYTLKKmHDJG
lutEip6kKjB+K6JTeCmoKo3jKj2y3nrtyTuUShVWfhLxT/XkXMp4WUDmOkzwZM0o
gESiVmcNCyRZEE+3Y8OoXtVXsAk7H/tgRDY6viFYyQKy3dhOFhGTQDxLLbzm4kLU
L5pPcox6eJGzOgU16g6srK5zxWxXS4LYGimeiZwMU3vq0depeR5De0y/VgZYGHfA
pkZmxaro4zwVMO0e0+qvLdkKyLKo8q1R/9Rrl3kMUD10GMrw5wOgkJLGMeNdI9H7
2ltLu6IgrcN08Co9zKRQZipX/dW/WwzD7sZOKkgDM2BrF0Ht7tfKZxVQp8sXYquh
N6yC8m3WJaXFzOEy4N8b+qYyPSSHg6mDkidxxSEdkqRDiv4pYeKzDEvT59KUyELx
ocF4QRt2KTlWWjYN4IYH+TKxle5ujAzGvtYpRjQMwLIbZvHa0b2XMUGeM5lo1tDH
fv2L2naAqGEhyynHijYB9I9sVC5UpkCQg6f0Kp8EXsGi7or7XY0S3raVWDcJwKMt
bFWNyyyhlNBpW9FHaCWcYMqSSmjx23olWT5xxaiFHE5+gPDB6RWRBg3gNZ82np1c
IUpgsfbnoI4sUKIi/EceEhjGEh8yfXgN4SDJY9j8B5s8sMsm4uBnFt2xxYbJvRlF
rY/B/D9f8qkgTGluQ38e7N9KsZelVRmKwmq70JeOHBZXMWbD7E/zjBgVgyG8jlRx
xKceKqIpdI9RG92oZ5fW3qHBT5YHUHoeNEjcK3JE1S11tiEsOdT0KZW4lLyDMmwm
U/FsX8k90LH7JOtqo7h0gfqEKkbc1OKxAPFNynOzkzz86EhYnlBbfpND3a+5Bbsp
JxK/AK8HAa9c/obijx8eJXfU7u6y/eLdp2qK9WsbL09b2xQiHDd6rtPTy5lw2S3k
Z6pjm7f8+5x5oYl125gdXuG6U3UQWjgmtdtUr5AjoSAXBjLoFHGq+p/BUCZgWU1S
OyPl0q6XiF2DOjx3jsqEA+D1/hQc77W1Cgr1S6F3Y4d7eVqvrcLw2CKvzRCoweEM
sAZuGDtPD1IvLLUWeWPVpQVjhHxfg4MVJN5JIr3FPadC6txafJR7CyAkKMFtKnIa
0cISIxVfTgwwwNKPFqX8dJAvv0jSTM4A+MKatkQycWT2TrhdGa+ONQidA3rdf1cu
LF5MPcO3/L/jWeLmlzKLwnfbLI6Q/CwZ/xEgWwqj/QJcH+0vuXIS04SvuxyA7C/M
yrgeF9KOzpqoKorsuAMg009H2Uos8IgD9yXyWrjP0tmkhrVEhVuAS8FI+GeZawwW
rycg28PIWZxyTZIJR4qjjDbYaWaZoh0MTdR8Zo8JCZ/MsXP+/P5JXiy4iVwx99S0
wsxnDpbUGXiMTGMLyvjB6ESaCuiZShwNM1xJgEKwC+vHrQ/8F7DkJ9RQREzhw1R0
l3AiI0KXc3+lHn9Ou8MvTxbWWDJtXlfHddlJo0b4kwxZJi5bPZAVSh+bPBLFSUF4
aP3mCHTa9HYKj+MK1mY7zXchIL+m0fcghTlYGQsZjDWaB0PR0+Do5HGUk0uiHz/z
P0zIvoTFsBTbYEcY5oqsxBVBuw9liACLsa+k8ljj/T9gk3E43de2PdiQe5vzkhXx
d/dKrhKIXMhlZ3nIOIGmf7C0f0cMgqdPhrvdLXBpMX6nRjYGl12uUKOUQssOfZ1L
ZdXNwbva66XHXJnmmlSqpx2oIa736INGItQ3BE/BYNWyjFF88+oMPiAUXKTRp3r9
dH8wqU4xRvUbspDQGXJ+lMBKoPwj6tzOdpk7eIy+3CS/6gJSCDhesagQKGLXosr9
lleEqfugrKU37oeJt7juwkAubAofvdeVyOKrcPRR0dZblnAwWXs3u+1YlkOJQdqF
QAu+2u8e/FQ8blB2kp7+Dj0ZwClpqCJ2s+qvJHDKvxuL+rnmuTwXg6igxwWr8qk1
xLJ0DiBldITdzJDrbsU6yR3e7eW7Cm6D/LqoIhJojKCZYPc9CF1Rmop/o+hvU2KN
oQW12llGDXOmw5T5Y8PPFebeSiTXox35vNRpfLNqPfMp8VjUEkRKsAJZyunujJNc
tZhiQxrrIrOTW4zuDQ0Oc9w7ENlkUMXhzdz3y2mjm7CSYisv845lKqEnD9PoIa/2
IrCerGdwXVs/R3er1qdb29MTOwLstVVoI088ouPFRUDAR6+SYr0E9p7B0Ia0yOXG
5tTXJE7q5x5KyBZAurduxKF3dZjTUpXEBgSzEZm+8CD2v17VdsLPQqhJQUs8QFwy
ytMp28H4TXT7AGVSG9AWk4/eQeRdchEguS3jevLEt0LnTTuLSw0VyJyX+LrT6zZt
4nKQM7HL9yhOsfWd59Dp3pcnKdo6A7b0zZp3RX7ZHOl27RxtPszulo+CFGFjhcFk
9nJGgfKo9lTlYaZeOewUIN7Xa1knTppA3d+vTAXWLjGMRkEzZv/qpS2L5mtXByQ5
dg9X6e5BaTmu2JKoAoDJ3riS6H/u7RxpYX0XiDp6or8YvoAVDZ+XVvTttfqJpEvY
tdO5VnXW5eGDN6o+6dtRrsBj9nW4QkXorBLZS6Q9lrPMuLKxjdwTykm8jm2b0zgt
fC2glB07Dz/ahQG08POgAd+mdxhde1JvVVcC56cQYhfuLlwAQphmDJS99GRcFjeJ
DG0eS435OBAW6YdHjTwVxnQZ7nwRQIpjT3dlHy5vbRcnoV+8BrFDBGVKdAF0X4KN
cgkeqOiB5cR6kiH4UMxQHNEYxfKCv0F/7vMJjsn7OHOlt3xXUh/JU0jIV8inmMr6
alkCb7YqoaIuUQ9mC+cqy0LvU8vtHL5MWqNXBtx7kAhGxgRq3SF42p4eX0IWh0r/
rBquI8ww7+IS5IkaMqY8A2+d5InRzgCoZx+PqwZusntJhRkHmmidJy65rpAqGze/
SAejERtSiL4ix4Kmzlh0stx4nFRh2wuCP4c1yrQODpH9/rIFuQLR/da7U4bZ74Yr
VXdFtDCOee3vX4kNTPXVHwwypIDe/lNSZroBGx3ZBkq1o3NdAQTluTMpd0gQyL8y
GbLoK35ltHqpmB0/RcfnqfLe2jWoACCSHVcR861T+dtTxl/5RXwbnp4g8RRPc3U2
IpK9HRYzkVVBf9dBiGHF//BvkQz+I0LlwP3Ed2aEcyXxCTAqLBhMQQeYeY+kaj39
PpPrVaTCX4SuAobQF9UrVZoj93wbOMuR5pkJ2MQ5p7qLXHnR8x4JjvjgJ/kaLMBA
+xTi3Dik9cHj0BrH0mpyWvb+ejTvKJQNjc5/U4Wjnbk+O1vMvl8dwz5JvCnQ4Trh
BSoIAXKSzJ6BNflkBEK5SUBJPmU+NygrhqASOgljUH2SaxTGt7f96NNAehdcb1rd
NZLp5U8n66u6LkzSh0WhYrKH4sbd0YkoJngS3QJpqbll0fQcGj4mo0TD5INJygqx
nhCV716pHFh3/fdyxXgkYbS4w8CcgMXOLfRO86hTk2IXx12kZZf9Qnr1n534i3G4
eujp5OqKfrYh5lhNcKKhvw5LvuEOY0N6iwO8YfCTvVCdUj5cAiai58sHUbF31ghZ
HBmJ1jqMmHX41bK61JBCCF6K+rVe8k1g1AoRvXA1+PSnzqO1FWQroMInAcMo2DMk
8M8DS6VJ6QpKrSbqxwqnBZhghbZ0c/SH2seyHgDRKxXrNDcf81LlqltD8I+K3J1m
mlFZ+kJScHMFD9Ax+MBAYY/WGbe8p81xRZpP6JVfzsLwv1bh/CR9BpVirwr9nGtT
piEbKNBclDHJtU+xe+1mHv1Ap3z+oVRo3wjNr2YfwGUDjeDZvcyHf5TRFKlenh8V
M6cLc5lFcEGYm3gANN2MiZYDjYBDr/C6UbLZLlPNl38w2mHkG082mO0CgzdOP22+
7ii528Ftfjp+/e4jvea07D9z3/Mj+rI0fX33+ISqob0+Rbvn6nkeBftXmpUepwtf
FF7sUmzWo9RS/2zwTvXNvNTzBhfASybT/LOb+3q9CNEPydz+IVG3whKa+JljiPyD
E+hG7yJBm9CAajr6tbTTyKH6xDCXrVN1hm1ppE/0W7JwK5NShUtrxDTtnJTnRJ/e
DbemkycdY3id/bNC8eMQB6Ji3p85tY89XHwxE9bX4xZkvlPotPaastLyyCAXNcWi
ISI7YV0Z4IhvZE2lYT7tvuCvo7XXlreFmsvsCWKzZSBFGRVw2SA6LwCbl8nDfLQf
DvBpyePsrz1AYom06b+x2M0eCLWe6f9j9jq51cjEoiRgtv/MERqujGarg0Qh23Xy
Zw+6sGEC+1QUEofBAMIYuH/jwIYlmkD00e3GM/i4OwgFCE1ovkQY3eudTSTogFYi
qPLr6zbQamV0rgiYMbVcLmovqAOcmkj+B+v78oef7qZHlnUIw66T0e6RL5TPnM/P
MGrP3uvxtH+OvVsbebPn+MfyL1I01VELxv8usKDEaALNEvynEgpChg0c43QLERh6
mJUiub/1mmdDhtLHsPnd6j8X150H13buYtwYPtojANeJ6BBl/s0YzLL55Id+3vpb
FwJDFOV5MSO4pwAaDj2P4rcCkMBfwdIl9N0OjoTo5dy5cezuKtbE0miFKAsJVW9H
dPz8iBTwNoUqnnplFa+rf9Ecahk3Qu4j+x6ITaKI19T1hPrA7gDkwEpz1mX0q77J
0ZwdDxqEV1V2sBL2cQBYEK9pwe7qmQEH82NFBrJpwcSbLRN5uX3L0ehAsHO0MQCD
EHqIAUIB8tyyiQS9FaBlssrYQ3ytnglF4Su2cBOlPwe2+293HDNh9cSNgQYg3Ivw
6h1IEfBJP0r0ovifP3/CgiEcmB8JiePrSpBXeJW15sDPf6PrMF418Z5Ld9Unp0+l
mNUPaf91zAPmHh+F0YUi7+Gu5jIYbFJyroGGnLWiDXl75hkyG74w+DWDXvCcY4Mo
phO3sykK/iIJDEjFYRXJ84mzJ8f0PBfV4mvYWJuD7SmRC41QzDr1I6ub+UqWH1xG
Yaq5Uus/TIkQdppRH95NoYr7F8avq8/RVt/oJB36LFTTx9Mee+qKiAdrk3cZduxm
R/0I4bLWCd2LORgnp1D7MjHtv6/oYztnSq9SuyJxwFaCcd9r/EsnYGgVzdcuc2py
K6dDUD3NVqBSl5xZXhynxK8jmh5Rt/X7WBRhJPrQbDwDRhWH5QcuYZISSePnidXJ
1PpY3IXhtV+7YMMzCaLOif31BklVnLcvHbAhkP+lv5PlVfUIJKIVl0qcfZf5ZJbc
P4LQ5YA6rh/TO9d9IlsXVmgxBsTWZ49hnmiSFBnzJxfq8X6S6vC3sO592i2FEsfR
4FDDPoIok48DTYI+UtH6jHDNnDajnFurW7vmEDNMMliimtrN9tPEAIvkevNjyVrK
Jv7/ZLx2ILnN0+jYm63Pwru9aGhAskuIDHM4rcH/W9Uai+mRj1s76ei3Nn8N/Dj4
vL7Gf/eVbuEXkjEED9cigHZJM4fhpFjxi1kcXv+HQTwOboWiGupaLfptEMiUYBSP
DjDFREOtJ1kz4BHitu06oJJv/HMOA6xtL6wka7GBeeKUlwDQ8h1LqtgOEssH/RJM
P4uJq23sATMLn5FpU1GlbaoykjlI+8+zq4SseHE+zdf5EgCFWUbXLXd8nDWLmQ/o
PpP+HhOudAv9upY0Lt91ezpno6jKFOwR1GO6YY+KtHo62ftvU7VOdRPE4DfBlWif
X56Zn7l4PH//XneQYTfEOMqTn3pt97rQxgnyDswtHsbjTwyeDObRwziOvTvBX1ZR
VIFAJzXYXCsONoQOrCRCQTmI8rcWp20dkeSNk2aqyNJ/4OKt0JAX3RNIKH/ciqDB
tzWSkdC/pOoUPF23Timi1xVKPDqZgnSX6v8z4TMDzg6wZzET2qSk/qcc2WQ0gkLP
DUHyt1d/MeOswO3xFmgvTHWWjTDb0M6AFn15/f7KluG0dUXcyIfPdpjLStFDBTgi
X2Ee217FQF5XodeTYSATYllc46eqPoSIrjgzraFceVbrxPqWfYvROLsl2P+SvToz
bgIefS3q5DPF+65VfCW33LRhN/3ceUusMjXVjJERj2yRr0kkNNqikXrv9FjeuzT0
diiCJ53GTvRVvUcxzXc3xsw07yr5CjJDTW678v5BYM8i44pM19uHPXFnDimWZGAP
qvqJzIiIyFD5vRGu5nUWKmMKGxiM2MMqMMQp2Y0C13/joMrGnfifgOCwIZYOMEHC
m+4EBJawuAKNSmc5w9TGk6Pu9V+O3JBb3/y6dRccNvdZdCnlDXodn6cHbF3KAGR5
67h6tUHeKdnPxqV7lLoS5HtQX8dXCWalOPo8LzMqvLTXUw94EcwEpMF9UaIw6Bz1
sAQALW2gZLl1qcEWjsEVIg+aQpaFAasjdfHDgicXYMpxSliTxw0bZi4iH92Ig7Oi
mJapu0SEBYZg//BkJmdZRS3rNBnAtIybDQ6hVmwSqORzEEveKgiUl9dq2Fg2qjBe
oF9QBYckWdgXANC0+rf1LtgGAQoEoIkcEumiow5kEhkJQ/JbsgCgdurcidDBJUUO
7RxZBDXFrwnPFNSUxHLi7JdMCZeT1A+cpZaxZl0NTN0jH0hkMQpK9K3O7ig3PmIb
yiH2b9Njp3OK/O1/UKgBDdSEKGBXRYoW39kIdlpDCHM3VLGx+6qVIVe0nsaOfC4Y
7IU6h6l29MaEBC+kQU27JSMSjN13Zudb8WyCPisy+/JqhRLT9WMofUV2LiVeYrYe
CsmCWi6sU/HR7ULUm8wC7Cft2gMqNoFmUDCfb/7bvAeoMv4enSMRtAXbgwU3a9D3
HGkmT9HSfj1UeUWYB3C8OEhHgvBLgCxeWKTCCXjLLXOlw3YnwUFVkVCNbP8bfdgO
jDBnxm+S8uqXKtNOnCgjED7+mDnNXF+QMu5zhzZQfxhZkuso7WE0KeGpMpXUPrwB
jNtibp09hHnCOvFUdb3+uRJcMygiLHZlxbe7wYD8jbsPQZLC5lTzRaZS1kBwdI40
AGqfG870MqvvrDHNBOhCOIFks7HToklKxOPB/tmmxOOyWGLwQ1Ya9GqvHi5V4Ftu
lZIegBgL+/REJhugiDNv4ZbrNfqM5D9pO4iG0kCrCIrr7nvtq5aSud35olQorqKQ
mN77tJrxIpcoRQ/0h7/4aWQioKoRPI1NfFAnoP2QksFTtOn3wOcPVPSf5vs+J341
jUTkyc/sOPTCQnq5uPiKlURAXMp9q9/AMOb3a7qjYn/h3wSRQMG/VS43wzFPc5el
qolAvS3AbeWFVPDb10v7/hbg8ssxO5zpk+uhxmrN2rde3K0cmA+D6K17AbzVXUcB
ByLGTtSFrIjUR+jbh2OfBP07YP31cv60OHqXQ6lUwhi7s838Pzu9dUe8s9cVHFgS
sHHMcSZ+Etu7txUqi1PbAlE8pQafkkq1Y8BeWwB1rEFIvVwyfqfiLKEQRTru36de
QOXPTFMtNnEmttv0Fl8gsmktm2WbxZ0+N7UOT/ddEad/VY3kVRlQDZ8US4ozCndF
TiSoTEpePTJC1v3IyNJk6smpSH83GskoMBGZeyQTopERtsslD8yhCxlZcjwzN91Q
I9phFUPpuqunT9P1FR4YjM9EaZ7eIvwOGBdL1VsLGTcbiwpQhnUEntK5mWz3SuX5
BsIzuMdCW/WsPTGQf4soOtl5hIY8e7lbF7G9mCMZbUnwCAmR77YmMxvx7ahH+NdT
CYlZoQAvq5xHkC+hISaR7+6paquhYFFbzSf4ov8RGpoQQT3cEB59rILPlHCTvUkZ
O5NZOY2WweUfuybjuxdDQ0Vt4TY2pbTozA1wIk6WrJh229VXJflCnH6VOcP5Jn2G
7nmKL3ifEixqqP/yvO1ygP/TQRwkrT/oB70y6nwyLnId8pB+dHlkB39bDVSGlNH3
u8/V6+68xOOq9m/dX0uxR9ZVPA+93bY6TOja/jwDZDpuCJY1q14VuCQyavemLEhR
XnwlqQJBgE5jQUBEqT+sKy85mx4XDF+Cb/P9FEX0DlMA8u5FIv/GewFVwweODluB
ftV81cYoJbQ4VY0NkM9yeb3ajXRRHANq32InoorGl+9J35JbSTD0vbfLK6jcHpn3
S0FrE8ubycM+qlfyeCSJVrovlwqd6wKSmLwYrkUGw/SSSFTdJ/kwqAPaoepLlchR
GVocxinNYIuxfmKLXieKNEOR8jr9SbgS1wRgRXxEhFuqqAgKsS8TLDazKLe7C4f0
/f3z4WaGx9MvfGOpk/tE+8nyAknTMDtWBzaqK6WrNJ12xFrenJodLgvOBfUDAXYB
gzodakCwnupUptb2it9A1TMQ8ZV2KzoDCBEf918GwHYfPLuGwOKWbgPmlhgcHNbH
N/AM2+aQl8EVfJG3eP1So6ZhcULSQ2yG+hpnYzkDXfjIX6+gFc3XEEixX4kUirVh
nPY+gWGGfjT/3hj5stkSq3FEiMT/+aVqQzhZWSfo3AYJlvz5AP9AsaZGMNb+qdmn
/qdi6gLR1ORB4YsaucWLr7etRRzEQ+385+gCE8A95E4C9N6sVjSB6CObS34iJdwR
CBKp7IRXJZmUYZbOupsINeKtduzt3RApBt15j6Li8NC5vwV7oom/nB+Gzpi6JCOW
iXilxU050arONOA506K8x3mnSXQ50AKlxbcG5xHJZaaUceNgth6EfjjdNwCkSP4p
P1SSiPSj1Kosrvbk5CeQh5wW6MCAEE6Uk4tK+KoSzXr5CdEnmqv1sYmHdpML485q
TXJEpQZo9FcPy+aZ3hQfxjBD1d0bWZAVLV9/fHdJzanHmP96EolK12z85zz4akDg
fGjOdp50Y9V8CwtWJ2NMv2oysi4UURzv3YrOXwK3GqQqkr9JaRJEEgbdrf/zTZrB
dNrPBf5Petz1xr8nCSvfXTKkDegEkl5vyIJVmqC9rVrsNbwOwhIgTyOZVMDNrz9m
Dg35m9vD8ERR5FwmQTWxCzIjGZn9utajEtx3g1aQ6nya6VUa/2yV8t+4tOZvwOb4
6PSAq/gsWf1a698NGVXVrdwqktqByLyi537qvivEyjVCknBlcije2H/TmmDdzlbD
iZe1GPJLGsZKUfFMk7g3uCHywE1QXnzDUX2c1MbZBDG0cUWy/0TqMRvV18l4K7d0
Lz1VH/vY+XAgAVLKDDMEa94X3U0EZ45J6HUlDfuDZ9pNEWB/jOPsLoJag0fdPWGC
WweoulEut0F05Y+TXXp8CKZmOjTA/Yztqy8FjANC2B7c/3mi1OJMl9PWOXT1XVCc
Rjo6s60fkTlw6+UP5fxGejy9utn6PJ/7Uz4276+byYLhjBB07S0gxs59U0OQZdYk
4zE0NvHJemL7dr5wM9CSbm/UqwyWlM1FZ4mMkX+owNa5DgSszokJUd2uoAakvYJt
kDuAaqghyfT72oDgu3JFoJu7ca8Qh5SrKhj8KpsLBNxYFNlaBjrtgzpY2t0PSLph
AChG+jvicPOI6aFEoO5+klC3Xw4AufQOcUomxvS4PSAcqcF+pjp9QhgVyqiB4Cv8
vVX9V7xHrle1ggFj0FV3LgUjefIfoHog5zkvu4I2mt+M3XsZnIKJK95D3/0m1A6Q
XwtaJq2azKK2W7nC4rLlWAlhbojmZKBkbjngSBPPUcLFFOwUYgwDr2H0FP8kgMIS
0s/E1EYNpt/u3LpQOCcDhXHdoRcy2S8zBjUzV2UIsqmaUzUFMdDXdWRTPeu0xr9N
FPDmjVBRI/m9IOYdUTr/+V9hmttKsHHF5roMW4l7XOxdGPQ+WnLsltUOYDe1kcz9
pzTESuHTVzQNVjJw92ENXY+27hqOx1zfcLMkhdUvf2oZh55tTpZjEKE/IwELZYXy
EaFWnYSGDVvL8UfTzLMPRPdOlE/fxl5XBt+rNdJSKV+cjcp9CW9y+rFAZopWrJCo
9oYLG2iNw74RBhImK10yoopz0v7w7pryBPQJFmePAaz7vrcE6ZG9rdFnOjQGJTmz
VBCVXkok6a6r9Vew2QlTHXHDxGPVKlHHeFPvMNoAzOwFKkHfD6AvulBkFSvTX+Z9
y9GzbpHmXujKPop4Sqtv713pqEpiz1Dzt8xGorawvrX9LzuOwnu9tM2cwfG0gm5i
jOxEpg+gWC0LyMdI7razVHd9vmq3W3+HvjgANqkj9R804RnxxkBUrjP3rJSNZdSr
k0IJaRF6c7/DZQEJHqJKc/IAGINM+pCr6P62eKxpgQmu3g9NfXSWuwzYRrL/WTrE
RQFrbUrovRu1+dkx4ZqzzpEb0OPGQrkbzSaDwAAt3NLA+1QsngHs5Iwu7q5rg9Ge
graC9PjXedYJ7KmxfIov9fYUabzq2E98XdIjPiovcgI8IJJuowTQXreavKnksJNP
jweyaP+PZiTO/e3/CjJ7yTEcUnmITIY5RoXvMFhBstv9pFMgutnDAsf4jzNaDluM
3CXyKcB2ufS0Cwvj54VxSBacyMmRB4ullD2NjhZa7P4uVeOQ2ihG3PBVgkqNpM7J
qFYCNyhFul9fVPiScQnniGTQUVdOcg7U4+F9Cvz+KXtyeEeOMClm6kQO4jBmfMiN
7B8gnrtEot+mYQiSpP/daH9OLzgW9v88P0bHXFXQjDZTjhWkBpVubN2JAKut3hBV
vovEvS4QIc4xA1284Zs2lzlQxGFp1eupV7v8jY0zTiIHaZwuuigLZhK6dOaGqW/N
8n9t32pCdHLzj8/gquHJ4+PHXnTPE81lD6I5oMhGWBSHjcBh7ZC0u4P0iTZ9gGH0
zC2P2CevlvEtE2PBDj7uaEcl05pxGHXhM0OuOR4HKooEVNfFZC1AkNFYcPRLqGtE
3lCWNscifnfjql672bSlusGhzwV8OyICsCFwZM0O2c4+vPg6Ix8Hr+Qp6fbyCsOs
igiU4KNbcabiOco1YTH4ABovuN+7+Mx7obm1OAAh5wPMAh44px2VDjcQmLGriIDZ
GLucDeD4kLksF6YiNgTKU3GZSV2UMMJMADf7zZnHuTkpIrw65VKttim09mOr4qC6
UL+Y48Tw3kKEWhsQDhJ1SZxP+2/EVUusTDO2buFpj1PZlj6+xtBlhd/u6/RvkSj6
PsHeiLiZyvFvdOqf5THXCL1VEkrRNLXMK7Ox0gkWAxonbjvF1WaJQlCObmihYvss
0UEyCB8p8DnaVC1Xdtc7VorO3mPPPIOhphDy7cUypqOEL7+YKn7+2YNxoYSnqO9J
M76z1eZhB24NvS4f9ytH3fGCplJRCS5lR6tothm8Vlo2sTRam6CIsdtyZENQktH1
sSreA2E59l3sQ/L1kY0TX9D3vxCMspy6yPSpipkvhwF6Kg5fWdXquzSvp4YZ1SXP
YuYSD83rWqyQcPrKFuYpvpRBvw2TQQNgq/tt4h250/qi3iWc9XfQdybpaQIcCK6G
G5dOMrdqmqyzgg8+1C+QctUoYra9+gb0VpIxFTkZWz/ckNJyuXRwX8bVYWG+Jfka
iCN1Mox07NCFkaT0Qk8LpYcUU9wDJRE3gSLB/TU738BAm48B0Ww2wp8FvoZuJaTm
U2j56567QNMgnW+W2Fy+wRfCAZx+FZ0tZB7jE1l8h6L1IYX+6aTgT7KiYyZuYV9H
N2uo5UWIosYovYk282tGP6Mzzv0wMsTOBYj9BMIOiWZR3YTPzIrR9RE54xmzjOMc
SCZFhlcLlVk3d40U7/Gu3Lle68/trFoDdhxe/zGvYyu3d7zUhLmkUrMRGBcBLnn/
6q4EcugoRLhGa5Tl1liwr0vv6iU+W8EHnHBXQXWW5p7v85AkM1Gc64osf7WZttSe
pFYqLtKd2ehDn90XaSAFQDkvfMO0HgHNa3jch75lOEtURk6w173bX7nL7rasv7Rq
cdLb2wQHjqCs600SoM++SLQx1auyMA/1fo3wUe/YD/qaUXz/RjNAqlRGUV1pri16
NLaA3sD1K93wlGGestDyUFaT7jiy+iqk7xc9NhpLf4UUC2H/JGr5Rnc2Mdo4RtbS
vJPdu6wMkhxwsPHG7o8AYyIzYQJcouFD4+F1Su66++o8OTwLi9YCr6wMutMRnBD2
0ooNv5g55egxQ/pAhVxIXMlhvgjOfKLB3s55b3urv8qmy/zqWvWU6bWVppsbJr3F
j8olyubTdXFSPc3IsAgYq1hi+w+GyLH4PAkB6At0HFR1ffRsuWyWHzhnn0/C12Bl
xI0nyMCcnGI2FGhPTqBw7PUuLImEY7+KgOxsr1pl41fIOBskgZSqdd8o9ei0Q5vS
Ik2NTX2rEM3dEf0+uCKXc9qzxjMLZu6Xjp1xg7/W4AfTWP/8qMTbVKlfwq5bgPb4
f0mehiwPerLTEDJg+ndtZky3I/OI/p4DcVteOhBm413fnJSGgCmf8TFu6KdzNM9o
Hrs2OBqKkZX08g6Xutthn43ynkhS8dh6Rtob67HPFTsYR0NDj4NHRrzicD5cSf8/
FX23/+RHyDkCx3rqiwzpyUIpCumv4ggYD9RRVLiIrV6YjvJtLeYn0W8qHB6XRa4E
TXBQ0dnIWYNRQdrv9RGAQwL+WAUeo9Ruov+3OzpiP0UV5dQaIngjj3+/Ok0IyQj5
vT4ClJLVDYZ+xOZe/f9v5sJSr3wpOPyhnzjyNk4QyJsfjztcYCRNOb/+8A3/zQAa
OmbcLTlIt1QYYYGl9dkvXg3Di0OiIBmEPH6tVZ/XOIHSjUdusmW3k2B6sdH/v7Ow
+3vvQrwrr4W8O4WHFuqUtCyXH7k1n9o7iF2eu0QUt9+ECm26xW41u9FuNCOF6LZk
GOMJEZTTpem+2q2pnIGoAxb4BVLW+m9eIbviHnBvesXr4WDKGABd583xxAemvtWm
ItjAKzcAt8WCGQtZAH+VxIyA3sr9miYOOzwI14F8PXGpMa/5P+D3f4gaF//gYJfU
JaNVnPqRxp5mwnT7rEPqHCVXlosHCVRJPRrXoXBMTFsH49605bzd5UkiNG3nq9BW
FlKxXMH2dIYrkn3cbSYLRvWRuPP9b/w5oN9XzmI/voKvdTEHYUtFvCrpL/YH9E5h
y5u/jwHzr+9PKPQYqZ3RbiKISLE8Frze9kZKaNJqRZnFQN7xo5JxGquUGvgQA1/W
Ms2pVSj9tZ0+4phqqy52b9FOXe7OPsi5vdOhSuEd/vOUBMch6xM6g4QDykg6lmzM
2tPVbliU4iierbB+5Xuv+tAq5UyVc2VE37JYWQfTwoXahHBTsqLxhKJ5VgqfBeFB
y5mBJZaSUZnTXHZe6FSMWbTzfE3xrfPNJeJvZ7I1tblZxsdzyJzLGUb0bsPh083K
IUGEcZVRUlkLiPKUIVo07fKziSG+s7dpKExkMynzglUb2Zs0zgT9oLuH159c6Rcc
jW9u/V+7PalkKKF3PAL20h9d9Xl+ls7wk3cP8s6FdFUVMDXCiS+2nDb12ZWFyPj8
qWNqoXxFsrrKn1xUI4tHBZ8p/QdlBA29TAxFYggQZL8fXP95nsDBYgHJoII9DOIn
gOY9zsVbAjlqd/6EF7/xK57iHSkZ3omlhDB339/9CDD7aohcjQu5Rp5gKuWBCyPd
INUAwBn7s4q5wqBU76PlesAYO4rRNZAgUEaX0R7m0i/sPUOtpzDgTScMpCLhrJui
cJOebjM1brSBOILR61xQin1Y8a/nsW7t7sbhnBg7pN3pgznnnGEd6gzro0JkFGSM
BidpzsSHSWv97iyX3+VeRDpa/wogB7RYEwgYj03Nri+2s0z1+slvQgNUqf7ZEPgY
+8AqUUq1neFqaRmqq8JrZ2v6Bj9SuNbFAuLKeOoEGU07UwPcEcWLeaOgHXYDFpZs
X6AZ3xxpIo1ITDYs9szmxdwaN/7xvmJ4qV9r+yLmJ3C4nirE6KhpQGx4OJXdUQPW
BiX9wYJaX+HlQdeHE6GJTJbS6shq3IKm8yjjSMAa59Tbnbii+eOir5eJCbt5bXmX
b1irH2wv8we4H/PqUu1g3PmcLSP49CQc490NwoOgv0nabDF6AsQx3QUDf5/FnfVl
suCchmbQ8fLjvYvCA1NNs1xmtfVkFWrAUeXObbsyYOCdUMANzufQ12heyRjY67R/
7/ICZeIvjj1MU333OJbUjYMPr4Y4HcuhmdoUAn9HGf56SS7vQ/XPzlTyb8rGbXh1
Y84u7zBF2J4SunX3RQluCcT+nZ23GVinxJP3dGAm228duHB7GmaDGx7Ez5t6Kuoi
wOTVQABpUOgwCrfI5NSkcNgWr0DqTlcBNWYA2E7Vkn6EdnrWbZY3GLLrmY5q4vBa
u5j8Ci3qkiFY/5HGJy9yvpq79sz80M32dZiaLBpVNEeAKi1mAUo9TLLS7U9kJmHW
qMOI8CTxI09RRAZ7aR+KX8xQvDwL8QpY6gM41H9hE61QYClmfEW2qmDi2247Vv87
fT4NbMwA7j8RTK/eX4o2tnr9jjvD2RUWiXWlIYZPrI0N6lQ2iiSmsg4JoFDSGs5S
MsNxEbjf4W5BFzBmhWucF/8AocVNL3zlE8vMBrJgZSndCs8eLqa27n6RwTkYTJ7h
hkKairY1HYU85CI4u0bBQlyyFUKtyjLrk+mKtYN1n7yy76rG6mxYQM+6lbYxWP23
VX8LBXLrkQDlp4KWvmltX9IKKQYWZitNnODs4M3S039mlr5NUrkCnUzTcgeGUs9O
5IGYn8MEoC8PzvGRrUJnwT3FCLSQmiDhi9gDi86FVZCM+IqazEQlNViPPx28VoWj
mPmjtVX9VQbBEzouUK2DgzzLXnWBPdSpdgullF07uIDwsA8CpgfucyvlvL0QhrOv
2h6gUEBs6VvOkV28YpHfKHY2GG7+QyOz3Z7eUWq48H73yW8qWhBSWRvAKOtQj1PS
CLM40iEPTi0Y8fxmX37DXok0jMXnWOjVyrVK3aIH69PleS9VzS5YxUYVfcGysaNi
GWGffYrepCOhd9kOK2tG5uJtAlM2/t3gnfOWfcQWK4WM0vFPQYtor6Gc5GZIcudC
bhS1gbwRNzPuzdoY2D8JqL/V7bM5FFN3eEK8hGr/O0MuHButeRviLmhyEQUML0Xj
xnCGfoEBkIKPmCR8EkB1WptNNJtAGSIfXaF5cB1vJr+63MNjhD3U0vEQBx9IBns3
AratMkSg5PVoShU4EM3vopey1S6+8EX1vAn1FdYtObTI4AlcpiBvAKda2yVOmcXU
iUlehWifplQoHtn4EQ/vjlOFDkEHrfc1Ik/wlkySVnz1nXn6WcXejbFac3CWZLyv
KbXshf2V3j/9loFks08C95tgc+VVSf7FC/fLHsMQAxIYTBpxak28p6bdFu86Hl8L
pJHLAW41VE1Pvrt96wHH32aiBjv3vxeJjUPnfWdeGLPFfXQwDeVMmlQm8uYcklM/
mSpmX4p7tlQgQUxIzeTfARRvdFOUs9wganzxnNXURgaNIbqlImj00bM8CoDRO68h
rTR1F8sG3jdYDh6bM8D2cRBsYdOuhVIizGYyisUTzVZ5hAYhW85X/Edkpabe2NpQ
Wh6yWnVDHMSfjTM1suPuw6dxp3tkZ/LgyTKx8Bq0+EGcN9kVFdbzY4+xm9+O7EZW
Tg+dpmFE8Jz/p2bPFdky2saOB/+s5z/mUNz20jFBjQDiKMJqFTzx+MI9PVwFWiAR
JTlrzo9h5yZ1xJT9euxq0VD5gM3VNnWk8CTt5tolzUfnxOFZ6Xch68dtK5S+sTKr
P7JvZaHv3plCYAw59+6T37ByKS9qJUhHn0OUvizR/BSlMkfQb5EJg7LC3WL5WLfX
FXotcMx0bNeZCI35CotPBq8a7CDsQ6xKK7NzUDeKKfalYrw/XFuOX5/YzOJSF5GS
T31n+8de0W7R2NmBV19hL2ye90Ez+ZvSsNZzTLYeJfIQlmWDfkStePUKEzyi5Lvt
PZdBVmzphHy0/0VaBsIRuOIOWdGmvVtAYIH+i7q8uRwr2G5DdyFCxUgk6ZjskHyF
EFesMsVEei38XXj7v8NV9TTEUrEpqfHwk64drlOBJ0I0GLcDaZpk2QA2zWDI4lyQ
FgEJRNMMGkdLKUnPAxmCOiBLjSlMSvxSEsodP2bHhn5Og/e+GxjM8+3r3gqsBoCi
3xCnKm2+kg/FUHyjCb5MQtAu7LHI8CIdiVssH7V1+iXjcvnDI2TJmpYMFPce2xq/
Py27EJ4h/L/Blg0xPH1UXZHl4nckbotlyUeZVZnbZAzTaSq9peWMjKVmUYFyMotU
T9yZYSuEyEL9eFGn3ui+u+gwxkvcU5DpQwHT1rf1iVFSqOlUu4nU5X35VyaQg0g/
GkHVWTVD6SeoteEOnXIfkHYrBn1lJwArcLf+9iV1C0kJMzteHPRjAfa5bssGUGPQ
tceMKkm8EfEkMverNMlrcoqp9bmMyitjWjhDi3n3kk7ndFM1/PmuAu9Rxr8f/zcI
Q7fShPpfiVXhLn+7kZ93EAOB5+T2ryi9dUtrPUEt9OcflBUzptXyQ5YJafbNafAD
4etLkt7CHx6WXpqSlsjaYp4knsjK1mC5mclDm93p/R0iaCQFxTTtnzbaYo2ZmqfX
sLvWN26W2dvmMUuUSqMzY7vuhaxW9poKDxBJ5XGNkY4qtybyY+2AlGy9TFqbKusa
Gh7P+5MsDqCSGumsHJfDg0nONB4PPH0nHE8NsPuINDTnngOkziOc2Nsk0DgeuKQA
LdaWvZvQFv3PjjZVOKV6HI/YnRtok2H1afY+4qXtSWDa3WXUKwANwyIRphlP7xm7
6vyN5Rzp6jY3I1s8idAyVxS/1X0nuRMF5vD5SQCYyFsS3EHNoUl43EOsjGaVwyIi
RIw9uIQXH2DIn3jlW+RuOTpAzlgim2EffeYaM14Yloa/uLiquZTEBBPekbcV5G6S
XAhs5XQA40zTWwmo84WrS51U5vKzo4YheGC52cVxGMB6UKZfbLoMbeNDs1EDOV9g
9lOyiGtchYDxm514HjPgh3hOQCD6I7Zkv1vCfZoRawmki6Suhap5IcTY9UNWnLjV
9sDM7v0rEJ8N/5QS0vSU72Zz+2/AAb/PjEj7zG+Cgya+5PNHVqepSxikwo2nKUKB
TTPfsli56HbTcauGhKSYscpTq6BOuSZncAyGBFy7oUv15iU8Sm/bj9I56oAMvcrI
hVtgYvYEucsXM/j0J71qVCGx27BAomW64adcPrxoZm9XXEv1Z2nIWB2VvQwTldv6
j2Bv7ww1WJrUOSwwzGnYJ229eTGg2SsN9GhkEmo58+zW7WDi5PCvrCs7sKqwo9TC
c05zzBej26hxocPY8UnutYD9sN3hBOqbMWGeHWIw6nOMeSJ3vbo+37HyKDa+DTqm
gurm6H9TNXtZYi+s36Tedqfua1Ue6ljyxDexcVJnooa2R1TG7/fYZtV7cwwOlBPH
9lRiSfndl8eWlfhIfBhlvGwNFDHu3NpEI3FL0I9+xTkmoHkb9gAWAnfFj1sgbXA5
/4zN2Io6usF7+QvCszfCnYIqvs9mwEaOfcs+IVZ4HkD9tvzjbB/gwnvzcDUL+bcX
iF+VxI/TDjBF8fEY1/owRiYCyJwKnMqon3MfHxoETFAg+9styQ9KWobCJ8wA0Bag
5nVgtTwb5vSD49nPK5yZzY6g80UEW3HWThlqK50NjiSEVo56fS7hh/lZDLIy50RO
tvaLzHme0HkPffQthJepgL69hbmHVI4JZ0jHwV1VZ+hyXqE1SzUZpgY5JCJ+ahjt
cG+9o08+SDi7UQ4Y6Pz9Qm9vBhKAjRUxhGwq8Y9bfkKADzOxfQcTRGAeo+tgop7d
WAyKBa2hC3Yr00YwbWsZxxdp5Q+T0EgmlleiAqT6wMZbMkDLILyzH1JASbgNDndX
YlpFPECMWc3uvi2DyQMlC+jm1W7vbZg9rFj2F+vlN9fxYbggFCVHIwbICRF9Fzw+
FCEbru9l7I0ntJMy9ejaGSV7c44Ql5xCyIjEjr0e0AQ99KlGuPIMGjEtKtIb8ZJY
usPaPSQJc/tO6hMCfVQ9xkbiy6++hWOey+uR5I7ZWwbWFugwyeBvGXYqzbHZOiNO
4G+okN/Fz9clS9aOc+Un3+P2kZRapln0RXq1PnC7FIF/YwZI1cYpgKGBnyXp6VDZ
OqC4AER87hMdIe4eIeHn0d5clT9oRVaPo3XzPx4UNHUaWlvlygwtA0GpxNGxcYAe
5CRiFfr/IzbgFRzmkO4l2oPOsZiEfCNuNG4NSRzp7lNhRFH/PMTEenrQwSoJHOaN
IFA7pwjae+zwK79K71sMllZ4pK/P2p44hxGD6cEY35BMtrFGgDEHdK77Y04qVFEx
6f+5zCkmpDh/GyK7umndYh4ozbW4p09SpT1Ho6OeAGdGht/wdgUTaWn9G/bw6msS
XwYQI9PrRtSjiiXkIXykG6CbAA81EPX7+XR/1GU3N/j9YZ4cH22J90HcBK1/kxqK
ft1g7V0Akum91/XDUMIa1WlfcGezx7d+0wMYvaek190wVmt9SQGc4rTG0YNlv0Xq
oiNhrC0/J7Wj7YzqLKxnxOBBaUm9uwJvqbTjUq88ZAP4VNaZE74mwMcPiXy6T0qs
tydaSI/KYvSQGonid7GMgdwj5xpxuyHvmbYzsgsclfXangavU+ifTBY+ria7Pc0A
TBWgANAs5z1Yz+Y1CePbzSSezxLcoIhYh9Wo0++GBPBOHC9/oWeXqMjqOqWioIpK
Wp0c6HxL923uxlxF9bKzh9ur0/Ay7ikyYwqBi2Rz7q6aX2b4lI4r52JpeZy7j56H
+wxSd9Mqgf+wIR0AEusnvlJxNt60udw3ijTErc+l6nWWyzzJLcxlMN9bYpcGooaD
57uvEgU5siTY0BTtal41zJKDgFbay/ko2YTCwr2eOxihMaIS/DDZ61Lpyt2uaL3u
WiigWW/YHUU/JzNVw2O58QTuDnbHf5XaMumIe+n7pF7CV3W4gYV3gFFbW2uk0sEC
tnsLeaqozR+by4g1IgUxuRPoMB8QTkenDuXLV9xbhhV3K2O56ak/KO10eKcqpMtm
rTf5H4aTwLaXy0nTHuxEwTmzQenU97n1Fqr0tuKyTVEHnkWKK2/GNBEUJYFIds/F
MhKCakjiOnC9sSgd84p3VhUEehx2EOxzpN3fWhZrfPadzeexXXbsE7Pzd/oleX4H
pwYDpEe3TOdBNWbmCdaBsozjiftYhAl8rleifISypPUMVFeiRRL0X/PJrSkKMXYu
ZcoQRmW09EoolDmJQz3CfgQcowzfxjIWaGEdsGP0RZgZ8wYamUjhtMa4yukYv9po
Ici/i5DKi+TP1VvgNwMb8J0Oted1uuUXfa2C4M7LUjcDoSJtH8X7Uz08TbJ8si+S
UgDej8LVQAWN/+Xn0TT0ut8dusaATgXE1Y3ny22azxk8NwU33UgXkwqDdpF2lIl2
ytEEer3PlHfO848SBIE8qpcFOwfNzPa1DMZLm+5V8Knn3QqxGog720HwgH4OeN/L
R/03sTj7rzbkweF10mPhiwI2p3TlKqoC1/KUgtEo74xvgh8SbUrojUP7PuQvlAgB
KqNvUBxBdUWc7+I70ll5eQ6ma9at5bPtQnwbXjpSkcYOlgpvZ0aQhfnNtVLQJCMK
brJ33xXzDUX07ZXz4ejHWKJ5tDxF2nhpH5FvKsxMd40hvDF+jH7cBht586klOlFH
4ODRPSuz3k9FXSm/ChXQMF8C9JdX/Adm5XYE2OjTT8vqblF4hHZYhvY9kFUC6qGE
apylMaXQMzb0nakbnQZ+sapGyaadEaDHlXzi4WgikzwfnQpfCV8RJxmWzrP6QNeV
vjjOigYIYCJ2RFCapLN3bQ+tXVP4gru9aBHMehUDQ0nQ5ip8TLO0BYmeD7cI4lyD
YskD9KqjaEPMZjhPx7gM01zYOdHrwmfzbJ2cn69/4ez7z0xjgwSH3JFGt6FupKJ8
sot/fVSzefjoCNyM7kpHbizy69bICxVaJNY3EqQ3G5mAddi4K+rPyhpj20Pg+Pe1
TQUdC8AUGh6OV20/tup9v1C8E+p5YTh6NfFR4LOeahsxRR0rSyaOTKmii+p20az8
C3mRiNKuK34UkjXCLOjACoEKlxMQEKOsf+nnQ1Fgc30eHxlYfBORy7IDuocoqpbb
ypU+fL7VzVvw88erlFtoOtDYz+/kFbGlm/Ux94I45CXjPndAy8v45GLR5TSkF3xe
Zd0luDgfrKYLT964G0zrc5ZI1srkJYdOLmlfJO1JydDWGKjALF3i7ydQbuq/QeFu
IvQXnjZsTzHJ+3/NMeZE4LNfuWSIswTiw0IOlQx/qS1upzPcWuqYKGurJa2zvgwD
kpkuOkOGbbNOZ7tETSXjHNx5oW+qILLpgWlh6rw+c4MTcdwL9JlTYMwTM8/rjBlr
wQ69PzOx+DBRtZ0oZ0A0mWNaqzPMsDqNRCvYokYmsCaFuXPqyislsnLEkTIOrlTj
pegFjBl47DkM1t1D+jQuhtNps5vFhRlyPWKSBhR0RYaIAKt+yKovIxtQobRO3I1u
c5POEpEjsdTB9ZMNWaGk7EMoUNxJIuQGqSFnIr4nlgg+NJMMWPlBPCYgrcSUEE1Y
uuhBXRyG/R/08lKaF8sbM7w4ZkADz0yAFgjqqmwlRaoeNK2KsfHs2yH5QYhxCmAy
7q4bYZXyTCrsQTX4P67u0rHQogMp2wWIzHjdbDIp5J9kwYZHbfMNb9YEDSq+BhZl
C8BFrc/2iu/UBEDNJd6X59vhmkIu8zkv7JgA2OcOk1QmSD8+NZktR7LMF1zfkaYU
YBoDgVWCH4+n96cRi3FcpXNEBt12QkmcwJNmFROplZ+QttY8bJzBgRJ2OIshC4jc
l42iOfR7Z1Xmtn7T8r7jGfclRhRHNPxiPvy8ZfOPcTqhwQiYtMSzffCJUWucE0XM
FBTwcvq0z3YHyq4Udf8NjZbKLVc6MsO3SvfPscf7FPVZu9ZM1j0/tSYqFiYP6yjh
d/MuLf7/+cnY/DeHcc48uLpIYQVw9COrkiF1r5Tmqu2/uqlq2ZdWxiuIY3uGChAi
Sfz8mNua8JraeY6uTyswccu4k2r5JSjgiL0Sf8RcFhoD5QfsfEy+twRCxRo6MLNk
i7eb9LnhO1Q5DM+ogtHMVmX0l/71UOq3QDqzguQXokH/4YrNHN9FTnnWf+0befNo
4NUPtYV9Y9aF40YR7VvrvzGZ50A9koa77xWPxARfs7yqIKsNIrosljMO9QCp6f3G
Pd6//MLtvvHKdtvCm5X+5ZNEu/VY66RSaS8mPkg00q6jS0QJWGYYsSBedtnBmGLd
6tAGLDCZp4fFH7QUOOYLB5mK/QLcp0TBWFoSLupb+U9jJ8YT1nOn+XAzN26J1xKr
qS+xZ54EiWez2ARkWAHlj68Oi7uY0+VlQ6YQnRy9K0uYQ1lyk2lXfLjhXXfZ4GkR
FXmD+w0Gdt9Tda4WPEu3Tem1uCY8HXECUKNJODiuWZ3wXNUKf3OHz5xEg+lxe11i
6qSQIbCuGM+j8nx41Opw2wNM7i+edPynz3qNZ1wNf6RjamPe56AMtMwxhTfOhbqJ
8N7E29cVpvGO/s8Ilm7F0pFLQ7kGlGbTkdntFEhNoYPaxrG4sdKBdpL311bX8PpN
P6u6WCw6q0QdTPwUwLR7jGI3eE1o/IR98uc1tlS33dpfxgKR5SagRLmeoOola0tE
ooRpbVR/bFB/tSkUcVZ396I0GsBI0K2/vAwhuONKGE9Bfrr3Gebl33782hQJqacU
HSkn6gfelHEcbCrSU84VxmqURN9ueyGkUVs3AyOllMf+BWIxEmWXeOEoh/F2pimz
7XEz1rxPRZie+J5c4vBIAw+M2yPNO5o/r62NgTc+9iP+hW3IMywGXermmoKx4fxn
1MgtGcXGqOhoNL+rCSYANt8xdqP8aWeZzJG3dDKHgekIP4vFVXSoBdulCh1jcyFU
rNkHVBmcZaS7HZYGK6GOTFVkry0QcVag7mHAGjdxxx6tzL+8lg6K5Cig2HfMTTL7
7PsJDgkkBqGDAFfWfjsdowHOS6WfGPZTc+Lx5pxqFeYcRk26jO6aJ5pOThAsKPuU
PUC2BWQEEa8At5kdX8VJWtuZkXdidRvmT2K594soQc1giX1PYBYeNwwq+8fV5lpT
HIWmqZWgsIzscm73cfOLEoBczZFGqbomkCRYvCITnSngwFhABK0TKQ2buoawHqQI
G3H4yVLzdSpQJQmxIKAKEgr5tzmGGPRPSr8iQL3wDHjfSO1ZPgRews1wrT9pXt42
PVk7fm9Nuoof9HAfgkw57KWvT+8PBroH44d6vhCcHUaa8AZy2AC7TcdyFAtxNkqX
Ywq4+p8GI7e2hQRwF6YbGXBdXR6oSCUJ8aR5wyqL5A2R89Lft7i8xJqDAsLQPiad
7pFeNifH7DVRBGpQD42ybd+Jkzn0vTXldyXX5BVRhCZdF9WmgQIYPPhx6/z3Zpn/
Olw74m9qt7ovbDk58E8SQSOlgZeFXKyLv8U41E+TPrXohOWV90ViE+osW9qEMPR2
pLxEHIc8e1xiinTD7btruVeTfJBrznK7Jt19jG3PCMySNtEwIMtclwTZmH6MJbDS
9Ros0lqw4ct9/tNgb4b5E0P+PexLMmlABYFAZtooKJpkcGPkQlvJm1xpiyiZ128p
ELZs1x5avAu+ng8fryrPSZSet/IUQJKb2o3lXVJ5e0RWmnLMqvux5UW1xNFIhZup
6yTbtqqXTf2Q0shaxXY0WAcmGNC9wFlpA0QytN66d7bwixTJkte1liiSaofZzlEx
SDskz3U5YxMyk+C6EfdbBGZYMikQjLkVaMGGlspf/EkhTzIziltswcoRBeKPOrUJ
+/Aqm5mGboyrwN1yxgQz3br2hnOlDxXmtuwrCha4OuC3wE9A8DvO0eKRoljSe97v
OZCl/xZTA9Ws69ZyNdzw9EDVSH5XyKed/ji6L4tG3yzV0vc3UI8Ep03R+Qvtu5On
FM1RjEN0RGfsTXPaOvG3h8WN0tmpZFwbTxM5A18JIJdPuh95+Hc9BJDOMWf0wnMO
zGtNDR62V6ZE1YoY6aPwiAM4O8I5rGfxtwGONPMyzpnpSQ05iAjPLwDNwgaB9fk1
JkiMzGoJEoj0TCtZOgoKW0KSK+7DZTIBGvMZ7vdO2YkGl05H66cdf0cd+sPuKWc9
JqM7D+nW3UCSJ5xqPSTZzXkUGii+YCglzTFNGNPLPa3FZBPe87AMLiEnwlR/cmRT
TEA0hBYZAPoT7kBQVALEhpDt0gHdcOR6O2BXmWvqDArxvpmqafglhM8IOynN4KfY
oefpfyspuQ4v+R4ZpdJEne5Vdq16VNG+SNfUltIPzlgpua+nj4IjyDVUPUA4gQWF
DihsYyIQkn2n+V4EasrlCRZTGWmMch2/qL101EYgxgzlXOcD1NLNFOsZ1uaxoHy0
6TfFQ4TrWn1qKLKpAFMx2vfC9IpI28rPsiVIyXJlBONBFUw+rESTkAo1TlKL91L7
rmQAwII5TqXMjNXTQqTzlNcGmQcJHfXaPBzD40L16tpwcvTk8Aa/EqR960KYnYgC
ttbNRiS0WOpvj+gJUdrCQNILC8ahpuHYaV6VVjqzRjjxMaNeTzz0GaFdk9vidlY+
hSXTEn2QUfeTZqUF4rDqT22UuiYnn48IY5ikC0+b/GEcZq2IrFPTVIOhP7xcfIaK
Fo3/O9scbM8attVD7YQXD8IWBrwpIlTCGow/wSFDi4fwJ0KuZV+v/wBbctpl2nkY
xNL/DQ31caqWU8m37uBKlUZj4erIRLcTKsuk811DHEK3HpSwVbXnUQgkuSSM0FSN
S8i4caJCtuDpGpM/b1JRwy/36GsvIIEtEdE+PRyjeOgQqSF0iOuYpoqYQdEUSYIT
QP/pkhW+negSMAJzrQ7HRsAcrOjfo1FP4lZGijI83Tlu3LoOvyqJTveRQmoKmlWi
0aSi3H8MZBcLHCBzOnIMjI+7VDZ9JG3UPEjok0zDS7WFByL67fKIuLZyn7iGa8aF
j0M/ZLOja4b22VVbt1QQE90Si5cSoCDJNWq9Er/SJ8rNUJnoEUA0mWGnUiepTko9
3JVqnG3ck4pCoSOVWDARUXEfrz4bWR97RePraPfCZDpd6bB1uUoLus0yhIuRz9Sd
NEk9uMz+zgaH0AgWF8KEQ4iaa+fSH1jEitSKdSKhMgNakksOInaUv8vNjswvl06c
SpJUQTSl8MxlXkMLVAUKNvjOzo2gPJgJBtJKqT72kssp6JgFaEZnVyd1h5OPO8Pp
VGES3W6fspqK9MkcpJfiVxm3LDGkcPd2LDwj29SgKeQ99CAr2aOLsNPJZDc+vye8
gp6K/jbfhz8ALVZu2wz2K1bhwbvWTmMMJw1DgV041zzwAXLxcpXdZ6k/ENxqM5L3
EEnVpZIHwlsmzRP+1wSX86DlJAhCI05Dl3sEtI9GWeqQxbqusOQIraFZO9hDRoPx
Pw0vzjtj8q5+rh3TizpGGG/Co7J8ERM2//Bi/uMZlYaesNWJSb3iA+FEqR2afCmq
8KjRkvGfexuBySf5ztPvRj/s7kZKOAU60zBpw0Qs+KSNI8yLH3aI1Vg8zUWaCAL+
OLfOq1G+e9ttR1Ys8QSkvXz9ruH5jCRTTMEhtTh0gImMcioQU8oh7/a9lFpRmaZS
6ZF3NdmzJSpEHSK+ths8J8rcDGiPCvaq2vpdcGwpEHZPf4Yzlf8baqGA1Ax5PGQk
G7TVpqYebN4eBTRUNeomWnY4tzy1+lBGqMmpAeEKMJLo+1RihMHvXPM6uTXTrOM1
srlFPY5ZG+nijNOXIqaOn1Ofu7rnFq1aayGiuOrXeJC87p5+IEQJX7dPuIwC5uH2
rxSKahduHBCMRCJHKdUQxBc2uU4iilAFfEb+oFQx7gURLJ66T2rOUSaLNs8ECZLg
v2/XQB0/rqzKHn/eWsQ2MTdXz+o8JuHTM45uyJbtHjqvrY4KYZSI4wS2S2Hz0gou
8wihqaiwvJTynFG8g9T/IKRT6Wcq9pcpa5yXfCOuIEesgGLGj9mAjh2WLD2b/2Ms
TnqwkdiZYRT4QEF44tv9BSyETQ5MxJKdqpwTKeMTgnDqdMXJYnZl8NLPGZa+BgWA
Q9iQ6nyNRAsl5v5asdHxZBzljoGSdSAxahQTXGrDPydbNg3vlaQLhsEg2KoXB3n+
b7PKh2io8E/jY4HLGhe97vzpTsFwxDTwrxkzlAw/B8Yztav2SkVjRQmHoiASjmcK
u6DBlCDzca2vtYiMvoD5r9t4QanfiBu/LvloOU+0IPOaIz9tYHZM3mdpabm2UPrV
jJNbyuZq1WCESGf2AoZi+YEq14Q9+yQj4+xtWUGrF668h85h6880kxoAqsi7P0xR
038E+d5S4PPQWDN92OPlwmmhbxXVjDvvHZsvf7HEe90idclsk58hcnYvubsZ7O3+
Or42dYrw/jORrCmkluoUS0JKRWLtaUXNATe6IyK488d+W+zxQp6K7hqSs4LAQ/Qi
0ARy+ci+1ft3HMKtXWiOjeFgM6phIPaaqgBa25cUlfI/fHDip0lFlkgk7VCwYgkN
C9UDjsn1PE0It4o7D8N71jIQRaWEjeA48X6Acnqk2jvqtv76aWLXDng54sSnvTpk
+WoQjPlhlpG2Pk0a8S5YLzefvCUDJGoVydNJaLDDoqQe+We9mLucldXcNgMzAg+j
5+FO/SGy4fdTlRB8SO8n5Fe/UGjtmlhulqWkfYLRMSAmaifZANjhzxx5+p8DKw5M
5v9via1c/GptFbeZzCLgxHguLqPFa53cCMBkistU+Vi4+G3MED7cRkyQQ9cKvdoG
m6AeuwX4CRO6j/p9G/m4F1/86hynlUYtprkM1W+Hze1UjwBXiXW1/Pg3Ygi2z0D5
NsM1Q/OPwxiKPjtGTiMfYB9GVekL79MnEPC3fEXC4LiMqTFVIMz6BN/lKoZJygjM
1NA1a/HKcciDV3NmUwUt+kBNIOuef7iKWRi8ydNA3QclSkIMvCOtCdPgyBP4TQWE
9nX61rZUBFd5xZVEDChD4aF31C0sV/PvwTZ7adLBrWUWek2H6wqS2jyt8YW/+wdH
jCSgc8k/RpkFkqe3rWDX9YxThG0HwiJno5awRbv63jp/OC6thmOONKIvlh2+2shW
snlbOj56oE3fBQbiKLg8c5MtDbjBs72j0MGwJUvSjnP5aK1bU/6eoMdgbtPImpwN
PNcfg9bAm/9aBgrRolm/HytJVOGxvtLLT4yjVZeatC9TI2TkcftWORPrrhnO1hZN
e29NVYvlUCvX6rbh1rEmlChZa89ESy6uxGWGcnAPA8VRhjNA9QR7gJT2fPHa/ldk
FNIhCBd1rqiNgX8SN6cQi5ML/uizta5sYwSucWTeUV4ddMjl4h8lAtbVvj429i+6
8wbNMZxErMD02ljpmU1DU0j1kUfoApxJyTA7iwsjbnV0qUatPJP4TOHR46TkBAj+
lYjTWmS6Y5Z1C3aRrUKdJC93L03D/KHCEYSA6qGIaMKRdeQTiWKcF3zjrAegtp/Z
ZmrKRIZWu3zFYPN0TB+2AeaMluR8o2RIBqKyuyYDaIFcfbffuqQ74w2NIR95W1xd
SqYsRYx9NjHeSMaSSkusK3i5zdBUP6811sV6ZlKgXXTPTBIBJiWrSHHRXlBWQHvS
A4cmV7iIKCbdvPkFHzC+mqEaO743UbOYOeeT6B9SJ7An8rCG/fGx92hvyHCk6yRB
jcfTPmnP/u/idkNksdb33p1pdCW3zty63K2mUVke9Pdclln13yPZLNji2mB+EMOZ
6bomB49GKL14PTGqndmj5Uq474DokRry0mKCll/RcT5VM/VnfePEdmKL0ETAbYK0
LPXYvP+OEYRRJlM1zonmxvuLOk7LRVj81RxRQXmjeXS9BA1LY2wGuMVGRnOh3g0H
TofHIcEPJKs4XOGb4r/i/KTQjWcsDGG1NbAW9a9tfYNVNKFRjy/tbpQhY5I1m8CG
13xW3m3YOL7sRI4SjjKmFj1UtsvrJ6w2Oz11PE592fh5oCqenb2nn3K7S9zNm3Yo
bpdPITx3XrgXovcQ+646s+Kd+BCgfLwVD3WtUmtaDmujbpkGQU2qiY8dbnjdWO8K
TO2E1UCJ1UmJw1CWhdMkNuEL3MN5GJchs5gZSa1acv6RBRM8tKjf8a29A+R64tn+
r0LFQXaX4Q8uCdA4HnNh0IrEPhBuOtP+W3pcTc0BYFFCS7HmeWaIz14lN3EyJC9S
CT3xm3X+R80GTcpg8H9PhQkGrLOr8nnqOT7yZjyAiMgxEHvhPVjiF2Uvop2kYwWv
tqh/ENvGt0zYB/AEWCkm9J+J71IFSwFadp3b5jQWtpC+KUiVIBvyKK6cFr9geUZr
75m9NnBPDG6eS9h1lWx2b79PBkiNmv8w5ikmEWRVjQP2G8fy0UnN4EsNl/ozGEPI
`pragma protect end_protected
