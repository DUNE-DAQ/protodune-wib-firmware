// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V4RAH5qkA70G1NREUvd4tbgm4SHQgOMgjG1tQsasrvSxQ47NuX3hhm+hds+C0qGd
rU19v5MrQXcqY3Wgccdtg4uIRjdnvKOM7m3s7gJB9pJGTkldwAJ5OrbtA9DAoBua
OAfBPSwo2ZS9NYZ78kevdlR73VqtdjQrzUJV7ohYMN8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32976)
liPjoMBLG/OoWLn5m7eZWIdYubI6eoYJXceNJU0tm4zxJ2PYP/J3dTSXJlbw/LkK
91drw4h94ci86GRO+0THybfHYaulT0jOrAbWDKr/nj/jnB+NHW4f/Gfbey+2ijTy
UMqU2Hg/xDX5/PZeemJpb5tEccDr2JT+RO+weE8w19S4mSRSLjd0MYAPk+hAKJF/
EeTfTtjfm943ZzXQ02FHo9MtPmljqhgA7e3CUAfLxqSQq9CNQVN9OjpeHgSwvu8U
eFIB+rTM9ivbBNLw2Ud1GfUYi+yfoBXtrrIYW/uwD5OhFCAXQYpNNdijXt90adb6
RadjJzezHs2n15Kyk3YUDlPx5f3OPVkgzGpFprPU7Y7mxehmXXAzjQk+ZvJApJ84
4S3r8d6862g3xCjTxIcWmbF1qQt9rgD8e9b4/iGmc+NfwG1gHj39sFr+VkmhG7U8
QSFAJn5k08zzaO6CUryvOK/A8XrjfkslY6V+3iaLoZSgPMKuOOG+7rCFmLt8bq/Q
f38x0FBd/YEeRffOEc0wRNI6zsGrdqMvH/mEnp7QlzCx8yXC9E8hxPYVSWeAHPEq
u87cdBn2FihDqwPr6YrJW9HjNmo8i5RDtgugmij4zavfc6qEzIrQaqMd4UYN2IKw
WWUZSBgi0MGLgTQWXi7bXmPiG0hdTtABQjHxF1GuTT9+ajEzQdISxieRpagiX3Ob
XeSzzShikf6DQlJExf9O90wDFASq6BSkccFfODkLy6sRV4zvNf0pFzG05N9ypaSg
ZbpT3LasVW7BAIFl9OT95AENBTnBHZPp70F4w12Am6KHJnZPlmIL1oYFs051m1gO
X/yWKIx5pwQvQJT17vzonkKTKHJVBHo4VAOkScm0Ul8L/H/R8mgTnZBn2eNb9N7b
NU0Fe+AwGBDmAyHOL/s1KXI1QCTuMioc3z8TnbWW6P7gJmUH6/6JaSDL2u4wWLP4
HCPElG7faZniEPYntBatgfAZ2ZKI9eIlxkkwTDS7zGWDgPcyDo0vEj0PsmE4gXSK
YFe/RmqaaJp2HKLly52xwQydj5uM73VgXr7eNE69zn+uBQXzL+96DLfz1vWMHgVW
+Wdo+KLHUXcgVGI9isPLLZn/Z0My6MOuebLFN39mu5fvcPAys90iarB/NKgRpY+a
+La2FxHenW718m0QdqrdFSe6bm+qTm8y9dZFk7XfoRVzP3BYLRjYeFmyuRDWuN2P
l1P4SJwhIHPFV6n0scZhzMI/48PXcsztgf6xKZQOW7gppfv3qQeg7ZJvqxIR0X96
oYNqUkEJ46IThPRyhux1577HhbkUBg1IpRGesh8KulhaSmaIz/lmGLJOAgps7+8p
8CzpA3mKJXQWXf+d9so8phDKVtluRtHezfspokwhLpscm68uR/MeoM8SgXpjquhz
CBUwOhC3ou8JOnKh1zmvyM8MqavTl5zNBIC/cvcwxfjtmRR//Y/Hn12PyW/soZS/
L5EqXLCkhmMsBWRtHHTF0OD7YH0c+OqZzhPW3rr46si3wsXC7bJW2yGEQW9ahKPh
Rv0CEx75c5hiLTupVMtxITy2NohDlTC4Cnq7hNQ4wFzdyFzJhaDPsCjlaUBSYFLI
azkcO7FXqnTiLz+iXwD/N7i/JXzckS2j+iEDc6jjt3GQCRYpzVktvti5aPuZFeD0
LbDNPKOy4ju9r57L+6p68TfsBQy8WvNWFgHX3UxGxwkPjjNx5hkK9iEYqcCaG0MQ
yfymqidSrMKAZpASfZS3WMBUtLNHN7Q3Jwh6HEw47pqPBNkb0yMqIE9R+rKXat3L
znB18fXBavW6ifAsBn548ryIIJevOX+Qv9sJbQ4jtinz2sAJIdKoINPzWPFBz7oU
AbVHZLra12uHh9KVrGwncMctyo5WeHI1eMgGxHK6xjxs14kySjPTjQC7QdMM/vLE
5ppup2kUmhKTPGKGnfqoegn/gLlu8a8AaA+fFKgN3kNEHquLAu1wzoPSvpYxYHG3
2uoAsvTPF/i9+/IzSVV/0n2vGcVKWeFXlmbNSZi3i36ZvyfyrM7umn4EdDj0e/cS
8AJa7cMiEjiNsBq4bpqkCbqmIDUIzttT5i51SjkdeGQ9nFLPHjNnEsJZ3DttrLP7
6Roh903fnhYVj6MkG48mh0Ik4603YbySIy40amQaUdpax6UMjkMLzCxBNKO/gaHR
sJNpEnUF3l7WaLhfS3cO/FYOEvXYh66+DPSs9tChlaYxgGTriHB5idOlvrDPCiSh
b/2owhoGngCdLkRr3eLbI5mGtE4dt6JVj9Gk5lTpiJhEFyyDu4p9pGkMDcr+zywD
UPnFemWf0e+4Yz9gcrO20qrLfd5/pIgO2oKgFURJZ0TH9yV1uufLCWwTtuvRu/ek
iuMx99lQdhlTaASghr5BrPC020/lkIfpSaZjHno26f7mApfUIHs5/u0syrvvwM8r
mFFtRj63dha29fgl8ak39kH0IbTSL9nhII+wBXTQDPxMccdO+UP3vPjpq22Z30KE
QJAnRmo2p/c1Jk0TkCQsx5wYxSBnY0nBjIsEOeAbWSHmZ2ywdjhtIVklzBGbN2DE
SaDVLph7Ht88C+fTq4a2qAV5QELCVPF769GQ77WciyCJFrViRHzp6apCkZso4xAF
rkrkBXvv34kFOn5GUsf3bFMe9nbn6NGmPhetZBtmVy8QWegEyQvWptKzcZl5obU0
GACDVV0gHpcEBonD9FMAdpb0qIatTdDTER1kg//XaZ09LIlwaYZkF7vQG9vhyLfM
OPhbEoxcy8fWIejO+l2fQkkb/EBwGBLweA41ctZXXR/u1nl5B+fg/nKTEdWEl3rO
p7AX8enBzURHz0ryzWyP/odtZ0/z8jM3kpArcBs1ektELe6Y76LKa9IxvzpTBPfX
0Qgx5JK0aj4TfJzTEKQDHK3ldXZANtg7F/4tLv8USrtA0Fl5sZRFgrrrczcEckvm
lxs9QvlSCroPwV2kmc80KrrXW7jW7PISVDFzSkXtCQvSceAK9GmGixcYepuUZKQb
p3vPSI76UgSK2YnQQh5Gwhxe81A3JgixStQn/gNYMba3XuNs4UzXjSXOPiPgvzk2
yB0eHU/bSdXFhj+SpgGfbctekyinEcTPDkZCQW6iV1OO9s7KKgaOX8DUFXySNgNR
HTJKi7ZJL5YdyVD2ZrbnkrEp9AccWKr1zOHDOXw/xp2JlAd0zyyWUn4jEClb3XBu
DIvloW8c+xaIhuIVhmAkDcaNEZTcIu5nW70UF5QDX2S5K2Ed87NL/emKZmnRu6MV
fbbaQ6b26HlvYj2zGajfa0uquXLE+zIKcBl2+0P61k7IS75q7t/Iq+Weik0rjTvM
PBBfrYyIVj5Dq1zd7ueNyJKxraz107602+dC5Aj4lRyoiHY+4XbXul2NeZJwWVg4
PrT9115fkJ+gHKOk4g1Fnp4J4aBd1ECSR3slmXZg4vjdahT4O/+tm0Uzt9K6fpG5
kXV7OiHvzE9GA+diM1WDOFQ/3YROfzF2G1J5DPefGoNlz5WohPdxMJ+D3Mu+JyY/
7hP0KZCn0hcztnhnJir8NQysodz3en9X3/F/u51U8mf6zGkrnWe993Vry10D1ei9
dispdHAuDUkIA4Jgz82z2ZZeag/ojeKWEle2QKg/5ZWnwHuy5VjKHjAIxZ90/zr4
HHG5ek9DMvpgWEXIm2TPYReQqeehcTv90LVU8qpi6syx5QpZzd+XCs48+54D5Yv7
FxpuDc0Hom7qzmKuDmxFEYxv5Hg0VdivYo5/5vxIqLBuXuyDFIgiDVPGWO23WyW7
9QJkQotpE7xgEA4WnGuLkt30mI+hdBPd0VocGACi2lNhT+HAFQHq3CbQhmVnUgCK
U+QHc0lnQbSRP6NGuQmWrbgwld4Nc7DASuRJYIcMeZWDtSI+irR9Tk4E1mtGyzC5
tILzXzgdgy+i5aO4DGCSW9uHuYPHCOLvyQ1NIljpshr4/4WQTeZdASltUJ4iK1uC
8OrmdjOja9FVzpDplAGHg5hdVOiEBt57V+AQCDxVyKgYDyJwQR1pdnjXJVZZ32hs
Pc4UxH2BjhHJIPtVztYYbyZeZBhRz7LnutPuKeYfdjCgNJT0UMQb3xvKimiEBT2W
krx1vPrznybdUq5sIZ0prvivRMpNVJogu7prH7IUFDFYNmleP5gH5nGeIIERDrKe
3dg9AF9qWSMotwGKy7FpY6KADG1Xiq9V8Spfah0P/++zFKrQ9oOeA+qtgjJYnd2P
sS7RpPDFhCQhxjfy21cRvowIwGlpnHHnbgFi+b6yPgOhYimV/ndiFILT2LnSOj+k
BBDUo1XYclCFvEdAxv2AJ6Jg5qAVOhriHSgX6xbe/zLALi4YG3vW8kntcQ0Q8i9K
ZmtmrgnFj0v2+W1/3t0LTTi0mg15H6V1eRSOvKIJCLgKdFcwMf5hODGIWRVvUCjT
m/N3USSBP1l+bdJpP1KbZoxpxPhVCZQExkYT5tnkrglwsZz9vwgRBbGC5MzGGp6H
fV4ORKXmkKoDQ7E7Rg2Qkse4VoYRV3OhS9CqWV8k3x189QBTZ/xz3Ce83pgKhtxo
q08LuhFJkXWNJAPjYvx+VDomYZWOxRQCXHU8EkM+pfjIdEp5Tw7NtBBpc7fbL42U
PvNO3G2DFYfbufmrKhBBpgzsiD53BfqKA1fUHYaOPZL1Agy3bDpq1b95IsBE4L2W
aV5Xbv/eWhLL+mZGW9jGCpUiwLcV7atyLaiW0slo4H+jRo5bcTG+AW7O592XayEe
9rDrI8iw3ZLhbxn3ay6n9Ul3/+SxkjpjsFKLSbmMCvmpTijCkKjEm4AqXDurClPI
H+aMVB5Y5l6WiHTWmlhTRQeExrHwUNpU3dpERszjF1BaBLFx+9nqry7/gDL7aicV
kUmOcxmDEi3FfgQDvCek7027Rnl2cUwL8MRhry72qZRJmj7rGyeYRzdU5tYGBNCE
dt7Kk57ALEadKgbOeYw0yNCdao6fUf45j931Ux29CdVeilk1slxav2u/Z9Ur2LdH
xTcYNQ51CyRJFwSKeajqz8OfRiWW18DQqXex5jP5q0+nq3Cut3caiHDAwTQ7m7jx
C79NXJ2cYYjjeqi7YnLWBlZaWu7d7oCL++3KvQJdnYPw0upiqtrwSDg+I0iWWwTn
BXjuyi0mQcDtFCIAbatU7PeYUh8sXF54KK1M9ux8w9o3kK6Y0GwmsOMgAtBsQAdE
SQonEB921/8AmCjJQ8rfUz3QZbnO9qj4wigIbUBgH969o1DzDDBLMLQ0Ikxo52+T
/myPNWwpa7JsKHmzsN2VsaaSjlf0v9X7nJwqpiaU5BgQ9ogeiF2sCFN0nHOMlSDZ
DtDVoMP7Adm5exzc/bevwLS7U0dl3KtCjRf+Kjn04OMgKXuSn4geXAI+S/HgdvuF
mhPrL+liyCqYQ33cQg0/AJM2GrSJ/K4s94suUv2CD24oKksCo5zPliVXmRbkUFKc
7PxSlK7rW/LEE4ylr7PBIzw32lhd5Fy1+k7DV8UoFvikaEuDF9/jVEeyMGl5ApHy
Y4evzVjg/OE7ecslzrwvcXETqYzztZyQtBA1EF5IpPWVc0kLXjnTt8ZUcEa6w5Tu
BmM1+qB3/s5+TaDWQfu6STu6MJuevC9Ul9tF/6+d0dToToSPEETQ+cvdzdZjc0ly
AF19vSEPyAJt5rVDcXvde/w6MbY2i0M4reD7KD02xg4alwFNkzshLe0t1y2G/1CH
M0tD39SzcUpbBRzTYbhS7DOPprIujkMCrJbHRcWUVxlEMCqjJd3bC31R9AJnxC/a
fncOoftB9wADq71BU1EIRXEZzUFW7ThW1FBJN8oLswaI3OxAZtfbmQpZV670MBTh
6a9gENXDHKUbtmfKxwrOHNvaNtznst+Q+m1laPPxKG3bMb5ebZz6hjb4OfmoZt3w
qRUqJE4lvIcURI9d7B6Zzs9fWXKmRase+QHLSUQwTsPWIEzs6DwNQIJURbPqhHRT
K1vbFlzE3C+ZInClvXwOeX1lfxr0pwq3Og16RQBW7+ITMMh5DE+RZwIm1nLlXbQN
sJyqGvkKjFo32RJMiQjxwh8A0kTCLgk72x53/mm6kofBIEaVxDJkMUAz6QaI34nG
0vPBrQdFKr3czfYy/flZcrxWhT6Urng6hJ1y5mUeH38RLPTeqow9N/f6XYKPBxh9
QwZ1AebS2ruMMWR3PSYmOlP9aTWmrjxSZYDgUcX+GkTyZIBkY54NH0/eFiuHnsm6
XO97HMYZZKBtAhs3fqUDKddyvObPB3XlxRGWANFcXOWaUkk76MycMBVr1NDlmFTC
nFqzTwuyF6sKexl2v/pg5KQVzBMqAOoQIgvz8HH8+HEofEJtoZrzmiurZo97wd16
Ev7egK7ytGIL4Qcr63cBzY33hKyl124tx99ZVyzqaxoeJmppHnw0lQC8w9J1kCER
MC1YOA9C+0LZAtLXi0aGimIBib2gM8fHtMbTbDORQPcx0T8wxcuZQfVx8OjpqWWW
XNVxiNUYMzqeZDpAFmERgEqL0njyT6R0g4ohTtSKLYuxL5UDdn1JohsrHei4X3Ih
dpF4m/jF9UQ+JZjJVSrE749L+7GcMSvbSNO6fVHCYKdRi6BFF3EDOHMkLLlViT0d
Ur3wEPk9cw0KnsuDKtS/8t6RYDywRn2iUSVINPYzRuVXIRWD2DGNkLkgiusNGN6H
PsIhEGHKZXuX/W4GPRVvfrTkUdtbL3krtQmskQxxhhEo46jrhxz0zIaJd2bVlL0a
sJzEAsTXtIqcEKu38FOUulRUxgaUIt0FU9qr3AW0y/aTOnPVrjjKxOoDUu5yZwBT
5kKcU8aAPN4bytlzkG1uN7CJxoU5HwcAdvRwU3Cof+rkW88Cus2tEMzoEJLPHc7W
KFX2tkOSs8uKe3CJ1KzMFl7XENdlpJc4qPPpjSbbsVpaDtDBlZ2aRjb16B/yYjiS
Wr4UcSTySugsLqvVLGj1sTLE0L3+34R+fWyT7t2SrUc+ssCNjcnZNzZNfhOzu/qm
+19onUMB20dQW3Q/bOS+XPgRvz4/0VJT8e5XnTCvBKn0OTstzXlgawH+f+U4yQhk
EIUFBzZZwEwKibVFDkmGNPzhdexHrxyMlT9S2FKoCItebGVe5n7hPeg4Wcn8cL31
IUpxeC1Ap8SA3N21Mh6jBUBtWDmVMr25fR773TotXFF1oSvLTUfi7zTbCvexnPom
1mvVjyUrYgtWtEcnJSBDKWeK4htE7eJ3PBEcw9/c0HoQe7Oc4hHvTUu8N/GVlway
gqjhghFxUNcHT4yGQRUadVPvKfCbr+SyONz8AieuQPFHUyt4g6jkB17FYHLnwXMh
Je6HFuVjoEabAeSmDEMofcTtKldsIX8+0sMo1+Ax+FugOXJczrq53mW09fxrMB32
VWA/4zJP3UFcxusaE8XyazcELEeJEMxJZ9cEz9YQrD3ATB9bPWIaESEsYeu4c/ja
2sUx8yRD5jaaG8/WGThW3tKfld2VPLOALGYUb2HwxDGfHXjV9ZerfsF00NEkZH8R
ksTUjnE9yfIAVTND299TM4sPj8Thpne0PlqJdKfE+lbATf+GJeSVro0xUQPv4yCp
VOChSu3FgTi+/fU19xGxu+HXZuyZmkqC//NXfd7Qj+wRUWFMaVXxlfb7YNwPGijH
SIo6GOOerusMIONelhCoCXyWItF+SgwNnKcMX2MQKK4Gih1PWEHiPrM825OjA5TX
qdiMGU2SYh+a9AMF/1sjDPppThKlFcseHrD54FgignGWQwDLl94bF3n6nwOMrU3Y
5TfvVdAAG3jVyFgEDYmPjoWWifFI5dEWidlVLUzXwqLV53QsRbF0WoqOGr5nt8Gx
jbqYBY5xSrQ+m7ONoYjlAZpU/2ukY7u8M6n30tPEUPpfsmcbDQ9IbyhE1mivigrZ
towpdi7niTtPYIXWDUDddZBWZcSP6kGU+476frvW7sGbKQ7//l2e5a9rsMdGEXXQ
qwU3osiwMUgBFNphXcdsiJx/Wj8RNNVECyj38iXtzXDLTYqe6Wj/WbZNdFj18FVX
3SHdV6RFPDfe11yWh/6HXiz6gWB4B36h/PwKl7+UJrGe4dDAiimAFjvlyfP2qIKr
2P5L2nwhTxZOkVtCB3T4BVDU58Jp5+4y6nSverWvhD8EgNlcZ2DK7WM/nrKX9ek+
heOsyH/QQ1vrh+81zgvsqo8+buAM7bEOA4dPJQFpQ0+W2iWBhtZmtfO/6kjFVrrF
OBQtKUECaO8IMgTAAyCsQ1ld8bEedJYlJMrNHGrki8/yjzjcqRC5a/kTMjkH+aOq
YfLvZEAbFYZILXe+tdK4xXQ/dFKNfh8XhnyXzVlZEyhQ7pHF22fIOGq+T9Nt7xUA
DQAFcWFBw0x2WKcIyeqieU+m1NB8f2NzFz5GSAZuvO6vH4pUep4xeQKnwkusfJ8o
stEvNvWdpkzo3jV3azHq9i2meXcTeYuzJVbjqR/96plId/wg1a+k4kOW3StGRjcj
D275e4zfDx/BrA1OUbHdPocueJzu/eTzTnlFKbdO06jr0uwiCxwibpB+83d4lh47
EHgBtpWcFwXaaUR0QjFgInN/9aHY6mwXzyCwMjBfT+DFZtVDb91nwrUr6aTinyDp
RbTeNSNYAvViSLFf6gPBWrpzmmutIp0wEJQ7GnLfKvgY0A0FzS92YuMEY43eB1FI
sMhfjwiMdiz+TR8Yn/Y+NNFx2QN9wUVu0fgWJAkV1CBL6IxUL94OoGd6OCr3lh12
TM00ITWY06qbivz3ojZF4YasPiyuTSQB1Jp34d7n8upM6LAGXUYAMmPvyXzO1JBh
jOVIbZJgt3Mup4cIEyHbjdQied0YHNOU+PYb+gd4H6yjGr9wiKafAF/kKVDSn9Vk
6O+iPo2zcwMGLEA1TA9CqCxh3BEWpLg4W/d5cFQmy3B9Lm/inNUEdRR5Oif4LuWI
urx4ffJ8+uahL/e7niUgfjnxZOXlawbtIv1i1hTo+aTBdqEBro55oQ82TVPF8YQ1
Lef9STN9ny0T0IqzkQZzpLHuLXIgJ7ehpOp5nE5pnOS3fPjXBCCtb9kuLxXfww7P
a8yOVvZOg7HIRP7cyySdMzmG/dteVK/F3G+WcTGx4c3X39Duqo0cNzjzVPrjZNel
A2T0Sj2w1lKp42kjndxpRj9VJzDYM2gztucF0wqeKoF1ftxPCQ040kA6jydfzcJy
bLClOmr7zXqwRkIByQwijRdzC44+u4WS4i2uXqEN00dM5iWLjSB0W/O8eu5E+R6w
x0NLfsxqsH4mrOF+b4md+hzEj90V/WAdymOXQPZXRfOuC6iudXmclDNwVnPTCkpu
rfFAD2LSwWDFUnC0XPZUEnAB10iOG0uKPeZDzKeDPhAgS7V2Zp4C/CDJ9h1z+V5H
AOx7cn2FRdbUnmXplq0CdudWDefvpRyBHsef/hMBWIUjFjYVZbF2U82iwNDW8ABg
qV/fZx7Zzdn4p3eoBJp4BjLQpw38Xxld+0+3ocsiZC1ifdv/VWREa/LdNGjPIDFX
BkKpzlBO7x+KRLGISjBwbMQOArBl1N1J/FNXW+zAFsrCH7VsSMletD59/8+pL6Jt
ksUHu9/ntbkedZV3YlNWqry6RUc246hcuwCMFPwv/tjcMSiq+IW9LZT6pPmXVu5k
vXCzuQr5VOzfZ2BH73i2NXAD98OPvsIWJLCfaJKeRMtueoi/svO2SEMxuroUi3m/
NvXkRHN5yfpHiMdCX6QHr0jh7XjVhBf6TEqdGP7d/VUt7cHsU/KN+UUb/ppQLiUJ
Q0Fwo1BAO66e5NpzIgJCD2txBJEHgSNXEcp1HJEbgsrFSm6DdNy/aDZdEojOlnhM
pkTOfxa90stWRbzbZSFUYjfaauBUqSOO2o3F3gcUrkh4zptv84YN913ZdnOCH8T+
R52qSEw6ZYZh2RIPUW98HuK0QFchaX/NATh5A1kpSo6T+PV3YSkTs8lluQDZXA11
V3e/1FBC7EMaAX1ZB9wVfWOqN+zJeiB+mTV+9ozmRewG1EV0g8ufgHQm3TV3WSmk
6kyQtsjyIPBopwZtdeLqUCq7J+ChG1PhFqnh6Qnzmjr5iQKnM9Ir3IhdUdS1kFUK
bvUFnrvF1+V+Y8ByCDzQwvrZxBN2DF6EKypp4PVmoR7KuhJM6GUfm/Uzo/Gw2+jJ
xkUt63fwAZmFa9bsvvatpxTbSRO0gJ5HMjU46pqvbBOAz3HFohYNmGSk0QE9IZGB
IDuAcqZmCrr8qae6q/CfMdwQpcSZVy+D/SBtkt4kImBgmsQllA5BMleCcagZQUtC
olHhF0xZGtEXEMbZx5jCqh3+CxvGBvVrW037Gdr57J2wOvThjaX42kSV7nB5bhuq
hskbmrjtY2bg4j96kTB3DChoLNfVGnrUzO90/1wDwM9Bzx0eveWm8HdTTC0ISrqM
Bs7+OGQuCEUFQ6EbMekTqDDZ8UpLhM2DJvgvqOf6jWf/Bejv5GhF5rLcJs9e9dFd
4Xeu/r2RXlGQzvYevpJJ+e/2mV4oUiB5h+mpP4qBBj0Ig9i246ITrYQmlOB850jW
rOf4EwG4A37ySCDsbh7FQyhkxjjG8AU7hL/6zj2AL8oyNIX7vzDMS02KG/Xu5i6O
Ps7ZaBDwZmGgATYmwHVN7Pe6vzGOO7lMH9BB+9fJahVweWyZzyCnTk16yVJVWYCH
1h0bouSKGcJfDl4Dt3NH7yUlcIlKwZt9FkBnqtkD0ESjktgko0Vu3XULT2e/XblS
1U8Q/ild4D/FRZ5Hj9elS5ZzHAd4CbGQ9bJn6CaCgXTJev8ZV+VO0ioomz0TNCR4
XxIzSh//nJn6AuAKrP0mcEEk9bY8S3XKz4FKG1uEy3ljQmMA8MebP5iIaTNcOkq2
6UOX6i4ZqpXXiqOfd1MAknwmY6tp1lgcZaFtQ7Nch4LCRSJRX1aW7T3L/krjJtEA
Wpx1bKMpvUy6oUTUNx7R7N1czipiJr3RFC/agcEFYvU1a23pDaLJeuzjjSZK0e0a
h5xU7v0B6EwjmmosNstGvN4iEfm0cISKBVoFn3pQxr8Q057Hso4lrqS6qD4POnKs
hOaxn3Ggx+za4lxhI8yV3JqQ53mafpqYg3DQvFYgaeqHBBOyv93ko+bn+QKK0kjF
S8uyLbi36DUj1UYJH1z1rpuFOWkAwhQ/EKGkX2EMMrKX1PKWSTmPedVVICZUUljG
M4foVGq1W9tdWL/Y7FFaJgzCWoOqHcxl97r1T7GkfSUupLEo1hBZnVOFPLJrbrru
chyCBkoUX90oMZqv0psc8Qdttao0r/nqkChtYpyHyqSlWjUkY4iZUkegwdzulgAt
WIWK/J20o4vy6cRR7siXx5FYeJAAKGqEWSAba4R7pEcw8O5BWjn8QrN9KUmcoKq7
e3gDlfhJXKJavmzUBzp2KG/yoaW2LDXMSQZKK17MNe8dtj0EoD3fQ/G+MF3lZWed
V2Kxe1pedvw8Hdq88JX+Tjsc0fLq35+5VUdFriX7IqX9c3xh/3UnVWQNfJMjlmHE
Oycjro46wpMwAvwO4qyZJAqywMLOzahSDUTQ5wXJN/csF3j7kY9FxDAt6uJyI4UW
DBUi2IaO9oWW4lJ4zDjSLfv2waBnWz13IyPWCWvJCP4a6xkXM/+KjL473oPJ96/U
+VnELF5UMYN2QeeKUejRizBBpflygJFYwQHPLIipP+S2k6N/sY4gqiObFakdFg2R
p+OWGW0cT1fVrZwTjb+96FITDgEL5sZHyqf4UskrW97vpfiRiqRXIVlZi8SU5tE5
zA3x+FFEC7C1FGlv0gCG+INuk+M4tlhOCwSz9xPHYLYxWmN1G1d0MlbZb/wLeIBw
zX/gxQ7PXdSFT9T0kQ4S9XlZeHQkvEd/KjI+PO8n0RxEwI93GxWCRxMZZI458hBd
l0vdhmcKo2jzlaVYWSOSS7oSSCcYsRf1adR0NAvc6RPSdyL+EW9xJoY+lvvLp+rQ
RnoUkBSoj0irgkROO33cB42kUaZTLLQwWFWjq45/sClV0tNQxbIld8s2BuOQQu1Y
eRCRaq6YufSqgmEB/KSqMPwmNi/nEs3c1/1d3HU642ytYCW2n603YdtsergxGrse
g/hAog8UfXleKONUBMnrU28zzoba34DelCrep/nYiqQfyqAoRzhrwA6F9Vwg916m
ooOCdd/yukkX5ZeyEjyODEIKvrP9NePJpb8mYVC4ZPJrMFD5nVz9cIqa/VFaHT1z
gHFvKi1Kg0hUOfMIilxeQERNyBJmJHt3TOZFtG3rvKVMtDVeksZU9txvUFNYafOj
EeWgp8Ucwry6rFKbZCAjh1/+t/+V1Zbi3vVV1NHWBTvRttn5uSuaqCHGpVfb/Ak4
FAhneWL6xByMJzT4Mer6pXHxBIdnxbbFXgAiZeOdkV/aTVf/N4sOhnhijBGbFQKD
R94HLk+4CG4nhH3gtg6ouWLcFJ8hfQe/qcyxM+cZ3tpB20j1FixTnQ3mXv5Syrmh
asKgCPllKrl8J01mWsWifRyoCNIJaR/mfGztb11DaoXyv+e0V4a+qu0j2WR6Blcc
Vgq4tNKH7ViaraJl/HkfImX5pNwLAEmGC+vEwrgGagi8Nv1U9dxfTknZQJ6bztAw
KbM4tssIZGhp9aYVYAKR5qU6GjNT456xiIAbTrSI8y5QZRTjZH9Ts7mIlfs1QnFz
nJxGrXeTJYHS4adI3e4e3Gh3sWeNWTumNuCcRYjMvpipbuCshQ3u8IyLFeXjbQcn
9+omMXpkBAfes2ERKjKl3bhlhOaZh/wVYIidYqchtjRcvCX2O0NoIlCqZ/zbAv8o
Q/LQ3F3TTnCmdgt34DL58kgAau6AwHK3u1YS2nnjBpANHVWepokbJnrrbX9gYf1x
/B88he31ghOkIMDKVKKvc0jKeIL6Ln2UxD+9sDP/WY2BmM6GwDjmAkqeOzKzJVPL
yk/sIsrR8l7VaRduqdTtE0wmQJf+N9jUJTMHUOp8h5JPwBfByvRiF8efnhra4MoA
50P3WEAlSaqG+jpO+VBwQWZOKbLi3dh2l8lIrZag5pgYKADjgueI5M9o9pCYdJVt
BxHNV41ZVcyS4zGy+Va+26OLfNcbqihMhnjm3Ss1h2xoVt/JRg6m1q0nJm3tV4PS
oGBe8KGretLrTrNUcXal1dYv/eIqjUYU0YMkm0Y2j88XvHznTia6b9D/vRstnn/r
4Io7sQLwLtCYH/zIVCLGAI/5O1srIosG8if9DRWXVvJODpWzJJAzva2T1rmAz0uM
G/2+G26EVFr30ZdR17QtQf9qOZpNpiyFraohHKTcH5Iw5T6Yg6EMQfu7nAXRLGyQ
XO8T42AgRIZRs1PuXqogl3OdZHF5MrcEWn7iAm92g14bBeQdaD75l0v7fDZlO9SK
adkERgy6mIpeITwjhLFA62DFvUvobtO7CcySEzR7htPJwQ+zeAe4uNLtMyWFywwJ
uJ4+VlxTUYuNo+U64pIwngGOiDO4E7izxyg0+pGkD5vxjmk4dWMxl3qZt+RvZByt
spndJ0KcHnmIf0MSfr6HxKcXsWIl2heQuIOl3EvI+rIJCCXkle2mIsYES9uCIjlj
cpor/ozka7E0BSqV9EjpwSKSE6SjNTi8HGKurn37dOOnzMvE4WtJYmr3ySkLlxMx
QAyXh2T7a1lsXkt1MYwtA9eoKjLojw5jFZ9VbWBWRiBQKS1y6pCUps7HxQURj79G
o2PtqhGlW1maB+PKwN1RMRbcgBxFfoOGEqA+HSzuNrQhDXLw2TfipmZuBlyPlpOE
GOUEziwFi5PLL0/EZjWGBCz6cCtbQryXUltDKTEfvaPcU2XsYe1B/tn4RXH/d4zQ
LSpU1/gNmKqb8ghEAR/YlhmlryINo2EVool+NoQDnAeStv+aCGYiSU4pA4wyJI86
1NyinCmNW/Fw/OMP6ZttCFJCueWsTsvP8Rl8R2/niObliqCBRJYYr3CUW7JD16D3
izusjeYnR13IFJZ+QY3w+SVZTE1Wk/Tl/vwKod+ua1Rsjl1SlrIeAvXlNE0jCG3I
+Jp4Vpc+NYyFiJ03suvZbSOVOaxsuhXvBsiPbid0axzxa07nGpOsBHzY/G4n3SQ7
rLdXCwgt6fzzcUxAt+f3OFVxaxpsiSLIUnQ6KsZp/GwvzvX3ei51ODESclRjxsnq
cAxNzYv30cvZXnkSlFtNrblKUzie2egb3UL9B9O9hfTeqWGMYW3GdtWXe8kjTfC1
uWhZNMn4sn5GNoOg1OYg44oXb4AaFPXuJHYe9aotUiRxxVcNfM37MSA4sdhF/X0w
gJhSlgNrQ/R3VzIjRBTLrOWYTwUzGOOhAbamBJvG5OBkDePkFw+gwIiBB+Is5iKl
TKKzIXmpuCXCobvvPAitlwYosPiwqOBz0GpDzI+7SOKFf/WJ0jMipD1Us2HTe6XL
4OS+FLMtCUBU7/NhwnROFptVaEj6mKBN64yHxEP9WAx3d056QQk9QHC8wTYnvmFU
KRxNfTDZ5CVX9w2q5Cx0Mllp1hWV/ok7yxvyKrMz28FAj4pphbK1b1rSqOjM6Se7
rrUiE6/WM0PzgqdKI4XowignCIyYpLLfJ+kJSGEf4RgIxYdC6qZZkWnd30aqLqy9
F5r58laigi1NhNTJryEQbJoMrS9QxYNgeaIPsgxTNmIjEnJnSPtl2nbN5N3qScBS
rA5PVlNnpyvdHUY1+pAnBlbFewCUWOSKoY7EOKfWM+AkJAOPKNL5MAcUVm2xVRM9
rk8hYFRXfj1wzS87I0S38neAPgRIZ4foVoi0kyHlGP50WgWfwpQMbX3SZjML89gZ
sYa3SBCmwWzDKtoLTYN5DOUGvLBF1+tJ/b8eMaMQNFE7FAu+QcpVNmQqEvMOMCpM
xcDln9czEmJ7jSXynkEZC8jvTt3qTDPlmH/6MAR7nn4kfo+fLc34gsqlQBO4amGM
P2Ua+ywnoTTUQKyF7d3NXZhql8o91Dw7xG7Xi+pGsozhXIulsEk8lyh9J5HYc9AU
pEAYoo9YrGvXubZHSwWL4eTEy4uq6K5ziRt5lT112dU3Ac/VAu9Q4F5TrphTExf8
W5iBmyzeWA5ypQ7iahQbdLG02GBeK49XxYTjI3DUTJM1awI1v6jnf1Z/STilNM7l
BwQnHLkpthPAqszQ0B6f5lTwb1tCEUI1o7p25BgDL32U2VYl1sdqVk95rD2QBYDP
F2cwQ/1oOD6apLbvjGK9IYzQL2Ftgyn2AafFuIUbKf2fG1JjmTXZt+2kLcu9arU1
Ai5bhgV7MXjXF35cNkUShaclzNQUrTS8AQtcEeBH5kn3DcnBTpUJAXnb/M4YfeJ8
r0js/Psw3OyatBaiGupTWvwWQX7zWUn6kdg9gvB8E4xryQLHfKPx5WYLHk9g1GWM
hCiIOTq8ilRd0N5Titfz79fWJzzDb+JKhgVqT/3JUWjQj6oeXqlzaEC2+3uxEPJQ
ljQhaB7DN9w6NKj49P6rPveoS+VL/U156eFZzKDy7kvDDhfeNUeSUThhx2qGCh5b
aW7c5GVKpDwEqeL6QvPHulzNFGtLgmJB5VsiD05WNXRtjT+QbGm2TCm3fmTRylGr
n8Tlvdlg78MlirzK1+asxlaJbKHBiUh5KCyrBiNjB6xMpEjGt/aMPlgvQfvgQPvL
++jkmytZlXlClnFpOYrmjbIc8LAJRuaFiJ6OPobhhE2FOcoG3Bz6LkgqGwW6uzCX
C57ZgBsBcWPLT7rvNq+0HG0yaOFQ3aWaqfILL7cPLezPp7lh0GApdEf9WboVkcZY
jAdJT+oC01DehvFIslQHTWVn7/Uvh5cBt22Vd0QOpQ2XgJ8WFOgslAyjldEFLw74
tad5x/VAx0N28FuYFm/CpRgI12/NFERgHrkY+SnmBoBl0P+5BbehGmsYAt0e779o
LLEccqSNT+MR9Xwt9ntC2rrX5/YSEEq4nYLG5LeHnO0lKkkZxe5NSYWDUHyVV9Q3
/GJoQIV4ap+f+6FSmI+lFoutoS4GpF1Z67ppxOkm9IZyIKRm1n38yw7TWm4VNDr7
MRYhKscy01g0ZYhevOFjZjfnGp+LGPFekEsMXsBy+556uVBIEY1VmjDnzVDSBnjL
sDKp8op6m/RgbJ4+4/rRCtTucoHGSMpVCaZBYkewYe08ADx1Chh8hHqxU1lJ+dRW
UUbP5mByk8ilbxxFmk2+n/+CtgQq+CU0wgEc5SeC0rp0Aa6U+XcUVLImqzY9LtnR
ND/j5XLCTPmYwiucnVjXm5ezfjPTjXkzOJOEWAE85A+FS7fuZfhkP3xT8rs61DPI
boPrYZxM8j5rDCuEtdra0WzIvHy5Aj8DT9l6D1RFhHcqpvUVC3o3JkYJfVa1TMGl
C3v3JJ/U0zPrhfWBEs3Pu7QrbRqEKZpe6W7YjdYZSzxJOOM2DdhQg/v0POvC442n
DZaWzLz1cprzUUTGma2OaUEBajREAqlPmLTz1Z3iNE0CRkJ6a1jokwwfobWbdqov
LK45EkHT3B2ItsDIn78tdixAGy25FiQ53P5rXAlCvCO0JGMPiL+x4xMjjrz9pr/r
VnHXYdJ4LbhnxGTZh9mJrgD04bqLO0SrlAKLFv6LeCbJWa4R2hqCWjHlm3W/brTt
td0256rw9ce143sUsuzJ+MHKp6MTm2kU26MHM8HzySi/9iiMVTsK0aSkhgEZ5aNm
UEc8zDNupnQrnKmJjJmADem2mBkbPr5Y3G6oMHnb6/EtNpRpJNhs6xxFYrqXH3Y4
gkLD7Gz3igERMQymjoAalYP4X+AWUaf/3m9y2bH+5YGqse4u37jnutA3eLVeAiDQ
sPl549ILGXk7gEaA+hwD1xla9PlF7uBpkaqGyCohQDlj1kikuNhyCroZTqxrLfUS
7jsG2wVgBSiM/rku1Ywd6I2X68feZMr2GeVFOoOyeJdiDiV/G6OZuILhBekGA4Fu
mml6dxl5vKkLVdi0LfP85t73U6hIEFlEy0IFCvqxwVgQ/+4sSVpjqQNupPxlxEVH
Kxn+FW8YEpiA3AuH4oAqMgouNT41jWw9reXcIuLogkEKZmSyiB108aGktgb3wv7x
0heYvqM58DrIBN0LH1J51UAyuNDoEwt1la4Yg7vEJpoD11yCHfdD1whdhu7dzRaO
DbJvMYtHxICEnWlawxfJ452nIl7s2EnM/23MT+Z/zysFVsLyRGxlAxrjavLIZJW3
eTlUAevgzUbpYXTe8jZ1M74J/l0rUwIpApTQeGoQfTAsgoBmiNQeJDopNeA7IxJ5
nJ2aIKLBrDP1bBuu0/8ZxjC9tIPC5dsNc05HlbhiEGMtm5tVS380mVtzhcUL/Ww/
MDdf5T7VuPQBKjQT+ErQ1tld6aOICb7g1a/5DhEwrJNLuh9g8wzPDRdXykRZSRNo
/3S6KZfviFk8wq93BgWd3iC9qMAVyCtYjtqFoj5t1urLllJgQ7HjhQr/kFiWdbV0
CD9S7enSQaJGyTDrsc+BqyXMknrw9Bjc7JbaPTaelRwQqsUFC3nZ808a8abVehkn
ITn6UF5b3ZZp/XBmrKkLDjBc1RxJ/Pa1KiccBHERc/QGo4V2feaHsmTbF4xr7aLb
J7zg9kYFB8DL0D/7XauxrbyCZYFsQSY1Xt4RMflZxyURF3FfbtZd/nN8Jq8nGyNr
U8lbKGxcE1Z3avJxunrV1jPlv6fr8a2PV24eelYFKAt0gGLxasBwZj6OBRKH7/2B
dXkiJZIV9Bp1awJz6pcSH+JCXPPdX3QZryhpPgIEqCwR/lo/F1/PmeQwLMfeTmUh
caGbVmG2irbtnu7znW663fnXh3ibdOrl6C9rdU++84gXJI6GYOtZhe36DftwmlSV
GXiVljwTK0aA5qVRcShVkICW5bp4TxZUp7RUyfxV00+vIeQP528X66dLXqhvPjWd
PT0qSxNK4Z+GBKjo/tYAGROzaKuomYNHL7RiMDJHQwqXeBoxAg1I023Ssi/L6+Bx
nUv9IP6ikFeVuodUeV8slNtyqNKWCjY7AGhRXsCrGjFEwiV65IRI9HYhxRvm3DiX
5C9KDWs20LfdGTJn9RTqid06QNgIMGc9wpeN4qDXZW4ug9gsIw/ZaqbY1lke4je1
9lfCIZYAkHtuCGHMvAo3CQYwSsUnFRnpsHqw0cxWrWmyHStt9UvEUOOYjTb1/dq5
IqO4Bd6oR9wLqMabRjSMKXetzrKcy7QctzO5qVgWAy2Z/G3b/wZJM9cFN0+C7Fw/
NjymFcn4SfSbtAo56I75wDwJubpyQlmDGYRXQI6SD2UdQhBDzsbhjMktps5b/2v2
rHgMHsffZlqQTMuVVvbFsFZn7fWRPWldBaKVjp62bzMD1VX+4lnfjbcz36hrfRMa
2LcdaenVP0rhMGw1yXLlBr/eWZhuKgDj1hSDzQOfez1KaqdHmjwIPUOoH9TJGYtw
eGFrqogMB1yTHh/hSdKWC01IK64fi6nV+efqAT42ykY+noe5sVLYrY69bgFppxWg
xSwx9AXHnEgYQh3c26AlSJ3/2x1cNLFTiGzzWwMgY01GNfz2jPM47BZ5KkBjU66S
dou68uvZUS4xofV3Kq43SkT9e6qrakeW/abNXXyaeXsOsGHmuyPRrrk3tKn9a0Ci
BVlNlSuYn6RP3ssVC6b7esJ0QOAt52AggGO40QIE/FNTxdvubdqtCvtSLDjYHCx6
+gYcAQNJzGgvo+iziqiop35FmkNcdFeySyUkHBkI+i7nFLaB+7AyFg/M/hHgz5Qc
AXPrrYDI5mXqEuFgh6weQQRgMzccWPcplTrnr/qSNwayF7uDjy0gb16NY3J7ov8v
N7WHY/mYFZq4zFPyUO/uvUT9PYqVI8QEIYa8GOK9ear6leNzY+jXI/b0dSBNyqDI
an6Y9/fxvHBybPX12UWKnYrRFcmx5lLO8UuR45tVCPUwSKBzOIhUE462iCsXvqqC
c8T05kLmtuqZ2tuKAMq2nzWdBjKFFkhls3xgP2igyBF55cczQ/m3FtmB9LI2vgw7
3wsFcVmClp8aCcMEYshTEisLoMvvAbv0yOpMm5NTfuzE28GTX53W0l5yEXR741/8
3uEuI+5jq/WvgV3td/rZi1zr+jkpE4HzhgYWZWzw1lf1hxo/K6LgB5BnDF/GxWja
GJtNFvV1LdWNJCnfny+K9NyDwZv4SDvtHiRlrc3+X/VuDIJWmYOaSoSS6YMb+L8T
+769U8W4Thzdnd75TDP/QjbC9jI4QEuw5Mr1dO1fs1RuKrZs+1fBNdHg2N2dxSZL
Bwgs6r0kRW6lrYRoB7H/OERnYF7pPqDBKjY2cm3MFt7psvenB7TkX/oGNwwy6tqv
w59pnF2M97v5G03cGcdS1nWHYQrzyksFThoNEho/aE87NOC880rEEpJL0+C240td
h3vtBHHUc4BM1cRNjsiHdVr16ZYBBZg76CgIpQBGeWC6xiUeWZPEVV72sBSoXHU8
A+ntGYKykBEBXJH4gtPEWpxPy1wP/hLxa6DFa0+XKavcpUELMOZeb6aWydTwXull
xFYEKHzxEQAeFPxS1IkSxp/ADn1r3AGA/l1M1yuNpa0iArayzLbaU9TAhjIBwENk
vge3Y19wFbSdBoSvKc1IxQYURLqxSFbRNm5A/C5I5sUH4sOw6Re+kja3zmYMIudv
zpol5VzL2G1+AU5rrIj7wNoDBFEwM5Le0fWSQo2/EuBB391kU3fqJSNPufAchY3U
E5WhoZzvuvSvwGhFdka/Ak2SblhUexq6Dq46H6VOSvYfrOZ+jkSZW75De+TxUTQy
szChg//Ujv7I9IjGvkibpAr9RBXGG2vvXiaFuP0x3WGytCtEwQFMWsjoPkLXRooQ
izvdSl6mrWRxghWezlcH3BlFRcPWijdDbm5XYSiNfDLgN8i6ePDYtKSVTqUnSIba
Wsn+0Ctg+GcYzAdYrQ9EtOlm5Ln6ftIbn4YxYdYxVcM+TUPIvxEHCZF70RGGzmSa
WGewtY34gFZ0O/ypVM4ERM9Yut4XGkA4ApPlzIqch/XGQACwU2gRIZCs474qeCXL
PdNzjnlDg+82OnWivjj8F+iGb2Emb9GEfJE+TiDJW0cfjQWpIYYeH8ILES1fhAU/
/pMf6Smwztp1c/uaeQNp1YHaZ5l+t5sw5UjRKv8b/jzIRCQOt7jPuaE6jXXeoH9Q
ATT9K/jI2CG9x5iU/vnTONppkaLntLQFqMLivdrpnM6uS36px4dHo8m+GQJMmQhE
e9e+/zyOt64BJ1VG5JV+zf/9OX6U85P4Wc3HTM/LRJs+n3lzzs+7P/kkK0pYZu+w
t1Fyi39xd4UBB5dt5dG3qN3GmguguQLocrVxzHHlGAuQOSqRIMbkWatenOGYquiN
doFOJhGYHLgK6X1i1QQzP/AgGp7hqZQRGg/eV8kWOPPtZQnqb1syMTurbKKSwnKd
g7i7ZFLYAElgLDW/h2F8hhlkzac7uyKq0RPm3XF3V0BmYAJH/QN1AuRBtUWSCi89
8xfxD80VefKVV/aR7kvbNU03eImWTbpyxswZLogHA6Q6v+YKCcKyJwudyy831atE
Bhv5hRGbPUZYFskhr/d4M1H/2RR0ft1FZjUgVTpDKLY516hVxbFKkuz5ePBayTXB
Lh5LAIR7XKu1AqVbQ1M1K1Ster/W1CdeHEfxq6duqw2gKUdf5sZEByGl8IIXoVh7
QawfHA5WuXJwQvsEQkxdBZvjEm2/LDAGMjHpT2SJkgH1M5wuhuvkmbAMFWm2p/Le
BiZXJm/LCSa593L+OBvHKZnCawgHRVKX/nn1Pd8TPAao3R1rerPdTPYzytqG+QzQ
h5MfwUkP+uPfsN2ON35wCsUvIPBGMbu+g8VzLO1TTDLk4K/PxvjLjzZk2ag3iN3u
yJlO6WxL/dUSiPQPlbO4bbv2Y1NTFVlDWRgoXtQLRIPsLGc51gItExn8BU+FfKBd
JFJvVlpL/o8vg00i41Vykh5xa0wIZ+PcWlHoLut8596JdK3UtpbnM3fGYx+R9riv
yaoNMwtrGi+pK7y3LM+Z1xFGgIHhzNnHVE6DQrzqWt3kkY0bck1bbdgcejh0yjBx
I26699r0m40s+3K97aR8GIT3brL437Ci4BWkvqQFHkHQHyS8JWFqsKx1BoIMmDEf
uDTv7nduxcM6XUHXYXfh++MKOoFFM6sgB2Izj4jH/0EKmz6rtv5J2VOyAaK9JOKo
GnYjdPt3DsVOdY6sLZzDh8BCv6r11Pr1kB1iCXnzjxgOOoa3u5t1yJaQblpKUux0
/LFqsRpzhDC7rle9M/S1+Y8WFi7xBHvmtWYd2Ikk2/36yy+hO33Az0mQKeywYryw
IMguipxjmk0UNeNcCKLvkgdQcEnpfr8MyduvaFB8ITCMQaTOp9Viv7b4fLc73o4u
j0nuxVCUTMd+12hrqz71gMw7EwTJdvr9U/mB0HHFrHiSvbfGztzEhwQx5dgOnIZz
MQ4q0q2UPdQUBM7R43Q8SDi6LZPgF3c7PXxIS8xR8XmNXXq8IhOxSQCdqaIpDk44
vOpYkgNf3seXF+qkB6IsybBbay2UsfVbCIu6VtwjtrPfxDkkF2AG/gMjeCPPJC6q
XtMrCWkR4wA/p586tU9nw3WLlcBTfIrzMkf4Z3I0UAY5OTsrefqutos16YwYAPYT
pbxtyMWsf6XIG2yDC4GFMC3/QQJvQJ/5F2WbmSGypGnLVanS2j1CtHDN7SRacgTo
tJj0tXfq6r8OLtlc14UY2P6Tzi1seBSleJKMwrfA7aw8KGDDKAruWycWpokdEXBU
l/6HknvCQjG8zSW+Af6ylzNAQfOjcJDP56MaAkEqJPFgwhwAD06EvjFaVmmK4phs
BEcUntQwGssTUTQ1d858a15joRPayULG3/u0W2du0tuniCn5JD+GhEO1BBt2/hTQ
0lwRP6XWpXrvyVXDZ/NXCHj/M+25ntsSLQwY1Fi5dVmWt2rrbeC83Aw6mjxvsSbD
Re72FgQuNZ7Of8yPQHtgQvBEv2o4f3N8fzDcdB/wv105yuydsLhQuVUJ8n2n+vyE
Ga7xW01pyExdB7UjM9oe/s/6Wum6DNdnOpKegSCrFFL90Ka/u8se4+g5N4pCJpAW
PJL074KcsUuIoP0N2WQRxSIA7J6GYv5X2XwackwX7jjWxC9zBn3rr/wjj2pH3Ass
jPTG3z+YLj6HG6NcDH9Ds/DenU8LupB1//pPgk1HHUwbUBeZO5vjCc2wj410FXvA
EPSVcZYHQcaKChwQbjuerwDKnXzGud1irgdUfLf298SiCM4HUWz5EWN558Bjj5zJ
QzLfqfPPzD1Qtlkx1Q3WuoLP+hkZ6RB+nkxceERvvZsMx666Jb6uonQTo0G/uHZ/
GHq2fCLr0BhQLtDvLvOtw7iW9iEIEI4TX8/WvCUtPkxeZO9V3GaDpAymdsLbM2MY
kGSXnm0YvsiD5nB58Kq88rRQrXs1Fz0bzJ6MJlM95R5kYq8CJ7bOCa+F81dZytzA
jxjs5lqD4Dt+vDsJ6cbdUxPF7rqufO8ZyB/xHZhAIJ+Laf9mixS0eGYt/GKEeG6V
B0cAyiVBuJCcY9FwD/NmeJas7CncaTgV0q8Twt47g1tMWpPe1Ayl3iuqASrSLWto
z/yhzySFcvvdYMJ5XnvcevMqiOwd8XjEYNLWe6pqxeNeC2Er2K1fU2n0k1qZdRBb
Xgd+L2/qxqqthxXvEZEWrl/NshOVHYVRf2NhZxCfd4dazvSo4+UvFC2/uuz2/5sc
i3ZiSpUo9gYU0lwU35b3cN/TGOnioakOFkr6VBTBc72HKd8u18MTk22GRG99LjwR
GNRP/mWmCqWrshYhNDA7drphC6n+0MWV2XMa/Jdzmv8caSiokMLfaz9s14ls6k2G
yxVVxxx55YBOunGPm0iw8aWURC4NjSu2BGaXEYW/2XLbN7I5nk0Vw96E29pKTtqx
2rG1UpzdrqJ4oBspWalxwyoK38+I0gDa1PAwbs7tc/XTv9/knp0c55U/fbrMyTBO
fq5knCegTONhmWuRGrcDuu58j2B0+XJjvx3GCpedlF7Mr53Vh1qEnrBkBCIVy2vZ
++jvQMv2PiVoNfjb0lToWmYfXvpD1kVjrp2wyb64ySQYdd+LKndBc21O3Gsr6KMM
B+qtBsnpOsLMWsDUNlVKD2X+sLI4h1J7K/lEljANCS7bFnq3JA5tfH5eD5JKiiBT
IBAlWzC0HfcpRFE0X0qOHec+CLRqU7YVzQRwJ3aZn7JqZhIz/AfwU0B6zPKKheNG
lvyE3b0Jk0M4UexkHKItabhAla4XDTDR/VPkaGt33uUg/AyNoFHAlTLxk6C2ISZA
vsDUE+EbJnpXazczX4i1g5aRLofcL0JsuDrHwSsOmC4pARPho5QY7+8GKSKP7peo
QB+d94nZtJPPX+uQ4yyDITccLxoBuq+paBeSwrn/z92KgURR5NDq/hcU7ILoUEq3
Ewn+WLf1hKMc+G5SVYKxhN6fJFfP60pT7R7gWX9qP8P4Npgza2pF96T0SroDJLR7
d+h2RRRKERQ+2n4sVonisSppv5d96VY9hgtx7gJBIBm+tb04SgTsy0oTv3DhLF1+
0Iiz/V1q5CBkJA1Pgy3oFnO1P1j9RsljpXA31WYOq02YwAWKCCuVCcv7GqeweyNg
eGHOkf2im5p6kfqB5KlFdt5DjkrYknoQ27PjJSVtitRJQLCcW6qBtH6LBAnZXWIw
xc6KH1lx7pcGdyz1tSbvkrfnfeJekq5f53izYK8YOM6LtgJ/e4SBYP1FHoPcXY/j
PArflh2bTV5c6eULTaZs2u9e1w6yXrZnQcNF1Y4AYCKHFxcDkLJV2S7eXc9jVYQc
dyfqj9ClGdGf1wtD52km5Ty53LokKWfIbh4V5IA7fYPoXKXazKIRz5PzOElY06nI
PHsjuf254fzoNjXMLokcV79fLAdtSqlYpQppGdKeib44hLDA7ZLo5nmplaknElLE
+/u7v6p8MzlDLi46/AqCVFk8NBklr9jhnAsXUoiTo8xg7XDp8BbuHkg4eg93hUpV
1XngEZtAFb+r5UyWDix5ploYraiCRAkmZJqFJlNPDIpQwEsiQgz8IBw6k/6sllPZ
y0t/z4MHIeN+hNIzyCUkO0687cBAh5xHaQ3guLkRluvKzmHxjoOoIUzZXoqLy5xy
xZNLYxCZW75lctKRmC2POZYcdamaJC5qkqpxe+WWUifSLi4pt9Ss9EFtyFmopilc
5WxwSMya69Y6OFyL+oFOOc0LX/lAJTIu1SYa+0g2vNvXXIVcrlHZxxmymiK/5pXR
VrzAr7IMWQcIS0TPYb//LLAAT2ao37HZfae6wPr6tnQDuBY9bd968LMLxL1B5xOV
Uf4H2rMvqOM38vMqdoRjdHxkCnsmh33iZOzu2lEVLGnjtrHoeGQqdkhxZ4xG2nBZ
/fASvVmhGCtOsCflW2cUj1yWLU2GRNfEjCKM0/YLkwSeD5XutzDYLg+E6LCX242j
I3J4Gpicbo4Z3MTY1F2Svw9q7gbb4YKtMEkfLIb9O2Ya3LRe4k+yEHY+cKhmAI7O
HEDIgtFt+BCTbEQIwluOgDdr+Vq3BIVtHvgbmTUsIIzPEqOHdRAsNC/xi6trBSMT
RvXzuU7rxVPdWYuNVEr66FwlEdbMvWCtIBjqR2EosN7EMiGkKNghBwKwlBNS587S
9ZfmN/Ke6NZcg2+f+q7BolWWn0okT9e2jdNw30ypEgcXgI3sfrFyY0zk/C+4kWnO
hLojZwxaPNr2465HGW1es/LCMARhuLUfR/+lzsOMr/s2lI5tZEvSBOaZUR8lbq2j
oBTCRKl+lSLwoAY4ImUse4dBK79wA64CvktidDGghjLj1QSQ3rONpzaZPdXdweBG
UJlCnzHW3tMwFf+ahhs3jV2CqSFk/1RLE+dqXaLwck9EhvqxRacH0fle8khzGhqF
o7eRbtQSxsWprqLriLj1Z68RHv/7yn5NPq3jyB9mmss5Ora3rZuetZh7o7ToXP11
H2TuV4PxtkIyEgZ95P7SAsw8Ilbj/eh02TQy8mUuDC75408ngk0jlIh/cHeVXCfA
xelwSAuWTuO4BoSlbGaS9wP4rPndIZY0XJV3JrL1y7wo7Bs1SGT/ewkT9JNMaRVo
Et/F4/pJzzQhVndiMfClyKdviDUrTQYHf1fl47+Tb5MMvv27JmbUJ2jydgLX8T8X
VN7aS0VscZPjZQ1wn6JPAngdGeippgUs5nhyFhtbMwwAG4gPRk5XpFDzZGbPXlOP
YbeIIL+/BELwigfBAf77DJswSKAknaw/Qv5+1GL9vamdZ32CvcB8wHLbZzNNiuse
gIrvh17CFng77Z3sVnJqiJAL0TSA4TsyTvRLHrAWqTNqXtRmW3f9pqQ9CyW/5v8G
fWzdvZvaBkNXL4vM5BD34dnQk0m51gkcud3OUCYEd/bTEatyFPmd4aicAD2TVxfU
9G7ib1j2Hs3cUH48NeFt3J9bcdmbJnekzFnb5sr0/XBgkZXkUCEOeaLMzzHo4Zss
4lFhJkFJk/Uioa9TSDS3KvsAMbeDRH2sjhMrXqaQj9q52dZCCWKH4lMGOk8zFi9b
QeSFy5AWjK0tGjyx6hvh5yLNtQoIvVt7XxQcY4fHfncp4NCHoYmE0P7MB7qkY1Pc
S8Ca1RJbZ1+0XINCB6pvtBa3CcSZhP0EUrdu5qqFfgdpuwk4DebssUsElEvKbjmm
KAaRFqJg/Q0uR+mwzagz/hpwsKupTyjULs1I/W2EgMQWV5Xb1BWrXBbDrFgXv73S
RYGU37H2acbaii6OwoHgpfTqLKAASJGxi2CYW4f+oGxlmWYCjwGCSWl0V4/V6msl
RCuFha8zLEXNZe6ci4qQmZsHJel73IAP4tGSz4i9XsAkJcMeeKBz99wNenfxLgIj
r3F+P7RZchvd5jxevltYtsjhaVJYNUhXySYs/T5UAwcH9qxQD5R1Ll2cj+sWhVkA
JLoLhFPf9O85zduEB422XHOz8HRPK7ZHwArHGZAiZ8vHPbeXAJlpK8V/6b+AKNpj
Iok/SYl5M1wrLAB/RMOyCbOz1rKA/rkpIVWTC5UxNTpDgbJgmpJv347cEzBTJJpQ
3MLyKPsWLP4o5Et7FJEb1I193nB8bHTCnL/N8nd2/kHTWoo1sP2fl039jf7ZlDAP
VxCAIuq7Qg7eMwuK13bWVD5wjBVMVv94YvSROXLEMIFUaODEhKpgX6DNiuuIPgA6
bXLOr7ZAyfLnDa+b3vh9YXYYKOQK4yLAY+I7rZejlxM1y4PsioDkGYstYnxEAt9N
MInWilAa6LTkMcA3u6cF9N88TJG7p9J0vVZstAeU+s/zGrPHcDA5OzCHXXIO7ofF
4bJoGx5hkfHYx9t41MCKP9plp/APuLSABQarkGLFK7JYrWSlqst/RpANn2Wn65wP
etbyFAbq3F/XWeKDlM7/kZQ8sDVpksrDMD3J/YUWA/i4MIVtffJiHo7GXu1qfLnQ
qdCVhhR4mKI9MkOl27TS2riK7eViOpxwl663d60kljOgOUqAvG6740RWYugKMCIH
UpgcH5yj1j375XLLI0dzvWfMGXcth0eItO3jvi469nEMHCzeYALozji0UiA54Qh8
pTNXAl6T5ta9+cZdbqdSW8MjPbXCRehyzhAHWTIe74qq5rBAUiNOW3pUu3vBG0tm
qxi6UMyMIfSxftY5FXrPznMqx1FISPcoH1dTEuPTfQNOtMlQatH8NLBOgNVlTCOU
fKzkcwfAD6jFu8t12y77mwCNxSscgcfBfgeNzP1DUc108vIyd1QctX3ylCyikF/C
8Ez9Hrj6qmlTZc7n3L2kRhkkJVP5tdNZY1XEHRURe+PdMyZ2Wfrpg/Hw/CdqaHmK
DBtYGQu9Jso4ISdMp3BQadCB0XS8rYuvTvzWyuDcr/l7GPyGDxs8Mim1REDMQ+Jr
qa5nmwKZRp5XvEiu6/FOjv4Vf4QBF6+nLcxctnSPc65BMvwRCsi7bg4DoV6GPSsN
KqgTEVaUKDTEc0HZ0Ot0Eev9s02k2pc0VoRapo50uENxEEwJoAuzXjr1l/9eyBr0
khmFm3QidGeZj13PCtnJPJNIzoNiEh1xw/ZgeSFeHzODUiRC6XzIKyuLuErBkd1f
bQ6Ux1+FsDy8yqwyrCdjqpSmtGlUkBJxJrkkYFzafLTDOe7LBYlxLjFzaASHJMzh
oZCHtHhCEA70fkCB7HQxIvprvX0/Xn+WxTx5hehG8hSgttHC1Sr35MF48MfvsdAl
JmK8b0MGdp1GGd7iokLk6XvdqqXYw/M9sAar1VsOhmc159npQ/M6EXfdqqlB3qxD
WiScpkH+Tcv+MmflRDfwoqTTplMmDd90UkiXQPlCgV33UZQH7ZdpjpZAtxwKC349
u8tgxxKbUolkJOHbbFSXmgf+J8g/2HqpGhso4qYNiHgZ2pvay8j8a65S7hUQQHw7
BvBrz0yKP3HkgallW4Mm/YHdkwnfjDQ5FWYzpOX/jyHGld0A/UBP/qA1rzPUMAKy
py0s5SSJ1xVlk1q6hkfNl7ByOVqGNDsIG0PKjIIWQKT0lxrJXjVwDFMJYlS0deu9
mh7uBhEgu6VLATXdR6JTvr8rDA0zcOFFPe5oOOpSR3cV9Z5ZJEDAaGI+bZPbBEzr
du4L8Z/KzuYq/hsfU0Guq9iFCIuf/tQmtiuKRoLVRHkvlzaagnyA7zHOD5DGtnCY
G0+ir+8fVYPAIJkbKKJYBH4/qrLzXcwgXm6YbaDi0yODoF9lDmZtik4yzoRhgH6a
iOPAi2YyUbNPinsX/VVnD1SFEIEAQe8i7w8rlF5X8jNGBv4UpmIdmMbZW946T5Kt
H5uIKwWfaWBrNxh9hF8POTP0yMOCyTR5UcsCVcvLMFJmSD0wvw4IeZmBX2SL6TBD
gzWqRZPr5AIMFYUlbokU8f7PZKZaJeoHcZJTQeIFrES2ASAp+G7P1gOY73LGRovD
eXVLZN7do7emQoJnwB/31A0g5DJw4Xe7oQ7ZMygZqs4zd3rpVKUyHlWs0a7d3gL7
2avzKzA3Xd6sGI00FK+vY45tID3NJt1BpCtoMxvU36teJH62T+M6p7CCQfI2YEys
MENH6jjUwcaxk/jtFfOhhK3gL2WfmNk9LVsYOlW/Zh3zRe+VTbsudnQG0tvJxxMS
7XyJZZ0Vb1ImZM8Lj9qDzM16I7GwsnV+FjJthZeQdwFK8tCvEHhMgcqkFcdJmE7n
ahQ8xkNz7GLwU9BDrTgB5lCHtOTLRuPArQt35LXXUI1RgBK5EizpdRX4Pqyx2xtp
dojflEmzkeauHTIuYkrooMbcUzCPNSRhIwTR80xwdXMfVpzKVTjqxz1YaLjvGEnx
B19tsb43dGRaJb1yD5jeq+VDkJPRSFslgxRCNMRdiSdLoUWWa/EgTokYV2X4Te7P
0eCWs/Kw/AGg1r/b4cJ8cvCjD8BglkJpxjgDA0Zj7ZnYLWIDhHH/zAtypVvE9Afb
o7OM1B4ck4pvPfa1uQ0ADXlBt1X5U23aOc9ddanZIZcLDVUN8epnjbusZrr6D98S
SkptTrrSlxnjwBAnkJwdyWKO/dGzO/ehf1W7yAoi8bRat8kRL6WU1AwsQqSwtXIX
MLkowiMV+s7vKuoAeM+zkyjf+FHg1ns6ZfX13Muvta2IIiNWtqLPYCFtLYaSNV5f
Jf9Nq2Xn/g5s2YdxxOjmU+a59O4FtWIAum6lZK7pANGFhROIJiuNLSsOEfJtE2AW
KwUnb/B96XnVgu5y2RSztp+xZ5vrVhOjftfyq1TU8UIP3xz7btrqsCKWhO3EwKWl
h3pRt6sYtHxNP9AE0Ma9d8IYO6UEdSi8zoKNJ08EGM+6plUXaD9X4uUuvzonxT+v
TXmO3cGYbB9LQHnT++0WYs6lPnDfNeQuXG7W20QfQR+WsRzgVBQ8ew/IgPD3R4Fv
LCAYaKM93LvJHvgd2hGmUWcF0DrmrjtuouaqEd5UCjP5LSylsLFyJzv681BJdWbo
L+f/i/ORm1jhqDbp7r+Zu4FXGLf7Jm2YASwVmX7Sd08XfGYqMic2jzTYoHYLG+lm
ZCpywYFqAh9e2xgWTooaODJYs9CUsWFDYCO34NVU2FDOb2O1K8HzkXM+j/Y5Jbzt
Yy6lonSTcykE1/Iy3acJ0V1p9CVf6gbz+YvX1VUzA2y4uwMXv83DTxMIIUh/BIt2
JvMq2hFps4/IuV8YrHgSmVDbjTdLYHjkkWkr5pLcxH++6rPVUrUOS5Yy6bLsboA7
DKvUpEqXW9LGdwbQjwVnxm1PXegLyK8DIAanCRBvggMmwpJ/tXjFfLsXpuIzlh88
rPYH6CyYmCRS4pQVAFPJUA1AjhvCz5e1aOc/GGp6MqbuSu99hvnds9x183wHNHi3
LPsZv2RWV7XXdl3MGyqDuf57KRR08a0JYq8KemmUufoC7XT7ifHcDCexJBkMg8ot
vqFesaWOoYANzmk3KcBARyrSByQAGlUCbHGvy2aVIqWLSwenWHXy1OBBE1+3ZUJ5
SdddfOGuNRSw39NOdshyTU9ZUwQh1HGvWq6M45XMHR1juGxpaqMiEeT6H/SS7qqw
fRpBEdxYgJ+rceFinB5qiQWK+J6SzkE1PL5XhiQ+z8XzdI/UQeh8op0lPsVzhWqk
dw6EqCMwMusMgEARahuB47ni/zMUI8I/9tna8dOkTf4Mgow+IZjB+STZMyzAcn7+
rLMcPwt9iNZCM6BpfLwGPOO5cIBmOwvoaq8m0MCfmz06YCC/bDNwqObU4prrubu9
QZcsq9Oa6wt6QzGP/GlbVfqaKFu7QbdEeHYsuF51U7Re65eiozwVwAAXlGQ/05Bi
K9Ge/5/OjXE10BTZbyCecP8V0nv4Z+cvLBTxNNryqi9XfhlhToXdsmi7YA+wURZm
sSI+5fmP3Wekw455i81hf+aJtcLl0v8plqJ+CwudZIxNHZjv95qkhzELyf+9l2Dl
ufX42wac0qstc/RYGu1KT6y8gf91liFhK/nnRJs6zfZ+/y7CzZ86i0Gug0XfqjWM
w0l8v4WcYiqGRwxmUM2+9HVyEx/8Fk/6sKi2sDyORT8WfkxX81csDpxqilzWsEeQ
ebSuquJZ0j/qDbOsHDgE2rFlb1YJqg/6/2txAncuK6F4jPKFRr8CSs9HKliFCCJc
lWqM0waKhsG7oxF0Vs2sA4Y36BfA5iVL72hpmdFPMQBO6OdBhHQjfJDkFSiyo8uy
L02e8gXBaV7HVWVbX6ppsuij9nmBvthqRTFNkMpz7EUlqCkr8WNkN6bx41lhYWFf
IVBOzKuWmW35v57EhB2ovRofQJx5UE4AQCFu8yy7dced0VN5ICSItD9wiaFGAlZK
D1FEWF4dXbKtfpsp/vyyVQG5+4O6AW9702djeeoXvm14UBCVuK+inyB8JP2CrEco
jjgzTVnEYaze7VzyqPf/vPf1buhRxj1NTfyytHmKJ/xnWp7CKLuJB1RxjD9P71UT
FkvGbPExO/9AVhIskkY6bHjAxUmU45NOw6TjzejPBxOct3mlfFoQuuz74a2gvOtO
MOla2wNOHXvkNvgGdMozGQsw08w49Omg4+LfE3XFSEipLKddTvBdsoujAggX+d0F
bEJNRgyFAkcipuKVLx35uQdL+qLRlAvw5PxZm0hKMk481BIaCLvURgQfLDnO4qGp
XlIsACvNuzjGvrCtqOAg+6CW2LiXh8IyOU9oQnKTCWBkSyUGy4X3xdyT7xC9J7O4
isGiDW7ZECgsmBCuIQCzgUwbMoXQa7S+qugigrIGYFsMIro+bRuiq+UROAGijdRp
jhd435YASjQHfHOXiC7Z14pdTqeFoWmbgRmCUkAmibtDLXy7iosd4F4BqiebgDjJ
rjocYZ2w+zfG2tXm8ycl95aY2UzYHzcGW8BXC3dmY7GTp5wxqhd7FmQ/j1ZVGtMh
r/c7rFq6agPzUBO3H71nk0JpKI4cP6STENtxnmdmkzN7R0LtwfwtHDESCMc/IiUd
xyRZQ3dmGLBqthP4rJCMwf1+BL4V/xEYjT/xnPfMQC/D4jSeBuhy63uNzdBsLpYP
8ixEJbPPStPwJIvQ2NrHLfyJn5mND8wzGyvIiOjUCNQN3YbrBk5PyxaHCFwQm8sU
9tTp23PYsRmDgwXe/sTQPuD3el39BeqTws72tWq+EiZMptNfbx9oVvbcY6VBLw5c
NNv6iGI4wQsNXJ/qvR8QzZ3E95LN6XBG8XggZMbxINJZWZQhJxxSbrb0ukN3PXtn
NB+YfEIWLgSKjgi+Rv9HGDP1q7ae/KfB/IApBz4BnXsE8ls4cFMoBfmXsjBafjyu
mL8CAWSDruJ4SUsuuacY7qmfmMp8GvVnt/BYj4LmNrTmUOv5OYben+zcNj3VzmyP
40wWEOGZ2/R5vsR3xUtq+wVXQVTqv1CP0qq8ei6RwSP+b58Qs3WhSTNj0wQa2UOQ
Q++AzMX3WpRSflSBIzIvSjSfxgDP/rPFxSh4ZG26MBUSAv3T/2Bx94FL9rXHfOoW
D2C20V4EVVdR9n9+NPSJDr5OyMkFqLJct9rNAGqLfqbmFWmXbzdof9LHVDJzVnPM
WTOr5+aCDdswcdTDBXOhKIgsQN/4YFQkm0WyH6urYi+w7zOt8Z1bskHGMCQk8LF5
HHmZzFfIvszfULEZyzJe58/OM1u6oo7FhqV20Mmf7yGrAuF9I+/bnvSwci+PYGTB
N1e0QU5lolAE0TWOTDi1DYcMO/dG8zpI6Fl/L54683jQMtSA2Lib7sgoyHmvi56M
1MIpBonhimms519KAlNYQdBT9N1mw9rlB9KNDRkhdls3UA1hVu8g02wGo2V+ZX0B
m3g5TNX9K2VfH3sBuUCldy84wep7b0CpvOlqW6HbTPl8Vxwpc5Qjlor9LKZJ27Tj
T7+vTr0Kx/LlH/CsMnDW9eB7euwMhUJxIjiUxUsfRzDlf+rtgpuaTi9QZBoH+cqr
9PooXNHG1Zzf+LV90MlZg50KWDqIvHWqTDmBg+fqE+ajskERRWQchq5TAU4fuXo1
UtqrMkeSUE/49gicCVnwpyKcbRNxPatWRyNOSN1SSNbpyiXtuXr3TZ0+A3mLQSmo
kheT3/xEqEI/gnvLyaELAZCVWoJZYo12S/Af1hbABn4o3c/Xk0uzya/n4/YLHSXt
wzPLM9tmoGW+iko8vJAOIZpY762pXImG33DbkRv0eJWKg+PgryUdZ6ZtsswO+YU3
BI10byBfad4ghKnFvcqmv9El15+3FnU9AQWTiH3FAti5eMOkefWlNwVPEeRXZcYI
72DWDelhfp/vvGMRDw7Ld6wweEte2FgAg++w/2Kui2Qf8M/ybbUQqeby2BtCUTqe
BB2cwDdFl1uTLH4eB9t2oHcpyo+sNV/PmnAb/ZF0va4L1wpmg5YRFfLmerAZZtU7
48GPBMXuHiFtStMlqYipWYqWUBjstm6/lD4Z3jU3Ay/VvtKU7uvlgSfHALcQ8fGk
iEciYig0cRvsZEamIyUNR+KR3Wifgz2PaiYmqo3BrkJDD1qTMhovNAfrfCRG00VO
iS2KWNZK0v51S2A7zJhIMRBAeGdZYvNRufPERZnBMkWMxSmKz7BuaLaTP+QGc9lx
XdBgTbhSih111J0QRNTu6PsSsZV8rzc32zMvnCJRcyfDbm+bXVEg0wHCHlVq81Gr
jRvUZFp/Bcvt9PL5g+FU/AVYZbyePOgp6fb+S45qPkWjIjVVWWEgT6ePMozb6NQb
6uz8O6XkdJu2gKtnBCFA2UtFvS88SkodcWX78zLrb5WpSaAgVh8xp5VWnMYCmI6h
UryY1KriaaiYTQ+vwPsFi4fzuIwDuqXbGIfn8v2dEZlxzW92hYP97Vh9Wpo9atT2
S4YHt7D1iJcmsJSx/RlCFctalIhJgBYTwPHN9GSWTFiXJ6lKKMXBBx3w7S52VFdu
Vvzv62h3iVUEAz2fVkC6Ui4pl7xGhzrhhh97kG2EeSc+oJQF0/w98G6dmxzwk3VB
gCASA8zOCVf1qX01P8qwShZPKDO2t28dhGnQMf/KqJ9Fo30iWtXNeyOoumzbCWm9
yCeb0icmAQe4IGQmZj+P0bwE83U4Fv5f48V3wF7eLtVTCywKxfPPhmDy2hPkzrFb
ZLUjM6e8J4hdA4UFr/bfqhk7RQ3gB96L8/IGB+C4bRMJ9b1Gs6Po6jrGSl6dDYVa
nAvURXUvJ7hkdvCKRcMr4Zvx6sSE9rCpsDdI/Yoa2eJ4VXgUosnMyAEQqTDe7BgA
BZCsmKsIT/83rV3/YgNuffSrUuJHYGxbj5c3vc29JfuPBxrxBIc53vclQ+t5jrRo
g6CfepSCuWeZl4rAwJDSdVPsQghUFXOjP/nCxx0GoR9t6kaZ5Wc5yx34L4VWINzM
jqnEwKOAO51fuMzhcbaEeKfEBXE2rbLwF0y2/FUGMOgQhDUKdiNO2O7aPfFgdWp8
4pjt13QEuoj5jVVHQJh2Ta+H3CT9rwfLds2yLMcI90OIbPJDMx39OGjYytOcjOdZ
TbNYH4waF7bC9mdnBxG+6TOLZ2ERiSrSZBz8S5p9pFaB99p50HMKnwK/lLwl+2f3
3wRGTtfQoUxPGL8r/zHyLa1L8C2Qpp7WMogBGV7VGOLjYC3cMp2D9lUlOHdBx8z8
CZRDbwJhENnrKEzZ+B0VVntng8458FlBDZ/UKYB9Otlu8DGSfauOxi8FSPcZ2fT1
SCytJyyyOFP1qx/+8fXdh6UXNyy12bmfa1KSL/2wPtDIDPRszhyTZThwh9YOcQEz
+7dVegt93wMFLwezj4ASbEntoIiEiDWPdcElT7KWkAfAf7DTM5tMV9znfR96yql1
tAHxku8MXZ2m85O+9k5UH6gOx6WwOzec8DlHIzd/17+nCFf4+/CTmcPJQcusz+jM
Y+6Vdkcxy3C34UA0a1vCAb+RAOVuZfOX185Uy5U0TparoDFc/sdRU5sFI91uA2lr
V1RdgxmOvSizfO5vof1QaGqdGudOhCH+x/saungPTsUgnEhBARJ30oL+QE/gCONt
XBZ0bbP7ZKnuWglkv7UIsytLhDoO8Z32/kl/eAUJojTMafTcpS9FQzQAv+JxjuTE
iFfHbVVnE5QYR8Yac8SAFxrWOdcr0Wgiza6FQn7f4NMg7XLGkxAGeAgm0UT8cqaP
8CnQZWMKXXz7rHmBfIriOI1+p6yjOp4Sfr//3owvYaGUx/HrmYkQRhplBXKJnsBT
qalvwUMQAmv4x4M7OkWKbPL0N9+7kTxbFDeozji78n1EBCxLjUvYcSL2QFzcO5Oa
qwFY8k+9AxKAk+4AwIn8ZMe3/k2mvBccf7r5zrrYbgfXP4UQR8B/Le4sQjuk4xk2
GONpCajylPCDbGiSDgFOw81LBnDJ7SyQW79S4W0HZq9eaawgcKMizVynyx7RN3JA
6kjCTd/lV08stP/ymvPRP9YX4/70XjV6Zy/dxw71R5VqbNlflS+g02aalFP0sJd3
Yck8KFtVrLx2vgE1VwP+HioZJ84vG8Q4i0sjzjm8ohSNyCdHWomIWHPjPqol7Pp2
SCeGY0QXT5h19ud1z4l7aS4vvwXgkB8Nf4rRyEz7CBxZjR7Ag30d5hl/mGN8s+/P
ZCYZD+r10QBgcKeKW90z2dKjmHNqMsbWaWczhYKqJBfGVXfZBxO14xG89PTlCCG7
WeE8yUVOcoV3CSIu3pZxY3o5rabN3Mwxde0Wh8fXFh9OARRfBnzsMQDkAO5bPgq6
VINXrCu7zBaJBON0iZVK5m+JLYQ6WUE3VUXHpmEBLXWvWv7ZBjATcYOcyJ2wxE1t
Mn0KRi5o8Pa6GECgENptpD6l7S1cpuSHtvTfb70Ludo5UAp3zST+E/979xLASr1Z
974vmjYaXDWKzZOxH78fcJ7D5aU67j6Z4VE6IkWXGAlBHrCPAZPnVHrmI73gpITs
tK3hJ4zgIGtD5Vd33EPYtaJo335yP1dGm1tcgbUYeZbr3K2GAUxVTW0wXAo4CwF3
fnmMXXnOUSNEgnWQRb5QJIAlNtmuIZBLMR2hvukL9aLBn3h99TpBeMt1ONon41e4
+E8vsZTY0dpFuyhN1/zwSNmsEo+Cxpu/eDRnZfvmHh5Cauvwlao6GyD9/YWbxzYk
vQu7zHnTuzovFY4cpNekP9Twc8La8blS4hXeaV8vhHfJtls9wc/gNdm6I99cQ59q
oVR1Ckn80isQSYuEECIhoOb5ZwCIDu7rdj/be2pQriuh3tm3ioj+ZPRgt2TByinY
WsWPo4CCQKUt/ajDiL/6CIVXWhXlhkFFYB3198a57Z8pZnBuPICsyw4zuApUoVpO
Pwqm8GRmiTKexOt4t0sNk8N1Ww5kDacPw0CKDvnaFKkbLOJG7XJfBbFVNydCqnKv
7QlJjyNVLsxo4VgndqJDavJfE6BqIt4Vv339WMKduKsJzevnh5Oy/Cv+I9V/gXGL
q9BIdxd1oL3s0xV1A1x8uzDXUk7dLfEjkYYmfIw9eIJviu9ghabe32OebLIllmDT
ssDEHlFst94qchXkyU+HbKCdjTmz3HnFPFOW7Qc3eJHfd94u8fsnG+Tp8UNGcITI
dZXOhLZWDi2n2dt3dSyNENENPWOfwRBphOAsJ7O/FmYm3IlnubVcKg2LS58/LOFQ
jWhj2ClkuK720xf5L3b9223wrobFGX33vKYHy/JL7aJUNXjPz7asyVrPLs43SWMp
npgPhjU+cCiRjyr/7FM8d1Mzrq2Z4pLYTebZI58LrqArKJnP2SYh2pvr9JT0ZoGE
MQnJbNemsFMONFZLb7Wjgcwgnw8mVc6vbykHXA5hCLSo0/ToVErIQXMYDdLOLKu/
7Szs6oQCVsT4fPD5g8S2ABfKJ2UWDKYSCiQtAeMt+E1JAypMK8NeFq2S1HKEgoxt
D1GuIZFcOg7HNScwfE/AkDcBWOBhSix9CX8XW7utbxHN+eBLiP2eCPph7clvGzJN
idrkmLg/Zz9SeIFbFXn+hGU4rDq02MZdhj6w0p+eRDg0XLquNBCk7b/UnxQ9X4iU
zbxSF1S8GzEsZDdadBSi8cLtk14fWyt2Jq18CcoKfo5xkAX00COaH9+ZE+sY4eGV
ZEf2wJPdz67SDcO0uGbTLwRCTsFMR0fE5K6TdhP8dc8HH5GkCjKxOWVgFu6kF8oj
EBZKV0PB19zpgRDoAP18iwthHl9r+0B2qDVmmwTzmhTFTrsr8au0u6pGtRzVgFGw
oDbQY5gtPGvIOeaBYL+pOBGbxvubgvKC4Lbx9Pt2MOeCC0DAQOVTAqerZUyaD2Y4
9jxvADz5Ots5ymtq19Mcaoc4GiHplexNmV/ctanxV/LYixjX2iccl0XUusxuXVh/
9OkeemhCqFC10KHfpm/gtxAW8Kf+b12qP0OzY8h7G1VH9FqHwVyUTrSCI6d8jAaK
Luh9LwpetVVl6DyrhosGjCChuOAfJ1RYt1g35rAPD/3nAK0OZDh8/SlyYvDZE1AQ
I4fPJD5gprUy5upmoJrKRkfBLkUUXEB/kVTvWbL9Q5vv9p3uJLv/NqPfkuwJ1Nzw
pspUNLqAQ7KODdNaqP+e6J/HSOERfMyKxuev0suMhWw8Htn4fXRbf340veJ6sXHA
vZ+ysw27Y+vQcJo75sQG+d9sLK2fpd60pMZM7K4cGR4bI211wt8xYWF1SOMdVvh9
oxFXA8evc5pB+NiTIfc9Cm0c3E0QTgod5Z3sSG2D33Sn+MdQk75kXaE6vSo1z35g
0grLhRf1m87F60Xpe3RPlNNJglKRqaCdY+zRH+QuBWPirddjefW3zzLG0ILyoTGQ
vnZP9N4beRFyte6LQv+1ptjhCyV/RCKRubT9F/QApWv8RwpHpV0j/L2pCG8qtDAU
OXB3VBRHGjw7HjL86T1qKPXhzQ/ZfsxaI890LtrXaeXpiyDYNRFqa4fQXE8mvC8B
wKku2QAjZ+bD9ovAmck1IjpKXVz7XY3o8f9BoY0Ovqzrp+VN0iu23uUc7TQMEYNY
SfwCRwClixvkMzfAJzgvEMvbmXkKJUJj/PP0WeiFkS94YR/uaa3aw3vdVM4biOqU
damwtGS+2R2OCTO6zDfb4X9th/31Tamu4s1Mya22fsZ/ph/C2KLxd/7DWXxKbhRA
bRsQzBtb5SZOfjM4twcnCo6/cb1fhJKzJ0QCpyiTsm3i8i9H2tPWOE/zAI84TLDI
pXylFA9EC5g4aOZ1YD31ep/AKW4GW7vfDLPOxBEb07u5fSvo4kWMSr/c9xDl/uP8
gmVnzHB9O7dkniZS6SzCdWMp96u3+3mxpnfNv1JjQXBJJdmbsvuFLyqyt4+IL5Oq
uFqlYTK0CfcxJWYWiDEm1YKpVkohKPL0UuHpdYZPXAdJHHGDIJ/3xJXY5MiG1O+t
iWchwkvLh0AENrSi6e5f4Nrql7Hpe95KXf0yjK0Qu7i0UVI4Dnnx6RQVl3e0sdMU
/4udZ1HTr14dl/xI4wj7kjfs/65SmacFlTDfLkLaRcz4XrhKEnAY+p3nIix6jsfY
pvKdPjpj7QaeZTT7lSWzEzda8gl0UIAgMar+4urfmA4GIYLO5O0yunomdPkPjjRH
X8r6fpmoFpvmKvVihgJsdeWiI6jOZrLAfzjK4WCBYNY2gq4R6xwXewika0Q0zh59
uHaBH/ZuC6c+WrtSOWgYTnySK+Am/r8fVXCLCY4yfxDgqst5F3ymFEjhdtA38coo
HkQuq9SAVI5lp4dEhg9WUMjoM24sfsoYuWNknp9M1h1AlaiEcI3aewe5sFmrRVLC
FS4d7QU8lAfshtzxYf/hdaVN1P3H8ALeit6UR7PUG7VVY4NYrBOM0aYQRbO6BYAK
GtcwBN+JBvPA5Kzen+qWRm5XecLZnrljybekv9MahsZ0vWEwlNAtBzTCX4QgmbNC
WbW5i9stZmgRvjaiR95jvWzpHgQYN/lAW6AHQUJ6rU5Bs2rcLLeRXX6rjwyyxNlX
ecE/AovWkMWkQ9WUHYt1ThdqHhE+yId5yVQF24qcJ9Lx4F67tLOS3eAGblycKZXG
19ElPtPqBX3zGAYd6tMJYkBPDD/wfxU1dYfeGxU/Gs0FAxz9w0QSHQ79UGby+ZrA
Gp64Oj+oiNwDlUQhmTNuWVls8QK1y1O7gNmmB3nNwWqcveFkPLnelbzf2Ip88Q5T
bANP7jKWwKoG2YK5R1HVcbslnnqU4GPHk+p5eYcqCphONN4M2khRa7UuCeakjRa8
TfJ5aHP3DzObQBWHGwtEamgmYN/V0/VfwX6n1BPe4VGfOsaauMo0pRNXIaHL6iLr
KbUWo+8JqP2oBPuLMHjmfMe24cdIxFW7U+gp/zCpHgGkDzB9UWjAHceckJBb3375
dZH2owyfcyjcrdU57uoLpR4N48XpbfRPFtBd9hJshn6RjmsMiwD1h/GrZV+D98v2
xR7QeyVeHxGRfsgGyL18orz/wWbwIa+cbYPDHd9JP52Fy1zISdaxHwnuVGtQq7PP
uMXsdr15cPa/zXvB5oufCTRhs9yl32tGcozmRtVVmmPFUHpZUoLYBXI/w+H4jy6c
AHUJXEBS4bTWJdalRbRQfO1PLVXc/6M9CS/m6nzQoo44FoCHX7QGIPprpPr0smTd
RkpCEYxiorffOYbLqx0ZcNcLGMQCNCX8SkYWTM39Q3msH6t5k1BVNtKF0aQLdEjf
K/FONyy9Bn8hxyZwpHtZRBRQ0kVn2SWZG+RZEN43BFVo+lp6tl96Seu+B1ZlpLw6
5qGcfrz27E8rJLVjPvGhaI2qoKYHZt9mkb2JGbR5axnAfKCXOoDbJqa7zvH6b57y
sCULFN43Y65TbmRtUEBh51tbj/QQxuxglKro8hL5DbY0BwJJHGY9kL17TOD5INOp
suuBxmTo5kS5DqU3HlapWYtzCTYYc7RKuDHLW/c1Ue51KEVkMparDY/ZTOEjNSVb
i9bisf5H7Dlfvymm88saCCHD3nu+MBVeCAPIA1vvIGjM8XhsrOmR7WvmtXa2ambJ
n2tN2MHq580o5jGMJEjnZUE1zK7VRn6mPntMcx0BlEv4ppoe0DNWz5g8FTWhCkYj
q/LZbr2YlmJLc7Tw1d7cWT9RlMI9nR3jLRU+re3FM2RwLHiC7pxanw7itLentnVt
zlFpq+w+ovKO5iKb6KlPmSOXfu4cd3rjNKqfWhAZloU+EMpUYkUQszyH4kRlGAdg
523N5yNqxU29Ob4PvuAIkTh7WpcA8m07Oh/AWaq8RPbTS6b0dMzHrAK78wz4zV8e
Y6pWcrFC+leZNBXQpbVorBu+d1fdRtRg7n1fGHa9A/v4aC8F1nZJP8Nfz5I/jZ3x
dpyA4eOFa9R+Xp2NBWAcnjy+Yz7SuYs4InFbts668++LMd6nfZKGT6NqNmAXH3J7
JAAcZvT9TGYDZwODC1fNtXgZrRe+1y+kwGetVNW/TML8b3wR1VDKeCwe8vBlNGIU
lovs1hWMvcaBhVZSBIstQW78aX/FsWjgNIMOa/sVEzkJ1fDTuEwTT6cehkMfts+F
F5BSFefDH5WsVIg2wxWwJ72ENoj0iewA52j2xRxMQOxe0iS5DXVCFd1WEmi0Erkt
xg2iTjysH+vlqJDImhiObDjxazubhE9qcKDfWTQphtr1iB4tma/AQY14nmncxF1m
EqdR5Lpmf7Gju9POgAfJB7nb1Uem3XUDtg56RweVX6s3oeyQpV4+Gww6tQx3KkqB
rIdIzUIybsKJTCIekBoY0ZF+rB4TEjmBL9XLdHZvEIexaTWWyJwFNOxSXL2vgI/u
+7bWuEaCMyXjXzGY6YH5i9weLBiQd3tI0M5yYIrPjA9fleooSLR580REHlJnYIbF
2X6XbsfVE72sn2GQeu7pIsi6qbVFrOCYIWj66sS5ixwW2qzE3kg6QXN91pyrefx+
Rju3W+MWf3npg9F7Ffv5b2DVQ5IyV/VA3NHarf83yK2SmFj3Cll6CzCjoOFL4bGc
dG/LJwrAG1F/vFeWYuGjrwyMPErsLXy39kUNkQiqwoc1d7r5q56LT6js15IUVQNP
Hzu5YU6W0MgPxMcmHn7hEO+NAiSfHn961nspTfZ7EexTOWdCY+Nu0roEu6YeCG0Z
28POo2Sf/wrHrIJFsLDs12mGvAo2RHCOEix2ACl5ld9SImt5JIxsVLixMfUWR8QB
xQBtEWD+3mW3sRL3WlulVG4b1ENvBtbgo60B4+z1AXkGnIHn2fvHYovzZULEy4u9
DMPiaNke0TX3qN6Pd86+rdmd/lEmPDUh+ZeeoytTiRYHBLJ0v9vjnYfpzSzerwDu
5JrA6RWWT9GDKSZwRyMNFiwodQcehmZ0da88onLtGndiPHhQM7ccz4Fn22c5OOqh
46hxwuoyRhUX3FAzthY7OKIiGmcX+3ZLQH7R3DqIZgLfNbfLT/7zHnzr7mZC1VYD
Mbyn8CUwMBuhxTIR3iaTgZFrB8vV1J1NyGl2z6cew7umhqSxZ+7Xv9P2UgAiRI11
FXLE99dBd0nU1hAuhkVN5ujlKCO7OObJS6lVPNf1YIWRJfDdnIM4ws2v57X0cpFd
9xK0xcsF0xxSuhoTCzivUQTg4SLixr8LDCmF0cjoVL5/3f1Bj0qYkY5+t4Y3Sshb
8x6lKzuWzV2NhVYX3TJq79UBEv8q2u2E17yNLmfnePuRwRGMZLcqAl/EVw6KhnCz
tI6aist8N8qkIxZjGFU9pVstdF/01PMWY0GuGPHbt+p7dzWSI6ufmPuQ2Qc8jz55
8kOkHyQ5TlC1VYlHjDeLM8xtfCZB1KaYnE1G8U/PpFaGwej1iCxYlVB5MHbfseF0
baIvO++rmbRqJHjVx9tdEtbHhu+26zlUbEn8eAuVRUK0M2eG403e1zkEvOhbd3fP
CBgSraM6c49dKZUt1MAobU4rClbHYut5TPr/0aNY5nNegZEbN186rB9Fm/oVYpL9
HChWL/sJGlA5hwr4zAUZmPacqr1eokxROYte9k35WzCKQs3jDK/+pMCN9SLADYl9
m1XQmaaiJ8/adZw7VVbhrG9o3HUUI5qk/9hT6c1YdzwgHM/V7LW7lmjXMuBz1+CE
aWC+dactDQ47DcM3rexDwcDcINFvesedmg7ZCxtr3+Aelav764czO0cA9AQBJj2e
zbw1J39rR4cNvzV8OGcACo7Xjl5PG3UyPE6P33eGS8Ji357YKCmHbLmW1z8Of1VQ
d0/jkL+OjtjBVJm3YJgrTLGFbmjmEQAkp2OgPZq/sjZR8eytVSF/6IPFwTj94tHI
N697ErhQI2OlJA9CFbkMMVlJtMBS2Qj5KGe6ATDEMfDYDmWWFH0+5VORgJx6HUBW
QGWA581OwOIU9EkAKRD7WFOZu2VdTf/Npahql/wPbt+2ey5wan6YYIOWxR66/4Dd
2odVX8Q17q/h68rL9r+zqeMpkJ4Chtcq7oTo2XI0/qeB7DOrB6mINtryN3D22Hff
BgWC3dobwZ9govoM8ghDrmjL79s3UsvLRaBW2afHI8F4a6o94l07IEzTbNFI5IHP
wVSVAbzKg99bDqA9UOg1UgRMgNdiFU5d+3VsrQx4NxvO0SBipS4l4lTY67H7GzR6
mDJnDwZjylXV3GM0ifZbihz3gbx39KcUaYjDD//rbf9XboRqmsm1GpW9Rf4PUHOO
kJxJ87raQNnpsf4mhLMxeFWOOse/1Ezqv1l8ZkF7jnFM0XtBcx/j+QaC+3sldes6
LsinUmHbPw2p5evMv4Be7cULHWsyuzoteZ9Q1W1Vu1JJSHr4kDnHzf0UWWKiZLl3
7kCO+CDioqJa0TnB1lL95YhGQSWUkqO6sHeKmXSvYKuCo4kr5htqkJgAD7MnU5TL
FOyjAxNd6Bvkyrb1tS8ncjwws0Jt2nedNK+YGWUn/E0pYI67g0dqEVC09zuw6n3A
3KkzXBsH6qR8tkN94cVHPd5vYDmIasg8Od5L2s1K+qBVZ652zoPUHgOpvFaBWd02
vFLEtHFlrK4Iyy7zEm1gWhKJ7rv4ypJ0AmySKAy6VsdEQNUrxCIxXpehrbZoVZk+
pgYpCOc5ST6OEpIA0rUE0Yx8qOzM90IOl+1N8sQUq+VkZGrnkceutRV3HmzSe7xD
NbSwNY8GTCjEUuZP1G7QN/1k7XNeqJiVpbcmxbm5vI8LqFFHaZMI45LsekzTXmZq
4CzJ5F+gpD5OnJP7lhMRfphkk0BkInDUIXqF0ZqXUCq4BOuZugxpIXyD2TZmvEmU
bUmmgpgeSDe6TtCpmEISeliIYR6SvUMYRS8cV+uSEP/P+GbYuVALG4Dju62S9ixd
9k2Uq3JFKBstwEo3W0GdmmGuJPda5zb2G9eMCG6ELvnijP14utMOB3JRjNRRyyuQ
VhcEFzkTsLE2mfXeKjUIMDg6W8/wq+KlnbY6c2BG9jb/icP0opesVEjWWGsRixlp
Yta+MeSZp89Mp16t4DdIsDYy1wUNNbsP7kS4zYZmDZBIvYBVtJdRhsIksZSSRBEv
DjhYtFRUVOk3iZkifQNv/0Qq55XTkYazSDsIyzPko6gT43CEKvUVnJxZmOB2oeoE
rov6+DSdgBXS0i1dVHEjdl/F5Zj61cgjrkOXNa33fssLxPxhmOJMGqVEXVmbNf7N
9XjDM/8ejVjj5Epzjugzc8ZjQzPDDXdbl05a47Mfn7dySCrrUWiLu9LDzui8WufK
2rwGM15QnE/IAFRm/OxETpK0/OfhSiHkYW15aKdOpY34tYCNkFBk7u6CYj9QopBP
EyvZ+krI5ov3yS4NPcOyerxfqr/0gmSYXTFzUCfSuKw8fPApShqn2Q0gOdtzoqE8
jn0obT6oGdXH6/R9fllnJU9Yao5UrvIraO9rIpGk4j9WqhBgoxAY8qkkdg/AqIHa
AfVxLV8sC7dsJbxQF+S4zVpI6NzEnOTuVTunl1I1DXmNSXsX4WLTf5N/oJWpPEKs
wFXIf2Re/PfkbIE+hmsgv/t6cX1dJIhObtv3dWr0cGxjhipV2gXCSu/XBKXzYkP4
rQdLnL2HkL01ZCypNj3TS9a2/lYcI8nft0sOtl41/4ihwsFHttBr6oKVBs9SREJN
oZwXaM60xoAKoZAtwFH8Dc43PW7iNI/x3y0cSAVu5v3Yq50dHYMUptAXcqFyE6JO
J2G0jq7fXI7BJOxrJtUX+IuApBoutgeZbNMtbM/5zPfCqd7TkPikj7npeRpv7ZnR
tYdrUJSYa9zck0aU0DRjbI3Q9epAFV12MmU4aHbOTkT/PhiixjCwwywoAGFPMmpq
WMJ94Pcr2qpeLtNU2PVhHx9BFQQXI1Ap48WKXCN/lZLxIgTaZqX40/Q8K3Qckc6q
Also67ttC8jxkNTPOHW3n11DlbsHW9WO8ZItNDA0CsmMMr9yxQkrlWrh7akGtviX
UOsuBcOeR7kvWcLOsDhG5pMkIlHuM7tI9LssqA3UVTfyO8f4IXNkYFLb/y2yVAWa
h5AnU8EuNkPSvixjESE9k/lTJOeSOI5Js4y3oKnXaCXXK5iTtxIOkey4R1yxl+3s
Av+PqpSER7OwOIwc73b+8TA9VCmr2Xn/PvGdGoU/AZebmk8D4Xy1SMpW1V4bFTPp
enLyjvQyAZ9o/hpgJvji/pNs9aJObK/zkHAPA581o2V3SIFaw1JeWm4grsdf7B6d
Rg/VABr1fMP5Wb87j8yzhE9bboI7kEqHu86DgormBdmnF7jGsFs04hBk60va9qFg
ENQ8HEleVtbN74jzLLFf6QqxBX5tN/rZUrHylINVlZhLpuddOWAqaQFiMOkeq5e3
Vfmy+Q34jxZ/4tYVD2UWTPnJ9HSy8nDX6KdSSRyHlGMKzN+ey969gvk5eDELwG+l
8JRZSO5F+oeWYfq6pM3U7ozcPKN+rTeDMKCmA6Q3xZTv+nG6jQVLtJgs8l6TOHaN
6m78EQd01qID45tOPsWkK2Llr/bglXeTbPk2xIKYcFyM6mrZSElm9hFo5KPN6Yoo
a1GYp+eY0DYjRTTmRxuWq6cFPkSP6FkWjNvkA/62wvUm16YTEr+HfyZhuu6C+bv/
XiEmY8tj51EO4GDeLJxWpsywOxy2nLnk4AU6rMM9ydJ109Vby6G0aK9bXNa0vbpt
5bkNHWXtxfkj3+/Ot91zEzzW8SzfrQq+7MarzjbFl9leu9n5pVD4BIcEtOgRDTrH
VrkCYk9wma7XJBR5h8/T2xkE05Lg47MtcK4IVO7eUxaJsOc0yktWxGuBXfEEAhTl
JCREwdtfbajXZtmDXCmTr4pyg1KlqUDtHcRx3yuVUoHVV4e5/E+nkwEM4A4trnGJ
`pragma protect end_protected
