// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b5dbQOP6x+Gm8gRWhxrQpbL7bcWvDpadko4WRyCcKA5LYo/YaGjjYMjLWbQy28og
injJp9PfIgJGBF8TkdWkzLukbsukrHPcuXTvZTQ+12kSijq2qjcFJDISGIKqKgfl
p5JwsTAPP9T6kxadVmcSaLDEFAI6aIXngEMGPXejqNk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17968)
u4npuH9NVQb0M07Udq8Hzpx3hclWFLKiJkcQH/nb1ccgrNBNN8Db5jGlUrhtDeIx
Exloks9OjDRDIuZZSkrk7Uz9tVVHICDYpvBfVlFDS/sjU6/s9jky581HnJSPjMrH
2RHa5poLBSPbXPpsz4zBmXormV9wi0BD1934t6pQcbH8JXnGWQ8MV8AuB4N4An5g
ebrs4atJg5nWZdxAu+bhBW2j8r9v9yiJg2zddpT11s/UseS+BKriHP8l3LHKqs65
n4crUviu8MV5dM6p4W1Hm4/TH1pU2sTmpxL0cueBaHUVwJed6x1cFbr1lH5y9RhU
4Lthv68BGNWgNYy56FmLpnlhQzzQ+hrVtUvmsEBE8scC/ev42ZzFvpST4Esa6aLw
XlrI8pT0usBSX9Vv25MOVrtRimpXhQBsKC8KlVlDlg/HWELpMqLcrfHHrJjzFVBe
TD0cGA5q0ws6nRr0r1a9mfq54NrShv6qKjB84AWn0BUsmLQkazPRx8laV/ocaBdy
dg87OybvTLagEoyUCCKtnnY9mE+v632AgC67hf9gf9xI5f5mZ70z+yNoVy76PSCb
XdFSUI/9hlvNt/GFdDAhhiwdaFOZgx2AQeMXdg5RjZYDqL/+iiJTxihOVTJ/gmvC
AjjO8qzDl2JfoVFmK/nVCefy2b6B2lL90ZsvC9QF4nZDDc/AHxlyTdFl9TYov5b6
Kb5gGrB4cObAN/v197Vx01jochF9OOkMRn6VbX6+qoN/wNAtvUCfMIx2qkul4VMG
FEgdA1qEoeHXnqEFoOdu8U8ETUBfa+QIJqA6LPA6aMruX80qtL/8dY9M6GjHlQFg
tnKC0y7dmTz3wZi94EEhqcrjLS+byrJW/jHpIJe8YZVgj1P1Ukb9u5wPGy3jKtf2
mm3j18Bx39GjlAQ3/5omniMyY2bHxDgoYQoLEK/t/QAXdFXVaE5Fu//NPST/ilep
UQPMDAQSCbbfyjOy1kwa84X5nrK70H+UHS0zJj2BReqKUeY7GU5KWWG93A2a1BEW
ujiEdk9rqucfqQkr/qgCkSqE6fkHcviBzD60hXr7egitcsGjc/mpClinl/tLFHXA
DGCKprPVrX5MsFnaTTKH/1Vy4eqaNrhk/wkdc0hmVmzzFyDBxj+bfT3LB85MaTjU
M1cMfZgt64P+En8cPk4D5YNhq2/bwiMLg5W5lOQ7a5Bd/+VqOEOaif0bVx1nZnuO
5hL7VtlHGzn7n0iXpf95jwiWOVVci7Upgp9Pidfa8Kp4SHGNnq7tdO6EOTBfK6Dj
SDIVVt+SC1v5dwMbLlxyjh/vCJDLbEPONMf7G+c+kC3bm267ziC/8HF5oVOzMc7X
FUhAuuX0/vXby1ahTYLgNl2whjdi5pI3oFIRzlov3LopLr2ri4ASCQFVL4f22SKP
Ggkqumo5rCLH3nj0Q3gn9f84gugAERPJUgNUx/tBQNhhLJvqXf1yjREGM28HBbKh
5T9SDeadKXW1eTTi+/F1/dRMtQGmTR3HLVA4CIJqevySg8qaT/fD4f6X8ksbYYZ6
QmHiWlI5xBheknycHokmH1QpIuLk2EWoE54ikBZ0kxxzm2fDsXT3bkkB8/QvFcuE
YW7sCI0s3CXu+EUcchShYRWXV6rVQnPp9ZsKwO+PSUS3tLujIr8dMi3QMHVyQyFh
NQ60uHjd3lZievflxhlKnX4loqnzDbOw2LQpxondFkrecwG4fI5O7/9Foyk/xci5
VvtPsVtWcpEb0I39D59ekDLPe20scVL1myOKjpA5vP3bvKtGOlowClfPKbCHT+aw
A/TlMX4DtBV5OqeRMZO5CKUGFnd81I3HIPIGc1KLgpa1IenlivNdo75fUaK58Duc
djO8Yl6UYBeXWwQ2sWxGM2FUSyFO4blwXiruXQ158T+s2JnRhj0t1n/rIY1WHTSg
VPx8wvt89NGQyUY6LWGSZT/Hevy9OSuqGov1Biq6coOo9LhrxeFQrndOR/lhK8jC
7KZ7vcVWBD4wZecN6KBmdZenSSw+XNb3emGl+OWc8ztF/kwa748h6pGtzOzaR0ru
CGKK6fleeRhL0NXaSzzKgOtXAMdQilqjV5Tsghmtq0q9zZ+F56OHxIJs/E+D+Pqt
CxKf/FD0cwSeN7E/FOXGdonh88/tPgEZwtpNl5740zhxAEyTajq3t85Cja5h2Tu9
jGMyZYXGeNhMp9qzPhzRN/BPS3NyFHu8tjujG0/WhqrJhInkdZEgcfrJxh/I1h5Y
tMPyJ03egH793OiRSuGtRSPo/2FogWcCzZmBoTh9cH34haSFcw9TMlRBfBAy5IjE
/BMBeaPUi9xvqXPUgB5+OBsqtr9xTaZTyiVhuGAYb61JpxFInUcX8b4aKjtcrWjD
f0Kvtr9wN/TH/J29mWVdCE5CnfijphMhcjpnT24easPpmbAzsWUkE24GzUNrkz/w
va5U6t1/LkC6G9hpjKeSsrbpbzvXgRuUmQpEZPkdkUFt3Opr95wQ888KshQHsggR
CJEpwwgQm7jaNTFmlz+XcIutgTFBOffxT+znA508/vPnF9nAL23OGzO2awLQX2wn
h5pHhVM5Gf39cKTN2wcNmQU0/p1Bxh4wOTfE8eJk2ERuYj6r5/TRGkDwbvo6WkQb
r2dMHIWjDvqhx9RFeb/HJTLQpubNIll/xDBMl4LDGN/TnlcGvYFA/nrLa2PLbBHs
z2lWmOo1NDdw8V4HJFSimKvTYaJ2e2k+VL5AexsCYKhGF9rqu42gm9B35nbLgBAH
WDzhK5m8WiB8kff4IcEJoGKaQG9a+95LD7uydENmgPGC8At69mu8JtjbS0DXAHcv
5J+vFskWNKrZlYoDGxHM+MHSsbm/Xy+Whv9ustgSSBsoW5chMFOYVJjnmoCuZ5mh
bPRFpN0jjb0XaxyeJE91WEK9L8DrjOUmT5izpX3SIrN3ApP+LXQo3Z/Ym9GIWvGh
az97oW9UJoXN9FdGlb4xOm1JzaBQvwr9+KPn1rlhx5JHqW33oHi2IiNhXTLRvt27
XHgcnQvs95j0ITNbT0r1pxQ9k8xctDnCOL9u9s2zfp6Ni0cYMs73Blnq7CK0m+nJ
FXq2T6dkt9FdfiLWWAOKprM0wiQhn44HFUJ6KcHcPc0OJZc3Bwrs43Q+qJT2jXIj
hnsNEDrvb5ABipqddNEZKLPNseMRs2yJ+7O11BIH6ZhjZQ+NclwrRJiHZKRdtLn0
+6QHSlrjS1JVn0zs4hr8LY/UdIcbXB1ssUY9FMaGuVlSxGU86mZxQiLfAdP2ZQpY
84Y8FMqVF6lMpOXLZxBA+x0oYXmqCRkAgk9Xk+gg/Virpb4lps8I9mgrhLlKT5Ny
InJ97oSxS0Q+HLvksrKWGeY2xa6vLy9mBEXsJrxUzaqxJ3Tn1uhiE/N79y/amwGl
6cEir0EBs7zWs+omjXq5rXX1hSqF0BZkFVFeUpm/aupuGsm3xknv1hy9xqHKFNFh
MiE9uFpvRC3noA5BkXdxrp0UP9OfoTkJIEDiumM7jninaRmArxKwy8ewEeFaqnDq
qw8DBr8wQDQCCKj1KwRYhXj0nkpVxivSGMrjOEczC71vqrQ+4vIURgWrQKOegtzj
5hYPD3Az3iPevLNRggswjana5B/cghq8IEkUrtsdXrS1PnUpbSdmm0UYNIUlFlU5
C6n3C+qmvM8GZ5Ij33EtKZj2F/FfDCaUrqwF+VEjfoIVWrma8meEna/MaqgyrTMv
NHLPKzqPeYTTP9Tji1algMf3gqpHpsNbbBXD63dJVvdvrOv4hlYdh2mNTtdI2E84
/G/BKjAwyEtXqI/vLwTUtHXLS0VCIVmi8LEo8UFZvb1GjGzGiOavWv1Ra2ONHyld
xcV5CQVv++S/hYeI931I7Bthr/wB+kIFvfcm4H2mjok7Xfxb/7KmXkHa2fSrKZkA
e7ScJ8AWRD4WSKy++jQDbZdxktqdCMxUNS/LYQkC0A/4ZoSm6hy+0luKNnAA4Cxm
+9uqDq1Q65Sxvhw91IWPuuXFIhSgXYqhESQQ9qIHueHUeFvbAiLrFg6hszFWXlR3
C8RemOvn0v3IzZQn1LX3HXMJXMjwU5lftd8uQ0bb7tSY7bkeiG7lKIkVKcZS2kbd
eXhxEeD0rl9XbMagjsIaptuy3ukGvUuC8qikJRJAKnZSmAiZgWqa1z2hxEM2+78B
rnXbBSoK5uQvKnP6kiXPwU/gNNhDXUiymIcW9ejjiYXejhzAJ0GQwA2vqW2ADSu/
R5IPa11HyhoSTgd02jYkh9CuLwkrFPf/+MvtJAg0W1EHHZMlVqYDIWpqtS0ksmTO
NyHi7OtVO7sO5E+jdGVGxtfcg0NfDXjVxN4GVhSoOYRzAWCV4WYiBIr4QocoFS+v
D7NzeVrkrMfqqNGjDq0ah+zqhJ1vHWeO3X2sdoNyXrXvHxyjAavhZcbQgQlLlANa
jF80148dA9ukVe56IGvy+bOeFMCmDSN2+DgQriC0MvhuQ1aPzgv02PybDE+0kVf8
bjqZTNNbiwGh92U5imZ+hIbISoOe6XClpmS8TKDt+TH+B/AGYKPzRwdB9yjeKE3v
2Lh1ujbHaxsiLnFWrAGtyruGHgRybdc6v5hfB0eKv+iYapJQpdeCZFE4S7wrkSkA
makYb1gqFlB6bmC1/EoEzMCvmku0+m3TPdipgsUHNDXp6BpWYbZMWjKIWGQq2rXf
bGB2YKO4902RFKquSb6Nu4LfVMOhy2Dk1EaZyqEs+AclpDkbLxqSh4+G295Ze9dU
G0nRQVAq6qTvTCWlKV8flNMm4SICkGVVeuFNcH8kvUb1zjyGJsSzr4SfXNsIOGdI
F4m/kff0Ss6W0FtVbRosbxdv6/5oJBD/OsBsqrKnZhw02pyN/rWljSMLi3Z6+dHX
5fuArQcf6QeSUVTO4/h48R2MKyd9V01vdq1g1NtfHopXhGoPIWh3PAEit9Aa0vE2
w6enRD25zHH3DuivJfGs1te2f7KLBtwF/juY8FrIjdU7wbXD4trQQzRcB5KLpRyj
RLDm4AoCof01Vyzxcj6lSgiobNKVTQatTQiXhVywFvDiS30ZAQvdGPLut6Km5544
L+o7tCp/twqq5+ziQybfLZaRfnK/GEni2YmhW9avRYWdZP4hvHVUUXZk49yIzFcB
D+gbwnRkST6IO4X+ww29RQbN4BjHr2PMcmepVQVFr8d+IC6yju444H3NOEG1M8wX
qWoobcpSWU2g6enw2cqQ+gWaI9qyWF9ykaZq35daErbsXAVTInPW+FZbs6+Prro/
lvnIMu+f6NnnIWXz+PNwryI+otJqmlCSWdvZ/XuYeNiD0kmsYJeWvxJ1qRGaN8GO
nOvVOA6CwzBuMj5F8ujNIv9IAMIaWtsB41jlXvul4tVb7i7bwkV+p9jL2Z5Cwq5Q
VOSzGLSWLOVDRXouP60DiG0gu63C9OQqduAzyKw5TNi88kF2q1fmOnYQvOtqiakp
GGMEvkUd+raEi6ZcBu4/9Ef4O93u7cZYLzmNz1GpEw02BGpBaZLCS5piiAjW/EyY
a+Ei3VNAaHAcDhnAqyTkB3nOi28RIYyoo4G/zDUOh4S15oVAHh/T7++yR/fBVspM
kbxEPmr2L4ima0tiyjWmNHBxHyRb8yquvLy07Pk+kgwTjuHKA68GTiBb2Puwr95o
g4mokOWwk2KXVwKxMWRAxJprfLm/B5/5Jl68LzxuJCER2AYqQLB22FZCLYV5QdtW
PRIK1Oa8tZ1ja0j5V3Vg2HMpsN9FLnZL/utNbPZ8uaESu3OOYVgA3DczlNuV87ec
4FaDeAZf2HXPBAijTLfy83cXfPpuvFNu2/Sig3bms0/a/v5Xf6wCigtqlpYucb1I
tET0bqq0GiaNjyejZd4cmVKMju3ftkG2oHg696QZNX4wtpVO42o+5gkeMPNNt89R
cksxa8R06Ay7MX9LexbnBQeFgEQnus+QI3yV/rZb4Iplbl+ArCR1PPx5bNPXDYKJ
qpay5s21HzMom/PesKvNpJmpbcDCmRCl8AgWkyzokaBJw562snCuePDuZZMOV5VO
EiGndGrsC9E8ci9ezjKLcSF76OcIhKaIqvoGTEVGw9e8h9xJDDhZpjj/FyvD09wg
Uq7V8k8HFvyeoYvaC0D47nchmiAMOleRHGwt0xja4caS14el9WwV5efxyS89CU6D
9sdLL70J2rd5gyneKKGHfsLh2UpMk3YDPLUit7eYRbk3gRjBnp5RYUEOxxgEXgy2
ZAVjfKyXJk8BL4FwDvKqRjFHxDj5OlnhZmeVimvi6+MDCTe4o05x5LLYQz7ND6bY
iVeVCfmPcRNBzUPWH1csSIfioXc+IsVOftfbogpeiT0peltlXURuMUo2tsc2ofnE
JSAYm08PVdZgwGWXsLqSORfhR683tRIsU/kAFxMpMRKXKViJ2R5ZK+3mHEMfYBVD
goABo5GXq23B6Br2XfgyyNH4n8RqjJBTomyc+joYNfOg5hL0qsnG06dBI0k/8PTw
uHP8ObnwLyqpGn/yRH1aBCmTl/fy+IM+ji9MYulaeaxs40BzU1l+9uZ+lVCxfGRK
VDUPZONsepbN6NdBJh08GEkq3gejb6z2zNKsLZ/dcl/8LDscoJ8Etzj/Nd9sa9wF
tpbHodndaVzGY/Q01asDdTc+jikM+MjEpvqL9Mh/ledvG3lPBVLSr2ENGYYFTNw8
AYiuSqQadeEWmYSStwd1h6FD9khS6hppgy6lzQwJBdfGkb0EoAu6wsJSlcJ7Mg3P
MwRuPt8LWBrmNmuIGWQyMR8R0t9Ob3atYpObLLPHEkUc52Yi8dXiB5+RGZ0M8I/H
qKvpmx7A+57WD0JAwDgujCqlZkGYaGcXv/IeF7k2PKXRTIiD0XuV3AzhJDVVFvwN
Rv5TZ3KwtY+9OK7wpBYmeZNeoaYC846e04E5hDMKa1cUxqBnd87xSjGehMWbd8EW
d1kcyoGrR4Z34rl3xp4aqtmy52UdU+9FvDh8shzYbxrYHbu5EgsUBRW2mJfDhwOC
jagxp+AFdWEIuqbO3I91a4A2/55HaA+kgMRhrgY3w+iqKXO1N3plLirDf4P4TdSj
/0quLCvZqRDDgPbDnsV6VQKXcs0r9jFyjwZU3kx289JoBuPyZ/x9XRBg+uzpSeCH
i5FwDULmB1DOiH1za/I033z4+Li5Ny4XmiEp1heIHHGPPLEPHuoqhYvM3pe7U+pS
H49xvLihlLCCzIzoFqitNyxLRbA00Uc2MtTS7vCKI2gyQlgZxIbBt+QOiP8v54s3
Mx+Oii23ZxYz2F6AUU2G1QBTeL1T/Iw2ZXOqPPUhoAmE9S/ra65B6kVys0haQ5fr
lb6AA6CqPAh7L0jwPM7/ztDhzs15AAvxNM5jBk2BxCGnsr+/Fwdkoy0IBVL7hbyC
3bzgibQVPXxJE1tezUqlNQWZCZYEyLn3xH+tgmtQF+V0VJpEljKvqKjD5hSq8+Ph
UaaygPzDRvhRNd0eH0rh8CXxmXFKMiKe+tZPgDuBk7k/H20EdUMitlzxoN/yfWQN
9QaKSQWLvOWSheyyfWpIFXmjnUUFOXpk40ZV3kbxFMbwIxd3TSF0trUFOK8vj5d5
D71X6978n0eMC17W+AoTER9V55of0CBepap8fToyc9q9rNbVEovvVmEmwEBUSS2O
LmGd2jaGoAC0DhLiUxAR+0hE4W6d55mN6KryjSS7Z5iXvoPudcnGm2N0KD7Wf3V4
UrZr6P6yc7lpu+AeoXHwdUGW8i90G9lBy7gIlJ6fSDOrBrmApNSy9DGfE8oJrcPw
51f2L4WXl2mrBFqp2LxvaU3habJIoaH56mJLUo5buobu3OfVkxlRCW65kp6Ik/cN
C3kQi+ydqEc85CruxIBXtrh06TkZpesHOTKkqfkaVZOtLDwPn4q6FTmFRhQhHKqQ
4J9uOtSym8zCqwnozT4n571yUz7JlzGgw+Qr6ShIJRNEh4MXtmEh+Vqih3K4Gdzw
sVd05lotFG3DCo3LeOHT6Q2q+lrGhODkVJwwZEAybNhtE1j2gvYcVUkszv7+6wxl
WB37EQfhOcR/hPbe1usYUNGOa8/eAELhdmehpVoxj527Jw4O4pct8CADdYitJHmp
v484s+O+Dy26zXsffmJiUJ2wgqViT/vkijiAYkCrok8Vo2Q/w5U944iz1V9RJVYM
VGADp2NoQIsc9BQTmz8E7Ni2pSmy7p2Ce4PNWIEEvGqHCIBuZBGV4XIkbzsTM+3L
jLyuWfk1OkYROX5006C8Ni2ydH0/4xK6OBTY4Ex/jEWjrGjf2K36YbFAyyoLA7US
Y4h1vFUzHh+xbAcJ/7GsVy8I58MdwKsAojMMnQoWhQhYYmT6f0QlL8jH4IE9f1+z
z62EYqcLfU7ncxbR9J3n7BtsHA36DlKEN3qaYr5mxJsBkAS2CmL4O+6RFShVm00D
3h3kO6CjDXa/P30hvNCa+wyMN5nmHzL5Ikz6HSo/rOF/UDMQ0LnQVBxfnmxOXBrA
M+su2pDXTDA0zV/UdhqZmL4Trko2yzCoJn2jemuUymFjS7lf6ks/VQ174Qgsu+KW
qnx8nVqtViRybDxprt8hwXJw5kPGJUxlybXVI7MG9+KChmEsvIlR1kE3Z3djBVjA
nSv1rW9RNlpHIMai5jha+W5UbsJe2rJwTEnx3PXfNEORweRla85PIDbKKlFfo99D
rUwmppMltSM5/BXPgDDJBT4WMBdWA3oYWqEtBLpqzKHBmrjC85Y9Kv41tToIDdzg
JoZ9kzJIluhhSlkfCCrfeJsXnm+STUh1PSeJvE6jAggwoWem92yRoq2ESSlTvair
jvBeeHouPK4eCzStBMZUU1bzycYOCcBO5ht7XvFgEMoYbzKZW/DZGJf8Rx+RLZHP
CW2UTMXk9uMoau/MLW+MifTLl71pL76dK0MkwYwG97tERKRmVIbWAKfPXenM+2vQ
kxa3MDrBeMOmX9iiNne9zezLOWhAH5g9P0h+wrSO2FPaeSTt3B+YeKCFBQ3suDpS
0ouyRbHJmlNsQVXKJOwh+xMRDAL5DZgAD0w3EMMj5oug+KWsp4a2BxVqYOjIG1FZ
b/c4VKeyUUQWcpfleDkGqUkHZkwFp3Y7CzTeu9QGVIK9IXS4vYhm9VCu+hMiq/rL
UhMe70UPBtHYTGwsQ2i0n7NTDdDmEh76O5VS5iK9ZYDPG2ZOGWlOTHiwyhj9Trp2
lA4Uw2jZoqhyjFnr3f2ryHEnm+cg7U6VlXYxglAj52ko2SNkycMabHPEkWArkOk9
TcTvz8dSkAjt9ddTt/HDkATsJ74Ea/NOYx8HoMXJcd2Z1vzVVpMrAKwe33/zQtF9
ph6yys2Ug9eqHV9MUxyphj3NckUQ8rWAm7FtSoS8OK5jvjVEIvbmtDAJJE1dev9c
vlwaIFC2QjjyBc/g8yF3UYImpXPkhYQPxRmSAS7e64YanS1gKjqaBvnbm4JaEVxu
QrItE20eKWHr7PY+A7zSX1mqbAHjhfEGoCg/DH+0xWZCAu1Qxq6fLOl6LW0QIX/5
kjpFxIOau9lthHxfG1YZvDod88ejQlaKfeRf89bMA+g/oyxb2m1ygXEzeDc4eeLp
x86odpJZfua+yg7qsj9WHF/Y0PKJWOlNy7AckFj3JiocVIFdB1opt2xWoVAzG9e3
+DhFAsfEszGkj1mzbkOyPrpXDiXLGVRiKkzke769Xrx84OxlKwPAu5nTJFhmWu5K
GvzRWxNMRSPNBriul666C6tbyorpNYol18h/D3Do6Ofg7uk4mtXbprrhXYS2UDzi
RUJXP+6zXvbUneS8E2/Y1dn+woHSD5sWrK7nlZvVnWCB2sgzqBhgt7uN5N72XJtg
aQtumaI+IKmoW0il2ZduS4CXYZMxpSq7oCPFmueX95nIQ/KEWln1YWanXqxNphOA
znCTres2dcHM5f2cJgkWClmLWBug9E2ErVW+yTcDkbKYK25JLSlTHN/92kaT/uqJ
oMfn8KYkfbTDwZS+rU8SZ8Jzu2Ayv2Dhy1FhdCnzhN5pN4n/I3cztBmudhnm42m/
WYRpKKkVErrHP7G+BfHZ8nlCLC21MyO1AS28eCdhGTKCxN3wgY/Dnb7zChYaq2XA
+FE/G82nNp4RWwtlghrRPJc6tLPHszA1cknwAOUeTg/shgE4Yjp6/js+Vn1UcAGv
ko6uAK/CcTSNAi//6XEAdcPEfdghcioRi+0tmoAXTQtSFZYuA0Jc2U2lfyRkRosL
1HUfKmI1IocHmOa9NNPdRUawHIrLMqSFf8KukuMgGDdRGp5xj5M9jkgCfNrI5ajT
X9YAmvZlY5lpd9GbswWTNdTAYSbTWvfcu1SxAhGKY2RMh6x23gS1YeI/Fzhks5EK
6JCJys8QRjBMcuo41AiSVDZUHegnYJKSWMArIxvZwqLo+F966MlBSw9MUitNpsHh
ls8OfZ5g8TjM33sxTgDV1aJMuvMsz80B+W+2g4WSPPumHu71x89wevO4NodOB4Xh
y/zLm4sAquCLeotT7Yorr5TdwySUjdVlm+eRTWQk9G4JoxqP/14FCVdGQcE+qrX0
STUnkk9ccnnHSQ+LebsBLvn5+J2e+9qrw/0JHxoyS/JRZOyDppD1A2JCRh5t0ENA
xl+Xe/PsRsIq76kpk6DTSSoDZou3QTcUPtc6LOWAmy6V2cOe3h9gwtMTLGgsMz01
ZIb7G13TpUtr8UpMDJ8EaqXZ6+8Rd9GfWt2f3OZUzj4Yc6wtJ5jnWld25UEXX5Qt
RrrYcc7aqrMPj3V4Bd0dAG7dlwMYG10Y9r+ISDeAn9VUnksY8In/Y3t65DgAIzYd
h1NE61vWcG0yX6G9zHbJiFVmyXJv9iCH65VpXD7ZXyjIczWa5FwtVWru+cQycBtc
cLt+BFAbtFWIoGbzFnrzQbPRe0eV778ydt5SUIAsXOb4Bc8+32NUvWOtZjL0lB1O
1fZyNGJQvv0Tegk58XsofovIvVATArqRsCN9euiVqqS6jDkrXUuPFjCsf9YwKHYK
wqRY39wHZbM7gEdo/f6E6JbBOaWf+3PWGlT2+ZQHklS/4OpbMYw7e1Dk3OCJXrLX
hXUzGF6Ek6YruL1GfdRf4ctnbYXRmCqHIfcUfoSQBXUQhnNz+oJVrM+Ilw3MKlVK
L3xxQWIUSsSvMw+7lndvZWDBnto9xKNdz/mZQF9zUGczRf/Dv/i+Z1d8FGmxXi9/
a1O9uuEYgQy4mxx5jd2YeEAwF+05iDZIg5OP+569yEyu3vtLYPWrPkdqmsX/83KL
URzJcdxi5oOp+9mtX04R+uLCJC/JoSdQaUhawQWQSqD0U8bP7GJ7oGMUYZm+0cf7
rhQxiUWwCiC6fYF7cVzRvOJoH7awPeDAC9PBHsez41f94mxv+IV9k0dpKetBL1VR
aGvMsCyMXJT+PPUf4Po6zdA7EpKkayDkT+86cRCj8ZiO0aklvq01W8KIUI0KW7sp
E6vhiAgEZx7H9ba5DUBP/lGqqACZakpKn1zG9K4GSw1TVpT49JYMHp43+EZBF5b6
+3LEBxA8HS0AJB0i5yuEztpmKOAw/g665gvHN6O45pS2cM/dWW9XqTRMg/npGNFF
AZ/9KdwxgnFRWVfbSjw8h91VtkaDdD1vBNx10vmAZw7Nv+exCLhCb+Tw3NBONuKO
P8w+X56Ds6WPb6K5mNXs2NEu9qbOOrEnJyGyg1AsfjV9+YsgKCbypBEWmQqqtm2m
5z/1dCEKZ7wLKuudWjz2xA2VVtVtVHPAh6DdkFr99UsVLN5ImdWf3pZ9ZXRu15dQ
mg1dLiAXfmIgDQaGs+iN+EeqQulXtnzSkVO5sVQJcZS43pmqng6d3YWhyKAYuNd5
q7yduOCPo0qzHJgVVuqOdcUZGph91k6q0tdMhNyZv4sFS1VJ9KI7rhFFNdWEofm5
hlAXDT3gh5Dz2ODsJZaMPVERpb01GxfKPPPldPbWugPRBQ3/SVlUh7nRbM2r4xs+
klES8CiaoG7Qq/vj28fSUmqViPlWjeXjfNk9hLMEFQ/ZN8kbRCZjl98vxAg4Ez9a
HXuTu9WI0AHWIFLuwdAnRJqXsOfAEs0Z5G2GAVx+5JoY87D0R32LLvPpeAdGOTie
hYbQjTSxGgX+J4wRMLZ5Zr7fA0acqXFfU4uNudm4E1RWADjRxQQQMtHwMY0Lgjj7
gQ6VkgqWBRMAWTImqCPUtiau8QAO+yp7+MjZwgAFiGx5SKT74tM+M390ll0+tz3c
IW3dM/Wm3cBs5Q/AG3GHHl0dkMdIiRUMFEx8MTcf75VuA6JvhQweXq9Ef7kJXbxr
J5wZWXZ4H34Vgm0OaDhutoCUnthnCX0lupwplkXvnbmd8yXsC0Oyt+zuxNIJPqBI
qyfDilJXcBaWZv49VQPE0623oJxLfS0I/Akq8St9D78Pvx665XafcX3maNrN0UuL
GqeY364hJacB1xrEWy/bgjEPovr7KHYnd2Lm/Gg1iL5uyRtFOfuaajh7nBV7jGWL
Z+XrU+4WUzj4cQp4yifnWv5UQ8O4EBMWwFlffdB8kxrxwZhtiaEUQLP+Ud1tAWQg
HhktOmjF5CAgFB8SZSi95QzpVnB8DrV+/wmdNeF2Opcj1YP1LKGuPt+VYXjIDZmR
mcG6SFd3ZMBGaeje1cUvyejO01FSx/JYpQe/O7dQnx3oa3cZ7WXLAf64fEAgncH2
pmbB+KAn/93YQFCkjottc5EzX9JSV+hANWjTCcI9u32Gqz4nVrFAo/mfYUeD2Vuh
ly794K4es9ne/slSdmbFeAIYERvxFK8LsB01zknXR0nEqTeJDw0gl7i8yfuDTX+m
4Y1mWZTD5NHKndDTU6SE3wWSigfKCBoEoMrpORojJlE4/5Fg6CgoD9S6tzZxZU15
ymhnGgZIFqSFtkYSTep611jDJqdLWerK4DCX92uIyOxSQp8hbVFxd+WirQFVwrE7
5RvcyHx/UkY8u32M4iLB9XK5lTFVypANyVoLu892EYhBJjmzn0opL1+PFeuABkxV
ABhby1C52BhqGLynAsbfsxr0C983krNEKJhxGAmJblSZRhoXa1AbbiyIQRthWYfS
riJuREpXUJx0PhT0CrvHu56tX7IRHVuZoxCjrSv55zm4caTiiLaayvKot5lBhQMI
BBsUyQhXtHon8i7oR94B5wRXxDi8x9fSZW8EVAR8+2QMors9hd3HHZA7LPTuIj/3
Ssv6uwdhJsgaFdni+cHvoWcLjw57DSsLyugStWACUJB6lH44+SCN6jjEV7n6GKnG
1xMzeG/ap67lget9I43YqJb/VE3frBenjtLnpbKlI9mHzPTaQVFDqcvrHKu2xHwz
hiC8xOr8Ygrui62r3yH64OiOaROy+RLVTnYt3ta3662Zw6R8UO/wHBQsxlxck6pV
0wKfv3l+b1T/v8cuJLnZd33Bfq7o5JxR7usLEXG3K1J9uUGxwWZaMYUiCWUYFH+g
HlTIHBA8IF8waRuvpy9RUOfI+Cy3l3T7/KVNUH6DmiyfrSJryqoHrCjZB6HB8Cp+
54yqZZUb97+ZmGcmJ9DdwYst7x56jC5V7XloGBZMpMynCbL0qROWjrTrKu1xoQ+d
mXO2yEalboSPqIoqaMqHQC8HGHF7ijuplbrCXEMRYcT1LqnPXXSqb+NgFaNAfhk4
91SkLng2yhS3t4FRn5HT+MwBMx2F6hUAjEKqq9so239Xu5oLVrjWdc/dLNUjPQ3D
MzYRJCYWSqd09au9sw7XQwr701fMCdE7mXXb8FdvH47MGYu/UE307zNhZj1m7KOZ
AElg3NETYcsZ1g6hfYaRv95gV0QSTN4ZbLF8oa/LzxFm9DGKcv63PaE2z8zpmJf/
akaIX5cMT01hPDQ84Y+IKJ4ardqD139XIhoJ0PqO2BRxQXbwZgPrXkGXWFMcmSWy
uGBg7FBG76P5Usz0kVrNsIZcnQ+TlxiYFqx6s2/rlQOW0jTFQn1o3EceS+2AOTnN
R/31HL+c5gGWsTYrFEi0/xs3kzvf3pOSgGJcl6HIFBjw3ON+E0/0B8y8OSeMAz9o
Ia3hxTrQ3g6FGQdXgSs7JnPWfpp7MB9dhyYhBJJZeQ08pX5VrujRzUGTZlU4obmV
WTvvxsX8lVTo6FjnH2AiV3Bf0lBS0mTzXDY7Pb0fu3SeLjiroMToGd+2fZe1/Y/Z
VM0FHw5eOV1oBELmu+tRxlAHUiRVINxrGRdhg/aQVelD9Q6RpojMrSnkzmB0epEM
wTnh9fxbeScVwnIBiLcjYrJmzmumWoh+qbTqk15VH4Pqy+C+vZNYTtGIqspLGrY9
DISbd1Cb5cP9ygJj2rXGjJlm3S6HjiCuV6lVdpL/TxzglCjhEkegjUUAc0KY4Idx
ZwIIyMTPhnfs6rn8Hxwzx7X0rGcAycvJs2G3uSTjz96OeE0rKBJQjhGsL4ZUqhZM
SfFBXSO0U2LlFGYiWi6WeHVyQk7bRoXx/osYQ0DfyYNbeDjznx1dBBmWZno1rL9Z
4T5hutyfRwombIOnDX0uvd8+lVacanpyx0Jv1neKRM+e+8GoEiIPa7E76I+zEWKE
aEc52msD+RC0rgvxx0F2k/rZ/x6O+ZKC6FNTGV3tSnb+dKkx2wiCq7xsdfZ/lwHs
eB0hpTdteN4TQq5ie3KBBImwaqdfw248CgrKbuSOkhOfoMcYJmJJ+qjqMfB2hdfD
YzoTk+GxXKbDJY5ct0UKTTvI3DNORTCqdhsc87Io2pA0DicaCziQpHAzyGZg0vtw
ZOSRYLIHDRs7n5Ub/v/1bjwVVbK5QFG7Eowkd8vpJviXd1E9lNAyaSxdjHx3DhLA
ojXDe9Dp18xkWBQHQ4jZ6LZIU9RITPjXqO8vYvWHerFaC8OtUyEuIRJomltjsE53
ybNkoekDjsCuIqeQ+hym+mOULpvXQjjYzbXiyyXRyerGU0POQhQZhTAO/G3aO+36
cHTBsaIvVdZUnr1OvyQ1PUJnI5fLhQHEjDTKI6qqMXlwFuuylcVElS4+NTHpDexi
lfV1GJFXAWHJj6ul9fsRdcBqWx5nswQ+ZNu9GrsZaevgaYLZwwNp+CPljIj+L5cW
upBaaDa/frNlEUVXSuR1DtMlYSFDElsskmqjnv8sBeSK468J7hl76LrZ5wv2FYVr
DRvlGLIDsDu/PfSeDznbn7CjrSECfYdZNAIx+UBMtOMQMEUnjmQapSCTEvP3UeVX
T63KCJzA3cJj82AR7AN9rTxYm6cu8IJfUuEHc5EAi47K80lB6eiWa7yqoORAf6bI
B4JDHLnM7uRGeP/UZI7ab2NxdKml40gtVnvSI5IKICQQ7s32Hzjyvg0yCjy62/mr
tChFT8c9Pmn3oMzCV+63o6KvXjhSUXYXVCntm9rc/h2HhHIUq8snLQ5G4zx2lNA+
ZVCfFadJahppBtVPDMWni+wYZ1/sOR+ejeVSSYUEhxUg8VIIl4FKO9pNUY2493G/
8iDvixeYVzZNNR/2Npjt/uiXJD/+8pyDH+V3Ee0fPCrDiJpKnFv8EmRVG5fQqEjp
E6KxyvxEHNNnkqKLV4UKbf2b9YgSPL24ewqVd+wSfmYES/QyCTB8ogaA4rPOBWX5
uKxbGIqFwnbwtfKAZorHigjZj/UnYY224XvYFXu0qvHVF1S1PvX6g65fyoE1mv09
iavt9TocPNruKCS4ly7h7EU+eVkWHoDtWQAhpKSa8FJC2ThcowPKyA0WwQm0tZau
2bMQdj5t07ZzJ8oA61s2DsDUDH5T0w0Eym69MOPmCBll0KV2zurMCdwRpzYdIKQC
Z5AFnb7RN8kW37BCC3LYFHMujRJhoVEAoex/NBiWsJd73p/h7EysvMnqP6lQhnKz
pcHljKnjc9k6cjdmOrr40AoRQvfL9YcEQXa4GGa/mJUA7qflTFOmxt6NtBBICJgR
af0nIid3ZdceRGy+K9ScS/roGnhT2r3ZtimpGuA+xglAGiBRRaW4z7RS164ieQN3
GbPyfWHU7h+4KzM+YdSglB/579pr9pY2Wi51KVnVHH/tyz5I6H8/hU7iBMnyUHEY
EfPm9rhul45CTKm7mP2Q/+9pwFbE+efD2687ERQuGY2BEHxjiYdS5iVDRdQ2CTtE
S+u8AfzJ0+Ld9xnP6F7YRlttHUKDlwhXBW5aq8vcwnAo2ZVbwt7cue+QRGjNRBGL
HzK5ByFte5tV15yL4f3c6ZXfy0FqhMOrqJab/CaRpVskXavBAUDF0nOvHl0+kFE8
5Uw8gh9A4YM1Si3OBf3Dowbji1vmPdwe2zqOccC+e3wTqmUxwTVxJHfXJtn2YLk1
fNcF5mE0wDfTz2ZX3tun+0vd0ofsZMmKXnyoMLZXlSVirIh0JqvfpE2+y0h6wNur
M5ievbeI/Q8qOTsua8zlIFl4CZlxGaiFZuRF4h07CFptbLNlza8ZrEdL/bnJOZ1U
20ui7BUV0wm4w0HC1gM/Mac0WxjVccOXASMcDzgKNIB5wGZ3g7vSxs0ubT0nP/OT
AsezPP1HIB0rso0t+oqEgPzWBU7IlVjJmFdGhYhZca6dDRAO45iEuZpq20FS0/9u
cFrpK992lUvVTERjz5JiuqOPFC2mfTAq6RjSvc4JyfHxXqNByzOvCrGIE544zNlu
LFZX86puhuKEp/qctdo5Z9zOawCPTO0xr1gC5+WUsQ+RF6Y3xXkMg33HCRdItcsi
hnpHTngMafeQ5uf5SZmF4zNc2LQoStjGY/BIBl5Ewu04WvK7oXRLm2+gV4wKPuUo
u5AvbpaPPrff7zit9qFTvlw0wnnm2xOOz03OSqKVeVOXEwqtmiXoxvzvTSUlGGIg
BGuuWgyn7DdLVvgt7vpGh+eZEzwTY+JMDwWLeBjMpx5axaWLZXUNo9bwhYpW2HnO
FglpU+38lqDwu6kkmIRpi3YAZdnm86xwxzXxeN4ALjZ+Vunmsj87ce6Ft1EQanoF
Qv0m9jkIrAA0STsmqzPbGlw3z7Iu/GJSzZM9psH8XqfSlIvsMLv4/iLdqqLoWq8l
Ew+9tglGnMzELJ9cWJuMotcOXZcaYgbYebrhxL+CQTSLe1vgHGP94hE2QLLyvMpw
u8FYaxKO6HKifweP6w4TgAiQ9q1HL4wZYIST+ugI4twMxfZ/F/60S5qBRQA50c7q
ot/JIkhl5Ym4EKoS6MVjpMzFfszepRUJ/1R8UBuaoBX/2KmnolBuK88Z2A2cWZZB
vj2qxb/MUQwT898AaSIpXpeKKQTLnabJP/Og2PUHNrJgx6t7XtzK3Kh/s9yo1W4/
IbqFmgtE9kudVoruNZoBP4cp8fs9CziBzX2sbuP+IxHhhsI+CSKAqaObN4kZ1AMR
buslLnh5CQqUD8X1e0FqKMseZaHEOkn8n3qo96QCr5uOvFH9SoGXq0loR8SifKyI
NocoNOsX9VNez0gwqlJanEvXOOP5e4UCnT8V10mLK8dgabmD/QP6Q6pxyYzGuCwz
ze1fdz+UFbfR/+LqXm3SpqkvK8qxyrzlQhfQLHP33e+ptzN16IMXHlwUEZfiGNJA
WNjoahYjYbHmgz9huOVAy2bm3wZi/MjxeHYuMFPo4LIvWpGrSg+gzCW5bDJ/Kn55
Tgkdom6d1yB3alK83smag9yQ4XJh2p3wqv9BxZE8s+R3jHOmyV0p2kRPhdH+sQOv
ajhPVh29AM0N42Bkls2FAqZwh4pp+R4+9Jas4j7+RETlvZXqx9frpvBUw3sTgbSW
LxsZ7nwCkg8A45Wi7ML3OGuCBllEiYcZNb47eo4fM8bWxEd7zL5mZUICIOZc01q8
t/ZOgciXLhwmZd0/GHo8b0s7c/gX3CNfxsZdpJASosWi9ltjp5OwddLbhSajY7Vj
Z3SFuD++4JE/94OAiKH5YxMcenFbtcUoEKKg8sVaxlXqGdFbHZyZeC/fGItXDcKK
/lNHeb9EJ/kLt1h6yu8nq7MeMFyD7PxiszNSgWLNkTXIvLUAvBL+lSSIU2gn/5T/
gd0JSa44+bzoh9FjXgxgHup++dJ278zRKjSWLfk6eu/Zh+etFZhhBPfxxEVGvG0u
0Wbv9EBZZ5FtnIPBQEYRKntaCh0LwyBZX9p8nM2wyEAo9YRc18NelnQB6IC2fw9b
IPqR8jCL66Z7dZt/jH5Y8nq8eb8wIvrtwYt7xBaDwzV0106hxS2MKesAwj+t9sw6
PF9WHdgcaI8Hk1YHcVDhoP0bY4a6OIbrlY8bnKMY8Ftjg+gnoZ9R6uSOEIcuonV4
1U2lD8Bbq7CNhBjPGDAxxSQbDKiIs3F5qDa6GCDp8Y484zyPHRAOFHQoAr24V1Hk
/aWeuqggHVpkg8q2qBnuejA/SbHd1341ZXQshVdKzaCY2yfKX8ZaJeZD/tp9FI4k
SsX1sSyZqIyWCX2L5/g9gU0VnFmmimLsWg01TJWBX0RP6dxWxn4cupXHQcvO94AW
bzNsRO4/8/XrybBvVsYUkLEHmK/FMpJLjNljUQFvC4aERsocc3PAKQD7bakG/z/y
1gecgucuzYRTmE249K3VTpQO757Y6jG9KQlpgHN0gS6DCBT6j0t4d/4jZumzx+Ix
hZdfNY7yhhr228Upa9S2B+h+YTrwWsyumEecoKa8lCmzznbjX8pog/Yhwydumxa2
XpcDFzKA6Pd4f9R66fxvdOYxIF1wBGJhsS6WCKpD33Yrhy4ShIXicEXqAm6TQL6O
VtUaVDHa0BUW1oY3/Vwq0yQCmENjkW2lr+xCW0WRXsv88TpWOLIqLTqIGXBGK/cM
EZR90SUWD4iWPVCI758ToxYG/IJgjOcbvRp5Ap5ZMJKxMC2lHeWXX58vhpFCB+g1
7fv9o2zqf3j9GtcBg1AfcaXKM5fAHJiaWbppwwF0FcgPBR1Tx9gsFNiIyePQOgUz
8LvTCA3UsjT0fymqaHeYiWkLrQk+Jd4ie4Lb6YdVYCJRJfZlhR+otDcOw+R+Xqh5
LL22MFx5l5VsF3y6koUfp56WXaz763zRxMzx/5Ur2xDiCH8mvnYV99WGuCr0QU3a
yZ/sFG9fl9GxYbZ4GY90lixcFjLOsWjdXyVUTQg7s6QBzNKbQ1rNuWXFBW9jRIR5
i6Fi+NbUCMHbqDNZWaWHBY62XeOvKpwKozENTzUgij5EGT50f3rcZAdpQquzQmV3
BZMsZ1Gx9qVX/3TbLkcKUR1dXI8p1ZnKzorVrSpPHLVSRZQCI/eou5Xotit7MwRx
hYXyDan0SzSZIBHG0zxD23fUPCuJImK+E8IGc5uk5lMX5OyOVMVtUcDrmYWT4cwj
NYyVvS6JKjlRnSJDxB4kI9VWd0Xbr+H5jVTiLd1sQ11qzZFfw9mFT1zDe5KK0je7
aPmkvVm19d1uge70bcNzqefanLQCp/KN3AUxMzZiwOlcosbZWM7FEaaB2RA6wUrV
yCwmMArdiRQIbg1Ja9GvLBbr9XniFWLEIp/mk2oGYhwBrW4Ms/xBxv3vvIp3FdI5
hu1dIrAx6oLDEuXm2zdo6gChQyMfx3AxRPEjj3IxKWSZhtsjKw2fJhtZDYBA5OkA
ZgZgZR6eSll/CTY5w+KYoQ2bWfdmJ9UYkZnIxSCum6fm6uJyW3r6xfF9LhTpYc26
GgL4EJUXiVMU7awLaroFNEa7ESmE1BU2LxexaXtXigq1+NQNY6nxysJ8mSR3EJxq
XDNbnJDqxMx6IpZ9S2gPMondQaHw3i0/TwEcBY5siyrdvVNsdsNGGG3yGhPU9AGT
BigQVkhe+w3H5Hkx4XRVTyrSIh5f9p/5LwnJXg5/jNOFWziykokxp/saf6Eqgzay
asg5M+GnIqgQYf20tqlK6rRbSi8J5lk3KwMvcZYPlbpCE58qmcV9ZxxBTzAT/PNg
pblfnrslaXt31z/qaf1xUQ8TIYlzXuV4FmZ88hDZGmv5NWUalrArHpAUSMZaoTNm
cRKjGIoUSpO67WPM125joOViYw6gxXoy83aSSCMqw7BD8+YtMmC3dQbF/g1eFCVm
4sXgjwrv9fbLv8WsXxqU2beiOfKAAksjf8r31o0sUybTTBkyxq5x5P1vChvuxVdE
6gpoaTlfFk61VTgI6zuZCyEOdqgBfmGA0KCQ3TSQCBNfUPm+fOe6OWMjAsOVrBpD
vVcMSxQs51UyPUW0fu3OBpf9kpEk+cbnCAe00FPQeBPW2s6uj4570MEhUCSDdmNf
FWYnRZ+3DfyEU75zg4oOjFXdC2BtJm+YkWFcv3rzR/OD5RHAd0qbz3pR5s4ADjvH
sv9PZ+pVsGlm029NdHRq9zRLzond3T0gbk1H9h708gRL2AZX6efd6YZXrx93FKwG
pZbX93ZFPDEEQ7yDM6qkiRKboPfA8fLp16CcFKKEPrPXMExfxaQTBaOjE99INs6t
PIRnwXKpZ4OgH69RG+pJil4im1J+kWBabbjJg8yNrjZs68PpG4Eu0i4LLGHkZ9qC
5hnTGRcaiWU5vRxNjftUDBn1iUxBzVxpT/B61XAS+/nV6KuVeWaT8dSrQO9wfH/A
aAQx5xYIyrkvcLpsu2vi+IzIBq3OnaIAl4VtLwg6mD3TrEkF8vjD9FMhVMtJxnsn
p+SqeJlnnFcNOmqB7zctnAiff45wP8h54+5WhFKltXNKy0SW4b4cUXCG6t9sNWFZ
k3CAuA18c69YN4IhhA8IHxA1n5UQxHPbqIWRvJEaVAkwu+HP2++RWmkam75vtRlp
xXJWEhBtZ/hMPIAHpkr0vd9dbiBu9IW8oO+kSyU3qy0Ex3pH0KOwK+t1IuJlAphA
n+SewxE1S12HIxMlze+/ERe6QibI4aa+xDIuZxQmUGnxFaSZPtJjG2ZgicHGYoeo
bUUZXh6QUFVOigl//IFEC5xZlPeuDZKEJMOrL1yY3gC+Efrlx5NEtxJW2XAQL6Oo
d1RDy6t1VLBWf7oYv0r5Bu1gx7iKgTZPwJ+3WEdQ7MukejNIuPjqQlmvRvEXqdfR
UFyWUvUmiIg3XdUmV4fL7T5Zo+SSikAx7DSc/FkfgNIZ7c1UIwmp5El2lEW/pLST
dYXcNKqNN8Q/jgJsN0pp4O4FbY6tNKJSgoNIsW+EwuWU3ZeXFMcAEP96NhALwwYA
g3xLXlKTL/qfg1FGBW+cFQvkpqFdYh/n45RDnecG4dxFHwU6jKkL7DHCltN9FLA4
YFMoZcTZACPyHWllAWO1R+ksi5/HbbSwO+w5ZOlIjlDMK9sLllqB+yE2hmAt0vdY
Ped1kLnvTWApfcxFEIcLMzUU75undjo7s1EnsapvSGTucJk3xCD846VtU52yy/w1
OAXKBHzAM2RhmBAODvxSo6NVeT1X6pzWPCayjwqYNjwyhvOaj+PGACjbSrlHHwQC
FUFz7Ej13eCGI9BvyPWPLEmSpNjwTredohxCBFzIQeIBdOUcwGv4tqAlEi+E1UbH
oEyRSmgT3HTMnRPlPJaShpR/dGlPsCrlAe64PCQpAkicZDj2vdbFExglq445k4hw
G9HSAUooo9AsK69zBMtmyBfdelUrcuq3paimiOBW1TnN2Ujexwj/L7jtfBDUgSsm
OpXnzmcnKbwSuXEMxstu/nUzt4+WZIHW1hNS/sM1bS93YJJQVqpwt4MZ0SxkR5iQ
5tXNl1BJXuNySsDvCALZeVJxeWzkDfFHERqAO+I68BEjTiOCNsgD3JqxZSFzPWan
wlpaXu7NR89HFfXRh4zcCi86sytxhkQg6qKk7NAqrx54xmgQF546+LWInSD43bsh
BQQs/8waVlD//Mbr5nRObIZlnhAMLDWuqmu4XdSvDEbNbqnnABg4nOXoSM/cKcQO
VFifq+xOtyBkhzPpo+DchiRqcAInVjFCv7g2hX75ofm2G/BsdIGmjDO0g4v71BQA
+awdYiT7dwNZGn6hzoR9kFWr92xLkUebDMFhhYpe2Yu/Lr0l5wyso+25LD1Y3XTh
EH+ScR/L0upSpvcJdgyaXHW3l8FaUqsTHhRbm6ocFB1fYxnw5BJOOz49zBefzkpe
oweyoER4xx1JSwibfbSwlSsExhOOurcbKoL/kem0eL8Tv/EKFM77QIw5ywm4mpJ4
PIVj5WvnmHKYduTHjwBRxk0a9nGcnetc3QJkhVfcjQfspUbgnTXSxyv0ZG3k6psp
b+59kW2FDJX46564VpTyhduBtcg57DDSGhgj1m3AKAEDxnalKbmF1gZX7dTQnu0H
syITwXP0PShEQvrRggchEfQpmOnnUjVUXCR23r3sFPtvM7taHEhmgnTSguiiLUmd
nDwDIpZ29KUp2RYQ43os6fuApht7WQ7XKX1grHg6cPyOydhM7nufW5ENYuRWXwI+
/dBTsjDOfSYyTAq7k3X+V432U2X50Pwy3la1Yr9YztCcfaOB2ExONQ8EiO7cs9ld
5EhEoKBXemuooSp8x4sXq2RDVQ26b/6+7tAYsAiFs0/mPQlB6srjgr2ABoxRoeUJ
S/6R091+ibksKlu7icsTShJkq/iU8d6E/UO58dkIrFBykFVfdcgSHzerC6b6XRnA
dRbRTVbbTI37eUDieR5aJfUT+GlmJ23iZ/AZ/C/xOIc7fV+KqbKGXBYLHT5RulTl
c9X7/m9UEGUuu2Inc+F55jjul7Cots+8LoVVR0wqzh11eOcD/6CNGY68VxJyruU+
z1H0ipV/safFNCUhGscbYDIcdf7wSOUxNcTOVhEJHPoQpnk+vz8tAZhMea/OFnlJ
EX5TiHs9Ey/XZFc5hXV+A0X0jhnDbEazQULTp1cnpkEJHeqok9jZu7d1JwO2Aib6
Z8QAgU8Lsm3rrG+YvEJmvs/Ca6xb5XFeI7WV+TuydpvRdZ+OsFS2Jjm/dhKVBH8q
DORMfSdGNFCH1YZoxjGC8UZYE/qsYU0M+VqeMZH6Q6+pkVb838SdLvSp12cVUl4+
vwat0pITOo7AFs+6chKOyTIqLkwFt0cjYnLuJN+uNJfftk8z3T8sot4q1Kr8Pqkc
wbvJQz/0iYNvVo6kFyYlKYtDHiV6W8B6lE7RfV20GZK8Q04B/6lEuIRsXCXwQkeO
oLUqHSxhMX0y05BT7N/NefYBFbNOyNeUrQnCecEL3b/9oa/YcqqFDLKYRf+rJJPO
5U5LbumUezI8extba6jnhqQSimyFhXwsCIqNQ8+O+YFytn4cqVKGteaIcSJHSyag
YWp5hTu38YtU+RJZ84d6ZNijPJ919NVe8mkByZbRpyAV9u9Fzgo0/3pb5CQjP9Ja
BkX5Z+TYIf99wLs4bNFPYkbmA1arjdxpvxE8/6Kd0sDULj+MIFnC4deMWu2Eqh2C
//1/v8OAqRPGb1oSg9A1Lbk8lWBCwW2x0S6dCJevceEXJuenRLH88UPSzTqS9/Wf
T+3KBn2pkCGr0vAj7TltiNZXer3xpu5hfmgPrjTpmcp9fccFjVwxGKT+nuj1xfG9
Qe9Zo/ILhuYWrFlKMIKQi5+ejcf0fupBsbMkpJQYv5/XOAuC74g+DMaARl7mVFRJ
GuXkyJtDs6UVQ1KCKZ9uUDkfnr1MBZLhtWMVTCUtZ0tLyjAWQVzSoxnvoyPPz609
cTEN4ySNLWEEZ0SjJzgz8aQJ6vMID/cSEy7yjRDSLa7ymX4hWckVQ9A2JmPOld60
k7rMDxOlRd9VQLdKb+jaATFbMywKzenIvikltn9zNpugxZFyBAfB8y5E/0MPECN7
39JeGyexclcNQTwi+J/kqJk6HdJkPjWseJdqLXHhwDHOwUp/kNsp7H0r4LtLQP43
bkQdG7ToWNSQv+XRwFzFAhzsO0SArYy8vFjmEZhOwKeLBTJEbNQjxW6jpo++WhIW
M2iD78LdLyOXaUNsuhFNf0dy+ZMDZnDQtel1Bgt/M+IthCrw7zyZ+27Qn8Prv/Hr
FCd8dVMudCoo2DDY03wZZBcZygm6WLOkLxVav2RvltdhaYjxqDshVR++bKwx9IXG
NoKZNxTvt+B9Jh2irJeb6u1pXc5Z5YVZkl8Canbe31Mg+s7PDv5X/lddwIaGdtgu
hkhWpm4FdDLLLOTTAgcOyFFVP2HqvQ97mCzPK73rZh3aMFQ1S7lT5L4yDbdx+kQf
WT5i1xAjwoFDPkQUPBJPhN/Eb3TmtarERs7D1Kjmhw/DjluFN74BltkP5svI3Eom
djZ0vo6z31W/6KcqLXHSOw==
`pragma protect end_protected
