// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
fDrK1v3IXxZ5VX/jcWK3mOsl/td4daKnsPF5X5xlCUkMxijEsVLT3klgAlMbWjLW
WcYJkAGFxVabAZ3/lCOr4zziyM7JYxo1eTsO2HYQk28iPWDCZLSbYCT06thiXSNN
x1rrSEn11+j6/Vo8s5frkpGVV/TFSS7LnzF6UqB8p8ksMT66SdBeNQ==
//pragma protect end_key_block
//pragma protect digest_block
0UTvVk31CpJIlJsPyZ+s5SNnt/A=
//pragma protect end_digest_block
//pragma protect data_block
qyRSpZAlpWkQjeDb8DTyCE1cnDjyrP4seEpxfhKc+5zsyYM9Ys082qggeLYvpy9L
Wb/CoFGruiopev925PUbYKXJAiBwbVIS/haDiv3y+NrbRRngFLiyZf3EBK0evYR9
6vf8G7YcD+pEIPQDpKieopjDA9ZL+i3MDW8HOSEC/ZN7CCrlm5Hs1ZHMeN7xgo0t
iYJ8nYTqb/UVp9AqZkd0srUQTaqMzDPnkYZCWKOCp5fX2uKH+hN6fM3QVPVZFc3f
kltjYV+2Tfrc446pJF5yYvn8jV9KYz9s3lcvUTHSQHY7uiDdnpAi8kqp/86dVaiw
AjoZBmmxmBVo/ZW4NrA8Ub06A65TcI6z3rh/ac/tz5EUM/QBdGF49a+mFYN3kX0M
Z7Wp2HkLGMBRIJJn3DGaSyyHF3sORiy+oUbMRm9vIscjvpjaGZcWo9wlvKYr6RIb
4q7JKlPBC2Vgb+iqI6CPqC4LRVukcbgdcRPdGOLVOGkYWYcWLcOH6anGSZDbnc9m
wxp+F8rBczLCnwXeKXb00sNGSyRJ76dvTyohS2BI9rOufhQM+WqEUYVJXltB3G0I
x+9ZNM2V90BuVdKXa4V+lNZvM9xHOPB+SvXXPpC5kEABs7sg7xwT4HdIYEDp1R0y
Qq0fQsZKq2h439m5GgH6mMof7icGgVA/hk0+lfK6SG0ukfU2jQK+aG715XaTG4vE
IFKVdBwXlX9wvemVGXkkxzJ6c5wcEleVkh+WuIRAdvgAQUrMwr/hW5JFGu8q9sFk
kZXanzv9daOFbbnEwpmExz+2hvGFA8REu2dRAFgKMuC1rn3RM6pyKuO1jKOWTmSc
HYKqZI3+FrtDykXfjZKIg09s4ctM9wPTpbm6LNV7ubqJZUYpjX0NMVzupGGfOr5Q
XwPlvous5Wu5Yn/LVpSevFa1N1NPxnGs8vbuPphj03lP79sWaUhLjz9o3oPYl3NL
JV5AniskvNNGQtohFjXG3eIbMH0NbjcVijYLPZqtAuaBsh6TSTjElzC9npvp7y3I
D+9EMcUQCyf/+GjGEoDxkyUGv0TmmNC4q7CiUx4Qarqbkp7I0kRLNorenfxLA9/R
w94YyoLA3Tkm1/2zSILutTw8dk2DwjWt9S/D45h8XjSip42/drd/lBImbJmrk8uI
9ExDSmaOM4yiyz5UbMF+BRZ3hfeiegX0iof4vBC59Ckz5cXHgMgC8DCgzTxxX1b7
bsCy2Ty7Pz/wULUncMBR9NZHFnLgE7XV64+aqWZ9SMISxldtUSaWEEjtRxsZY+VS
wmVT9N1x5D2EhzLIyeOlHYMm5QKtI/NxVrtuoDc4sYF4MTKtmLjV4lT6lvOSU4Xm
nGmBsoo0leONy1N4WY7ef4BEVTAC2CPvtmitnGRnmGhQmDvXCV2XQPVjN7ik3evD
69Tfh866rNQETZR8t1RCR7aNqLiZ64E1FttBi11FTvEjL/dNkmbzYWKuh53+yZw0
zKvIiQ5qqLGHpm25AIVe6A0WKAMQhKYMVCmy0Gxbk57cxMHqoHq+3c3diNy7SqsI
p3JlEhOdpLWdWlQ7l08NlAGSaLTZpiSn/jhFTpebininoIbRn+B7joupbRS3mclJ
FtEATcLYi6oAchJDCG+nutzaCaeTBQkFGBnitCjj5bB0zGTsiBejpTJpQFmr13Uw
MeLMSTAhbuDI/WXuXQYqomIQDCl6G0ngBARf4VmQPq4+/V2F9F60wWoak7mIppDA
ZklxHTw2XkT7mCHH8u8LVXb6xSqdzng+Xq8vD1a3aR6WrAPU/M0MfY+zHRsR/F6V
DV0pmrD2omVXBS3nH/F/ZYozI1Map9o8cEs/HKSIHhLOhPLPpsECdiNLNRVA39tT
MlJ/bTPPh3D+PMzrIX4g/QsSzPWU28YojT3J6yyMISF1juzeChAYlZmYspJw/Cnb
4QiOIaNbJDjZEMc56f05e69SXf8qVYaS4eGVaXBo60gwdAyJS0lrmtawVO6Ptul8
oFUqstqKe9tIOyDNWgC564THUTbX52PZ7kpv9H39Lnnl16XGERxGiMkgvrZZdkEq
mtxjX+GC9PLxCJNfRfQwa2YO4wnmJ8Abe2TlVYYgK4nY2HXBvraND1MFkKXBphK2
wGGOF34XSJBEbF36pTjhWYBorqaonigT9dNCc8mXpajAkoxHrcrxiENc3NvJsNa0
63D5Rb5mkEeOw0nFo1xDwJETx0i0iKTnDnQJZvO06ywsBcqfqDHtn1zeWm+P0X03
BkV6hSRbGPtLJKjyXpCMnDLDmR+E6XUxlhuooiADYGtGL9yB0xSiakU5kxxMp3l1
EXBpaauxcZpedhJoWzjsmZxwdXgiAMoqMhwLsXCOqidJtMRFKEa9zgmLle9zrpnS
lT2eXOMPT2N35OkJJ0kgYH2H5GfFP6PrbjhuuT/3aVic0+t0wWyNbGLp5BebzrRf
+xq31LzPEUK2EwP1FJS5KaZWFTnR+2M0nmXPGJ8jckaut4YlYfnYDped0bE2AfEz
eJGviEpPYkXnyf7mziamW3abgnqQS3fJdkLuk7KT12ybtLXAamD8JYBg0Ohvfppr
r2SQlF18mo/mlrPoLFxmJS7VzGwHnV/7Ocq0j2CMUZROvFS784SixmQN1sAJYpzi
af8mIXr/MSM+0FG/j1LvQ4LGry0tLX9BQqMDJOKZ759k+vmfaccGnixjYENGJa8c
5DSJOCVal4GigU8nKah962tv2xzVEgtGanlveBN8CDS6mHP6R28u2ISDnuuRLRif
0CqeqKPZP+fx697XsT+58D3iwcjlmcDrTpaWKPCYymda6NkT2gQX8EoglAX4x790
FuxAhFa2aM4jdvtVpQ7VMzpuTIilkSg1iBkVbGlJzpOyXTTq7yA3sMXy70aEQAda
CgWMrl3kYiOe7okKKAq/XHrj7dDsfFSV3Y+0THLUBnl+CwygEedpi2U3pmj+ApM+
WeqkphTEPpHujREr3sSY//ZzV40P2lKoRrhSXHStP14BZKHwAfCqgPW1k6+stiwi
kAiPnd11e6mry60tjcc/2OLsIcviXKu8eOSKDlDKhI/Ie/af+7pd3vPV6ytc4Lk+
6Lx21tUXOfJkST7w8APTGoyvJtQHyXQfrNTTu2692S2mIdKfNzbn8TNJWcrzFAdY
7vHb1h27WoCwYCJKPLprhHcWNZoB9ZEmQWEbIsz2p3ngbZKM8WIT7+ICgpVLe4DD
L9PyQZ8lRLzkxnXgrGejXSkzvEcORLLNgTfb5NPYTE1uT82tHYg9cPxGt+wnsBOQ
pw0G6C2N0zjs04eY4LUsmjdzdS+qVWDLPG4xYiOnzVgMu089B8ui9PeJ3WdN8ztj
IvmGmH92GzrRMoRcJi/3wNL+LfhA7iiKUhB19dquxRHzAqjVmY31LxhFVgI5mSWv
XTTNmCeVnGiWGfWYGAn2Pf8dWNJyaxBewjcFD1s2PCcYWbrKyqwR2eiyd9BhqIaB
jT2PoXq2V07E1K6qBojAdFck5j36BnFJ+hG0nTgLUqVxYnr5E+XbME6smwhMJwsg
UZPM9dRIKb04zW6q1/bsnjtsOuY02lFxUB9UbxbahDY8VmMY9BH9ly4NTXo4kqys
08PyfdGnUQtotfgpjXMuyUsDh36+PgNzAWGzwEAEF8HNjDkjDZlC0s0pANPXQK5Y
ay04R1N9B4SIFFylBU9H1/YM8mNJgJLq628UXMw9TTlLaC+4j8Xp+ZnNJVHMhXnw
7LWF3+YFo7bBRaVLtMXkvDTFjaqYQXws3ZHTVrYtTWbSOEQaXlthJDm0AL/PoYiS
d1KySzKuw1SdxjIU5aWM8Lin9imgaT0VuGhY1/Vw2UPMdneL7IvibSNqs2DBkF+M
xc26XQGcSed21MLfY9sm2GIYtQmntBLwpnloqQIe+K03pRSLrMjpyYhJ+IxK3X9Z
t8snNrusNjKzz+jDIUoaJaQ8q8lBDlLOhhwwLI2tyqNuUcwEgu962MkXuQFUc/S4
EA1tIkz5wmFDE++K3rnolUMbESH5WZuHWmmPAk4tsNxK144GpkolAY9SepN9qtIn
pZqAAKnhs7ufxQ3WT+4FwD8If1WNmbnO2zIC2h3NMG4zIubeBAwYgjssjv2Y1jfJ
bwN0PNjMfnyUm5zsK2NqQKI0vGelHurlXD+e14JpnGHvMFQi4GxPLfEamMoSfBaX
X7QUuRk2/aux3Qfc/RgJvueVojgnUMe7Rfnr1mFsoClI2PZQBUqATAo9VmFfelQc
YdJhpphnQJQZfAgGr7/2fCDRVpN9yt8w5ck+UBHehV63V6j6N6tH4IH+1usIVuVV
zsoPzV7W7ThM8pib9MdJLSIc/921cVscM3pF+m410erla8XETgK/eX5ZfAQ+6EUS
ZBxT+dm69n4aZ9sEv5n30o7fteHgDKIEGUwAuiNmdEd5Cxdqz667XZ0WiMDKTsWn
ydN/+/SpJpsFctt1c1cPrAkt5lGcl3EcLKg1pfMy9PlkXnMKf/DWOW8Dkk/G1HpW
mofN0kwQWOh+KeO98jnIb9VP/8ipwgD8e9DDPaeRnZXq3HOfG/KjCMkYPYxBsqZQ
pFvP41u5+Dg6JBtkrhBbZXS9ngJez1MCaDltF3saMI+0ZTtv3vKzMmzEZZ4c3r1o
Ymei/rHw+d8g2kwzofX5O8zh7prg7h7V02FX73lr5FP4vKRtoBzbDLPx2iW2Sc42
NHyuRug6i5wa98XrY6bAOAaqUvkfKEExEC7rHznW6tx38IBiV5tf1IDOxzeHC9xC
hyi865RSQv8IbuPYKLJXOKiYFQXYof2VMQxD7hewLdF0ZfqAlu3feWnDM//7yHzq
rXNYvp9p8BdmZgxMldo5VljpzpneZ59HU1T6G9Vccb2OFAcWeb3Bc4sa5HrrqlFT
z9eAFpCQrC8IV7HR5F6gSVd5d7Oktac6p6mVPjRPYeMnLu8EdfGO8hCnLyDnbHgv
AYKc5gB9lyA25nDpwtmzr26bueyCFH2jlLVTHvjdzW76qzTcF4/jE9XKIgTmoadh
5G2/nGLtpmyQZxzNEq7yaquJFBDulbNlkv4GNUEh9ENuo84yNDWzjTvb1ROoZ4V/
/X01p9PaQgd5UQ++BxE68jFRWqMXN1ATPfGeXAgkZzmWX/8S+PeoNDwCjGh3j76j
0fJ3C8sghAxVTWoUODRfmDKy6bGG8JjfIkQCr6RBd9tXDFXUYP6ZKVOHFzwK652C
SlnLYb7RI/vYoJ/y4DKq46QBkQ7/xGu56ZT8NoE+J02t/UQDIAHl8IUPSjNssm2G
AvwnqePv6YQajK6F3/mxPUBcSURFTaEMVsmd1KKiD+rFX7RKskvV45bqcoBP5PF/
tu2Xauy1fZUFJnq0kcw10uSehMkYQVJ8EoHIFJyNjxejlwSfvGNnruDvBHc7YMzt
fV/zJFXsk7IXwHPzAdubEXUqpiY3QramBCh4d8BWa9G0ZCcbmyojtNcnpXR0iH6G
KCUcAUJG0HoevmSAvcQ0olWogFGNfHgiFEHj1Q41UxLK62WLxlu4TkbbXcrhfsX3
Xn0kCvGG3BVRZyz6s57fF+6zsLoboKkb8nClxJ0HBHORtm6fSB0p71mRUbda/fum
xDKaAOCPiZPUKnFErq8pwZUGSymDDKviQvbbq0Xpo5JfXhT9SUvM2oEuzBR9OQdB
qvK+uo/IGV/kFg6Ti7+6YMJdflQFujhrqbw2IJ97LF3q2MuGoaLeCI6nwzJpBU5W
hZr4XYyixUjHKStDCSY0f9zyCkfEvDYltiM5wR6V0WxXY2ZNoBs23ppbf1OORJnO
CDJNqE48LqIDxoU3CB67Th4Cm7a6OG1QxgWoUtfBHr/QYmHIraia6zl9+nEKbmJE
c6l794kFrTkvL4NEVWKJ86wNOGZWRCiUhSKwlqxeYIwl9neyJyJTnbWtl2dUtvKv
wbHkwKJFafQqZCRBLszDVYs6HMS9WxmQ0Un/YgcoR5KgSnoJ4RwO8rJftsqPPMrL
XHuH24+Ib/8VWZtW+IjaOwb8zdhW9AmgmzZanaYLFjKsgvwCgdNWy4Fbvuydtoh6
EZT9hMepRr01sJb1txIFnMSJJmaucRELIWkCF0gWeCUcBnojoYVrAYtVEHsh/OhG
OLi/IHEPt6LjFDNhd8nUuLVr5LcRR0mWumleYwbUiMrSeOi2jfw6oxzfrhBlzTNb
lsShwt/PcgeOGwEnO3Jj6PP7AWYX2X/htZN16SqKhgbbGZ7Yf2vjo/suwl5nEM16
We0H4uyM/0gY6qnGfNDJWIkqfcwYa6cgtndKniMTuJJdmF1+BTMODEM2eSOPx4rw
QPvTjo024gML6kbky0K3IQG8OCvkuoD6BYcFc4MYm7iYD75VhqrFCuDIWfKx69+l
NbXpAPo1bbxNqniYGLfxGicoLL5/hL/TqBExAFHaLXPufl8VTz3U0hN4Gn5TUbVN
VdRCuRQxW5+wfqULYDlaTljhMsk7IcGZj9m08kG2sS9chPpkGXYCeml+R5ndKGRB
8FFzxbd+dWNot3xPhiEvZnNsy4iirZH3YILm0STwyvwlAVdY1q1sz1YFcJsP+X2A
SneDs+xZUKRx8gr0HsXiARyjVsvZMxQrmHclG9vSDsLI5Y+4yiU3WnPosMH+4XUV
RDYLWIlI1TIq55KIv74JGUMRfIBwGXOzfyHuJUosQbd+KKKD/zU0SZLLk03+sZ5U
Olxw0G8TlX2F++r/gsJRp/+osDBAIK5iP5TCNbXu/Mt6SpT0MvseaGJ/hOQ4cQdE
HTAhZjyW7TzPtdK4YT3yPv0jUvA76QSXSoO7q4s8Rrnqzk0HFVCoIsIw5yr0spaa
u5csXjo8JWyvsAfbHvXk8IX3b1+67/JtSfWgZDU/27JRXidCC9Z9V2zxFDeMJQU8
hRwn68OEkqh44Ai9SHAo75DZowqeZ6qFP859j83EVTlP02ZcdEiZpRUVU1xWgF/c
LXmNntKukBzKUkRoDrdDvgobIQeFILM9Lkmadp7EmWf79FjE/Nut03MAqvZVlBp2
v1fVSSNM49gplfFU7ghSG0NyOFx74K1VrpBAp5gMB1u/EAhI1RNSeaC4RKrWsfH1
brWGWELwazo/3Tw5FOnJo45iU3Ok2TN1ENTq7zskgxE/72nCa/o+raLSG6PYx5gV
4RvmbyeNsVwGs1XWRMJL5/C+V1a9aoUHwrwthJqflRtB+N17EaKJS4Vsv38rmKXg
pzp/bN0qW859YEXR5hzdAIUy70KBBf2/Mc0yA+V9/k2C0eHyMLqQO8Ldv6ERMz0J
SBklgXeH6lxCPzbGH/9GR5VOG13yJIsw4uANvvVXqiOB9FvKZsAny2db8m/NefUd
HouLHp9Y4lCLtQ6Q938fKvDfIB3oype2TaRgesij+voRGa+R83/Qw4NfmWtHzuxP
f242mShR4TWwTkz1h/jvQqQpyRye/QCcV0YIASYLURvp90DeY7c3Ni3uEwwXo6ZW
ORZjU3OUfQKpB4QGM4Wzs/NwiCO4dAKmAGy804J9+nGsM4OdnaRsZxiMTdbgNM4A
1Z4ICTgtwiDx8oK8zXrpwrRfXfO5me7eLukqEaCKct6ymFi01qO/wGu2bnQOdCRp
ArsLZCjD5fXwSABHsRiapV24UubYZvJO5at3fZqbqUoDVKB6yz2HSm+gbrOWv10k
fYx68I6o0CUYe6NKvVo6M272aQ/N9MHKWrVAFv+ngoIqLn06QqEt/+CirH0RWLm1
HvFlAUFF1Ba2qeWhlQuIDnRXJTp+78u1Pd6LS0sq+DDKpFbk6ohFT6+htNHvwsgV
nn+wOI+ANRU/p8g32I1vMoydX6nYqcy1VuFIJMQRkCDsG0OerNDnQ4IQWjSZxxwn
xp8kAEim8rW1C6cTpc4T2R4nGsH0i7zHtC/lSAwN7h9kC5v5xwsY38zoKA2Z9Ijq
hgJLcV8dWeqCnutLMPND+xwZFH7xvpJOibeo6bDUAMAvrn5Oj6jtqE15GTamceX+
n8ndYyBovBpP9Hy8O5IOd9nhoBE74wORr8PY9p0ZW5hqu3f/AbEPsMNG1kzloSQt
dmB1RO8k9zN8zaFU2dxCClYko6k6yroA6iP1Lj67dJtrLQc94sB88ZLXwkzqbYj/
2hncJBzZLcsCc1uvuPA6BTay7N76ccWyxZskg6S0UOmrqxnpk0TcRyd1iAoTeSS0
WtYlDmeQZv2vYWnPzrimrysa17AV3W0AtHm2U9rZUGevfg6+pujfqkXdLvM3O5Z9
XL91LYaO6JWS88YAycUfTYLKuLqMMdu93v33m6IGKz74N4+Z5UlgzwYvLrxX7Ikl
htxckKMm5Nh+hTckg1kwcGaISKez9MetI6IyPzr2ThPNUS5kmNeE30FhAX8Yag+o
SCXH2EpNQK7ArCH8Xe4ceCvr9zhxBhyuvZSWGx4t0eTW2O96VOpdn/uUTu/uyfwe
Ql1yDrAha97KszpeN/1Ge99M8RnHUvfEPG1f8Qa4QvN4k494tCrT8Lf3kWjhwrcv
R8m+Tfo+puek2qUOwEbX4kK1mfRXdrOTPT7+qjdF3uDmyXUXvYpEHPRCizJyrUp5
2I2ExDw2rJLTmwetidBXj44nXYiHfK/D/Dsc+e/lx23Xs07pKV3uV6Tw1KTq5AcN
pY2dzoAXpBvLJkcOjW8ov+o8ifpap+aEIxhQimLD47jHr+FkfZfIyeessZ3qYX4u
7NxJ3aUf4s2HlXvwXb13P8nEsaTF3GV8TnC+tntUvhraEGu20OuKvm3NTP+pXqUu
e5lLpcZWuLHleHLjhOr0PNOBHuTVHVkmqMorUwBHximLGFqaPVPnPloC0hu4stQ9
9oSsQz/ta5gvynsIzqEEPpe3iZt/cNmurqT6LDaDK9OOZCuUL2i1oK97RPtM4ryC
D/z924FsphI+kx0BhnALq7x1YHIJEKWgm5p6j31gaW+g+oUSeXJ/ShDvSnKId6xw
nJOhueAunWElQ7FML0DkKG8baq+5g/7U0troILy/F1bWFG4GYAUAd26i7anWd/sz
BGk6f0qRNEuU2NlGGCsM2A8YwvMFzfnqkEm0XccAkUyh0Ljl+uGdoXc481Oi1JGz
GWEo+sxbM/2h84WauBul9qTGddBZyIjppBiCirSvGmrwuoxo3l4jH1TnQYGY5s1W
TA4Z0XT9iNkfmPLGymOOg95mdlje306xwldicOVM2+uCbAmXPl9aVPPwtta6y8U7
P28UT999oIqZtPjh+/LQLwkh0122vwTF5/s59A5bMXANNqm6VWgrB4ATxJtv/HjA
38rbUJrGgejIxp4WJOgzUU60BKGUjW/9enJoX2UF1ZJDzl1+5ZD+YwR0Yw0A/qin
f/4IGpj9VieFk84zTK1GOcFgt5dajhHtpXGhw59Us61BICoz2r0FqLW9nbeV8W60
TNdu3DP7RjU0ghxgtC4Fz4OpBKTMq9474WSftNNHn08S9KV3kL9pvRthI/7QP5hk
yVtFvzldvNegcKnnrEFrByWaJplDyLQEQgV9Nf4iJaXWNAi0vf3cIecPAKe5hMKe
O1jazNG4vsnZazIPFzKYKftntWBNSvqSxX0swTBv3OsmMNHAMBLzPRjCt9FL0+es
ZuCxp5R2FMT38NI3x4Uvqm2qfilE+Ca3c+gBua/nEWVLk27mToHJlAlRviF9enAw
xQgfHmyAFqrr6oZUfXpAPctGZKTX6cseesjzmDoGvc69c1naPOvuXC7YqdvV38gB
IV2UocgdJR+aPgWEnpE2ukIP1yufKu+m26eFWin0aGBcn4uVGaKopm3DK/wqluy7
aXuiTBZqA5iun36kNT5OmN8Qd67PsmL5HIEpQ3rf12xPxVpf1uGLWYZ7+RjdEF0N
Uxvs5T1/Jhq/7cmzaS9QKiPsBv4A3mfN3LGfhBFD1TGSKJdpOojA+2TcU/f2uxHX
IMsEmh7/ntvPUrq3c7KpOPE8VAqdiydI+HF1WhBl/UanREFv9zv+G/fqanCC7E4d
yGgMmLugnWX9aFZU6SDe2bK6DmU6/aKBsUnRNDB3QGmOI6WSM+WsBUyK1EbrHNgd
DZM4lj+6kdDkpHaAFQhwZO1Dv6wmOrjnFmGTfdOvNfP0kehvMxy4SCYspKDKr+dc
rPYXnsGuLkUXkOoYMb29pK4H8x1QFdli9tTHte3CLuNcnLaqKg0VzC1wtAp4Mbpp
Omnt7XvCqxespjLaaZgV7TVmAYBJ4f9+z9o4wFwd1lTNY5ODSF2V5/l1bKNMb9eF
6IaZYtufzKWOUqsiE50220pMLDhD9AHstnH71yEWKW8c2zwTNfInc7XP0VcnWJ6h
ttJyI+mVO9DXirxTwjIpMubkSYp61TQzBPpnyjMHABImJTSWSpERmlH+GWl3VhFr
sYtb+Q6JQBMLnyEm7WAvnNFA2SjQJWAjECg4shEV6p2osb9hjeaE4tK2c/ILzFpj
CaBydnMuFaodGdejqXfHX/1C4fMyCIuayTL4jTpBGih6AYwNsRE/YGlF5/zWWZyq
i+Rq+P47ROUwE63lJEMsJ/CRN/pIESrFgPjYXlQ7g/nA2FVKnDK/vq2ryMxVsrp8
igykuYiyr4g5LjsBxfL2MFDoywGyTj/LLvuvqtneQm3uA8+OdQ4Ed6f6AUYVwJ4a
BF5pQEjbmmPzU+EQye60aES/X0b3KlcgHHiF1jdaLOCIn+iyo3l9btbBgS2qjZeU
2DcdFNrmpY0yUdenDDyEUMGkvVWXFtgcKNveZ94iZfC/45LIz4fqFUJ4iDFUySTL
+lG0UGm7O7hRyYFHcmOpXn4cBYVls47Ao8ftaPonWqM5vb/jM55dbH/y3y3g9X1i
4tMpNmsBEWOgewiyfdAXJhSoXbxkZV1X5vDWBDid1mIbDxbulMhfmqkR4TJDqJ0n
a6q+Z421ut1TPJ+6T0kNQtSp7FFBZFhZz0CI3JFXWF+sP2hiFRQyUAZlyiU/N95S
oXin51xdfHwqj3GixmAiS4IlOTWOcc+vZ5IUbcodIJ8/RLt5r1FfWCdOm+qECClk
H3bSVmd50W4yO6ueGBJfl989OJitrs06jObwL50fXiYSDfy4qlN5t2js3bkfLAzK
kpU5G33Pp5Ex8oP5weGu1ta/P28uog65qM84jrYhoIJx3xIG9kSnnNFx2UMg51n2
nW4UIMuDcLKiMkf+eSmVRX9/HAZFGhW2K4PV2Dv2cR9zxynGsI9k82lmBqz6vVRh
+VHSR5QUtFULgxtQXT/2DcJqwUQshDIgMoT+6sNZtJD3Kxm3khMAAKKmBc+rigTv
Qim+lh3Zjzcj5WutpMc7p8Rhow0y+NpkN9ydD2VzVJOXixz2A1/vxCcBMSGmoYvL
3g9ZPRAvMXOtfXq+7ypwY2NkaNE4N2fGIhJ1YvD7wymbPS4tDB/xwA02VMVH+KJX
wpIyCDsFDT1dN+QjnvlN6kHzomoM7FCULW/rce1T/cciV8GLZuJwxUK1PKIU8cQK
aiZbRCngsaTaYXKZ/hBUPJN42FDP2fFLdcsaY9bNoWrK2+pewuTSKSoGKheveCzN
xIv3rQHjnoQ4sDaXt8VgF18+1G/ZsOa4M6j0FsGNGQWWjGh8J+mFTy49UfkZJvia
pZ2k/KuAsxhv3Hk//MqUQISQRl0uUEfxfE6Dt86hubVKQQPYkO4kuo18sANT8DwC
Ih8+5NLMF4AjjfWUwmxdnuVAqRvGRcoCn8AfyWivp/QlM0mwcs6w9fRqih3YCLVk
C3BWcdINcXwXLF846R3cDeOWfkw2fYwRYUBDx1ge6RGW9E7CEeZ8UU+eIKqe9Xu3
CKNUorkp5yj5KxYzJF9+CRp/n7rHB8LyvyNNGjNzl83cqQ3tRNfI4bL4w25UtXR1
mNx4Q82uaXv2JuGZzOScl05a0f3GboQF7DZCZza1ime0nIzreUFmyoljlnJ9lomW
cEWVTrApSLcxuIyWzsFV2NC6YK5KJNCObEAYaKymC2EVjQfr3fWEBSTsgYWskTnw
uFNEomlFzuM+Dt4p89N+APiIMfKP80pyg9i68/dhh0QPFEbT6zNpmXRXf0d2bQ5p
gkd1i7dWU9bx7ThpJ0LAHY0/avhTJTPqNKdEYRMRsZncfjNqfBXtKktyMPvn0yzG
IIQr1+e54feQIt+EE15NOtWhkOpPS62loill4WRjv29iJvpISvys5flFh/Rz9xhl
HgzbHdNmuQWyqA2Y5k9tgWYA5AwF6gBQpJ/f8qM43erm0YNYoM0kFT3zu/5cRrdJ
36JQOct4nvsB52om8mM97z7GgzbbTvcJoN6hFCvECfaJOZevhCRM1LRVoUrCC4zP
zv4QUoQwJWDu0PRLE+Nqg0+zHrkiw3tA36a8cJ+6+eFcPO0wIjpJXR7Av+ex+N2n
6YV95pPMGrHTCenNMVI9s6pJAgG/GaJXNygL3yxYhxIoZrOUnkitSN2dHBidRpW/
Q4AroH6Mx6TEonIzhPQVz/0hGzqrw2QHcgtanz7399TsIViudIP+KZG5byMOqSnu
sCW4unFl8dliimX9g9kxSg==
//pragma protect end_data_block
//pragma protect digest_block
cE5dwEosKoERD8iGUMpLnFV9qtU=
//pragma protect end_digest_block
//pragma protect end_protected
