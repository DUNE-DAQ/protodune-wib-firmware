// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HpgoqCqeQfQdLF9Lo8yZVKnsmVa6DZCxrrO9/ViqMo3eBj/tbSMoEWowEuAIGotD
4RqPVd+I/tDoqyaU6uR1JV2CEKtn7p0ON0juLipflrKJkN6BiHUkkiuZP+2joo9m
z1uvqtgJ5ea/pGaDtXGRQxwd3a92EoODRNICxIWfMuY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12176)
AnQEwTDPTwa+pZiYNji7zGZ8oUnZDeyZZkp0gwacBJdceL5Qg0j8txgmBJdjIpwk
S4Qz51XT2ucBYZi292CH0hdd04VbhZJeAzjsBHNVrr276/RNp+1xKx8gOE1hJI96
wTAIjvXvcZI8+RRdVyVwuOQda7iNiQcNPbKNMkIacWMbEPcpthh5YXVC89iKITfB
yga2jzpBuenuIIf210lh0lrIjo9xze/9mDiuQ4KOVgyWfRVHfG8m85mjkRrziJ4u
DsTT/zJgWCrWz4cvioM0P1XSHqDOystXKfoiFcAsCJlCJGy0XUkTMS26fII+680o
DXl7yDn5ar+CXb25DkdcXdNUAWfco9FdW3yyrl2HXLnKCMMX2EFZ+Wy7QTlkHH2D
yNXgIneMLxriD8W4foPtg+npRpyk/vSK46PdGbDUHhxU0OUYd/u37l5oTaY7RFAP
tBA/8FAI5fkTMArTazZXSKJqgDrA6T9SjEuBgf3PDw1PZSVgMTmp5CcozCmMsOnA
bg01/J20tFUcBN+SwFBXOX19JB/2+UbG9fgT02hhSO3wiXO3b7EuB9i5+Wll6QWA
WwhkkLbUrRecYxa8mNq9cLwU8zOcT92FCBCz8dTMzsN1Im/zII/Fv9IED5ygDRNG
zMnYdSwsd3VmivL88tPFGZwW/wyXWjuyK+CQreU7nrHZPuwUbGxEtnl0G8KfxL/e
L/Rp/0PjnN2+BoUuG7I4xoE0/TuF1FWgjPKfJkOLJ8ROkoLvDYgDOlBxefvr33SE
89tnD5gJ7McErL3h2Gtrxlyvr99OCNo39exSM8+U2cA2i4nXk15ydCstW1VHWn5Y
H8riJ4UCwwuY4PFKzZKO+AjCcBHSzhJkJ1ZnxDKh+XxIVayFI2sVEeRYyPe1h0fK
32kRtDjXbduZoFwtdnAQx2BOhtcK4YSO6SLLVa/X23YwgIg97ONmtXYr4y20CAaA
/604rYhqtXgwW2uwinE0+5zmhms3+ctsKFdPzdgybejWpbZ70XWsw3Pxl08nZJ7U
hu70vIFUqUvcaYlHcny3bU9aF931sgpAU83V91TMMHeYx8uLfCSVeEkkckxQ2Mtw
F8Ab6+omEn0FfGNByewLYJ26kHpEd9sNI8CeTqKTJRDaPypSHi7Gf4qhqrIlJ1iJ
PGmRJTxi22umhjm+4A+pOog3vLifWAhBUfM7LHgJXuLSk/7EKJ9kfxVEe34q6Nbh
PJcwv2dxkSOahvU6iTcs0V3jgoziWsG/DPA7KaVG0rok+vot/XnC/nIJIjnxTCVz
7Drv+Z33BfQ8mcSOY+Hx7nrrRQQmtdgsCpswj01Y1pUqe19HfYV66SXr/Iim0l9j
ADHUiTxG/V2BPu9r9/vbc99gQaXbJekJnk9S/ZDMcBvCua+VcLH973/CTf3C71OC
jEcbe0jZH6nRvRN/u0weweJ62timFIksO+vEHwb8u9SjeJl7hYmm97/ofa7tw2s8
AwMEqexbycgCjGtAdlJ57F6kPSUzHjGt1YzNras4WxaEq/3812HBIkswys2D530e
b2ajaKCeRiorGr/VcH45er3U1RjvZW/dFnuFUvS91gwSP1mmyEqEv/OaM0SeQwWt
dhCm15u4sHA8vLDS3L/XbAgXk+oZluwiYcumuDFBS5kqpp3tz81OMoKMKiLTlRna
ps1ERUk1Dz74cN0q60MHmYRGwVzdK++PaDlPVerX6hj+/bHYB38X3RkRmMY1sTVZ
+JJAH7ekqNFjGQ92hbHB5ads7Rm+KE6pIktA6WL/WS0z4+MgurZlBGkH1QebEr8c
Zzj4d8fftDtrtoZnQZnfftBQGm0IZkOfwQ7aA1nEFugNF3pkixmyn7wJBZKCLibF
WTGag7QvlAH7g2qA6M3+/fLJZLYl2fIfxha1VEmJGplSBRinoyAVNVq5Z/JkHRaA
w3HmcV/quVsPOUaBY6GkU5+EksUw6MYKJMdDv6CJ09gAjRDroxQtD9RLPBadadkc
jkYs0Loc9t7ftcfReFJ/x9cptHEwzXJtUWrN3/BcoaKrUchDqIyuRwIniKOg/Xhd
oyZ/Bjais+3aLug5EcvLeOyGy4iZt9vgFsbHEo7ZNV8RWabypgIIeZxJ2MFhugbh
U2OlaYiKGNKNOaqwXDLyWlGtmE0FmFsl63tVPL2qkw/YjeGV12RT8pVRl4sE6lJd
aMHw4CaniKI9SwUde0GHZJUoBti1NBfx+7J/g3a2KfbYRGYjrD/29DJM4HdBsDDc
r2xp/caYrq/vfQMXIByQaFj4eIRlo5T00wBNjtkxaQirDtT0vGM1mUsnScQpdd8Y
EIicTjgY5p+Vf4TI6jOW0t9Cal/HKgL0cZFv6bI+pAvr3T68yJiZ28STtmvOrhvM
zx3y8DSGepZOTyZYVbxv0hTKnsVuejKhHgpkBimt4Gr5QXAQWg96x0VWVwJu6ihz
0Nze2CZYIYaJOyoHY2uRupSEI7pMz4hCJ+xAz+3U6ub/PL21qgRcIGXEtJJTl7o5
087lHZdnRZXBmXEn02cjvQwoSZ4Iu3RGEkR4yY8aN2UqS9K+cKGguxnBO50u6bcq
ROIi73kjtzKrtCU2O9BdqU4BIk2hNbkF/p+0A28drMlFF4iZTaXERhGPuw6+sXMO
9HA/a28Gcgu0QcJk4YW5l1jF0UI5lz+9kSOgYZUfr7W0YzOMyaDvI/OHn+DXbN24
zNLRqV/GAwVhc181V9qC0ZlPQzDHBWrCZfOd/ZetIgvZqs0cOusfBGbMb6nCoNmS
vnw47Y0rjlrddSx73rBKgDxU7bobxZG3XXQtgVrcy9vahIJslwgZoz7k0Eq9A64F
WC9H/luJmuh39MGASA4f6wyf05DiG/xGnMBCdBx3iTYMewgpodIiY4QyBwE5pzOU
Ho1Fw1UQMz/K9EvtK7Ed1ggcTQU/F9WFaLpK42EA4gqQQcm9gSk6ihKwI5xIILAZ
N6JBzJ3mhwbE8M+pVlH8+qd0ub3vsQRVZwoEjjk6vndH4vGBPoj3wTOM4OaxupQA
jbZuTllHwAQg5EUkO6EnfeHmgp8FB1sUG+b5IxrlqVad6i++CTuiMBZSoUxJNEhy
DiWdlJNdRvga5zJD4QOVUgJtDIAq2LBb8NB4izC9+IbOkeT4nN4aDDC8fcNi1Oly
pl0NYIzdqZJLCsqVWHRkkr6oSByHnkKY1P9HPqoY6++yBfqCGdpVPTgUxD2N+z6E
x9QR9Z12DINyEOPhAUTJ5uoxXaWuhGID7gKaGEY/rNLQgDP8xq5Xh5HQ1WR0FYMH
vmzF4r6bBbO2Y2mgxbnB6pj07a3+xaaObTtAHU7weS40kcQv5Yvcy5y2aQnvyiGd
skJBzOoCWL03gFneA5Py9+mhHN8sruBzbCX1ugxivdW9IMbg8ju+hJIilIwPZmGR
ZalFM/GSLtMQDLgIjKcYc4gdHzH8YOXWZrEKnSUbdvCUVQ5EI5IFnlNxEjXssYdk
V4L43kkwnw5Bhv9Yl4ob9oScEpy77l99456MGYMrWZBq0aj40lTV90g2wRyeh7uP
tgRZRj6KKB2F884uO80fJ4uW+NLC4R2Ud0OWGaX5ONk1XfIhLwJxJxZYUhMMF0S6
DpzuSNrGUd2LqvI3Mzzyh+8oncz2d2bue9v7dk4vb2R5V8v5kZmwb5KNAn2C/sCe
TA6zOqClZ8s3pe1Mmqw7iPpHF0GeuwESuTo4bY7L5lMhrCm2wgfMkVcnUbmuMIiI
rQSp7RtsI5GH49bxjlQ5ORTiOCuohbSLR43izqxQU1JUFkuLTTAjbJ0DLBny5kfO
cJBb4YzJ0iASp10lzQGUSSwd6ltO5rQ1H5cXl7fkh3LNwnOsQM1ECDzVLAWJr+O2
VfqPtXlWbkwh6CGRfTy8SHyZZxyEUaf8sy1ZZov7uN0lUla9HFFejlK7JlzUVtEo
+tv29jJsNiNHkfHJv6J9oNbgFF+OSK10wA36QXa/8wDimsepBFhceTIIMetFQ2sS
dBmNBvbay2mSa4jh+aUhaL7ufLEny3N5ySVNN7FBB5wx8JGtFMprlu0+t526HBxU
FWwSHaCdDXAr+7JELNXJKWq2LFPv+ehWM/GUVdRWVoyUqDkasm9yHqn+exSEAfQ7
2FnAoFUZS2OFxWeBWRxomzdKtsS24MDs0IVQkvvc/d53ZOYGK10OpPS/7DjMd5p8
f1EkJC0ZiTwoSxPDvP80wUTYPvDFCFWXK51vmLQrfgFtqpGlqBNSaXke7atKbruO
Ed0oYbmJFrnMF+ZN3QVA2LnjlVuwJSy0HVATOdgrB4MAEkxNnUhYVTprLoTapsOe
+8EQAxa+rK3jDQCyeuXMefg9PCxFHq15En9xLyZgRHjvWI/sEDD6xXj7vUwVK4DR
OelDB97dawgAzQG4v5HyTphoyUSeMpiuRtCx+32MDKcW8sgi4vrHTaAjaaNns++v
qIaV20omvphBSXbs1o4vtzz/lPIwj1AKkjodYftWNDD4ykEPEvLu+9coSFoCW3Na
mxGc1Y3n/p831vtpfWuMTep2gcOSJ0y+OYEaUWBv0Yb2FPspRzRgGzDqZ30np7fj
g62B4rxxh633iAFoV+v5lpx6S7Z0SKoED9Op4Id3KJrZQLq50Hum5TCIwhuDnCAU
TKfbCkY67A6LTSozpioZbbliVeHxVuNXIOMmkLpyp5nhWLdIaAqLYaC9ZwEuwUZR
aKgTIFzUUeqAqVSu62l4O3Z1Km6awB1DPcvn2cUrwhWxY/tGrkg9+QnDJMO6nCdt
ocqR6yDwFXEH+9V6iOxl17FimIKGGQaIpPy9J6oXyAJBSSDaOjJS2FovOZmBjRXQ
YfMdqrj4fz6XQGOtxoSh85XrZel+H7JmuOCT5NjHIqkZ8f5O8R3r/5j1NWnKpqW5
IiMsKhrh41LUmZD4yZgxLVGJbYDl6s/AMXWkNIvSAaoplh1PzXZPEmQXLO9EcaVn
Jo/AM19ZFYoBWTVZEGoJQTIINN0xr9B6+1rEL7Qrf3V+sTrw9zDUhgGWyCm0vm8E
sfblUs5+/pxoEpfAPvt7FkqSXSU0uF4oLvNf4Aj6Nw/+LAqEflkzLBAjkQvtWik5
c5WgPJC9XUfZTQ2/5vLGZiAmLxA4ebrff5CFm277AkMruTGp9mGcTns06NItr2Qj
rCXCDmPyGSL6jNWtPnUB54Ro4zmw5wBRmVOIyhEcn6GmHUOYY6THJDlHULjvRmVm
QZkVc83sPkQc4iHEpAkugt7h8U4xS9HYliFwdNPIOiff6RVk8G/744EWVOSUaN3e
3T/owG+5e8a4va8CqPEDC4MeHZEA7Re1YHtkfoNU2ssA8jMwWXEYVEJgSHQV91dG
4wBlgK7mmH17EZyJIBzbMkUE8ZhTHjz3eqtI+q4beWc5zoidTqfb6tosSStw+DBQ
vgQSeY4r15XwkSl0v8cw/diHXdM/y9BZPuK5SYJLeDsFAP9yGdaiOuki1PWFGTC8
kgvAmvOAoS3Fw5CT272CxDSMj6OBwp/CL7hkluYyeoS7cbgqISJUClCUivCafY12
kBXQY3bQkgaPKOIMnTM4J9oz3LpKSnDXmJ1oslsk+OHAJFdrfRgxTR+OmO62fwLf
Xfj9VbJLV47CazlPa3kK3aTxifHzT7xfAWTTZ+UnP9vRvzl18jbz+RMWPk74h+LK
kScovnhRvzZIyEZPmKDLCLP/mLblymhIUTEoGxJF2U96TqFqslOABWjBOZUR5jMT
bb0bZkZj9KPRMmsNbfGiGJ7M8ck2gngCG5FVUDFzvNCtGS1e9c3SpJVHo40sTNRX
a6ZBLYpN1aC5uBPsFD7XCXMEV5dremqhWE0IMFEE08YGzJhUCHwPqGmYpkoHjG9M
WFSryJKjsanFFW141UliCLufaTbz+z78tA4SorxaevnbD+Egq85C087MQBKL1U4X
lnVrTTop0ee+ZE9KDuy9Bv3fhndHJTQaYAHshVbFcZPvrrD5miyLrD97BPpsUFqh
S6GpzXz/EcijB0Lam4QQNIgAHAZIKQP055FC7kzkUbkXsnjEG2AKXSkYAorNJQyd
VAJveaofrUOoIn+WB1hmiyoTkoVIYoVuPHUzruHbDOj5RCsmoRRi8Ccy2/XqJVrh
gyo9YG55jNimNR9xjJRW5cXzYZakfn5i/IoKAS1PNoqBZExLywV+rmwpf1ndZSA/
aVlTUoTQaPO6N6lNVVMOL3glQbiFY3d7BX3jrrLjH6rFuraWFOJ8aLSlR9ugOfcv
LyP1+v/RrS8E0TqAyZKdsmU7EepbK8QuTkymbg+jG7wvuWg+0wHXYjEW4TkR4nbU
QY8GjgY9cCvAn9ZRb/50akJgRoqu6CzWkGwzS+/qbRbXEAoSRymCcrgqVMTZMq4x
9P+XeOazvdjN3akyTqq7OIdKqTN1Oc6heOmrSkr3mT8ENJ3UzBp91i5uZwQoINm0
Oa46+wmG5MeglL3yk+zH20TpMLf9r6t0+aZyosYx8cS9p2iHmBu+qqPS6Afme+JW
IpHgUGdyaczktep1FjAagoneH9uIUtiUikHoK/4rg/2c3yzVjrE1IqZdGI5d97M3
p5so95D99OleptZIwfnrxeZmCOVxbyWdO26DY4sLrFA1aq+0yy0bVEXdmxJaJ+4l
J2l6T9I49mEILPu7DMYbRQna0syA4rzDzgaqXJwpn6G39olvwipq5ShmrsM+B85e
Ck5jQJY9W2by7X4Qldex79h/YN3dl/xZQSvs5bgfqI4B9rSKqPTIHeQneL1gLKvf
cXYvam0pn0D2GCwYiWgYUcs/cpVFlpPwg7o+RLbjpNSZ/U+u5tGck8NVhGyUQlQK
rZry4XAqs335AiOloSjJ6suvY34xIbm3h3jZu7ZmCLnv93g5M5vX0j+T4SROhAXr
aWs0YGstLYDe6YRIHiawlKf5Q+KDcjf9u1d9fWfh4dcNRJnkVcg2DshopjT3P7Kg
vEvNwTWKz49pK1uskpn5O9Uf/PrkgaCWmKT1UaxxHr5tVZAqlfEMWJ66j7DI0e2j
WWrbzs4hjg3f9AeYvvf/mOsquayULps6k+88Lt19BPjAfZ1oZr+hAc6z2Bp1sASX
1HYAGFyLJkHhYbdp9GtWBpuQnryiT1pFDsyH9kyCL+ZgUEIKnyhRQfedcLNGiPfe
etWZU8tAA1hHIGnvzu+Aot7X02kDBqv05puNzLqzBJveq9eR8dLPckhOi/vkC+9K
1sV1FCK1WdpMq2PIcmf3FQaCKFRSIMEHDtVZaaho6+cpjJw9TrBf2vcVxal6KuN1
7hASl+Q73vaV9aSzYychfCSClgJWSw3AEsgfpGiQ+6fx896zmkIyi9WPVACsRnzn
yNeGfv9DhyTCDiJFwBccSBPZ4XzeBDr8BKa0vJDyn2wAo5jFYSzLOrX+iNCWodH5
KOnYY6Ey6aRM/P3SPBFmRECcNltqKY4IGN8W739KnjpykVjY2+AgNi4Cfk/azinR
f6Qdh0Rjlu4BTjwZzisPdwhiZ00RhNT9kmIzgxfAe3MfXQ61OhbVaVk0yBRVQwyj
CJY/J7tu6YRnZl3RtCp/bK/xO2ZRhnQTI+bKVsvn5yCw5C9jngZEkbCU6x78VLba
ZISStlfZpRhwUozQT0TKekkUNiw1f1e8SNpqEIzl5HQXzplPKyA/PeL34pOIgzwd
PBUSji0zUpZ650RlHe4EYHRPiHJggD6sRF8DdWLJm+Bo05Vi/TyqsVja+U/v/XRl
6bYmpoXbOCg5Eko25OU1SITFs3SvZKP3vXqFWp9cyghNQriv1y8Q5OR+HP/t86YD
V5RoQsqjahk0wNf5LdC5xrZ0Q41eli++8OoBHYTOxZwkOR3vsfKXMgz93X6xIxIy
MMVafqk4z1TixjaEGznx9/ysocuWi5HQtSKql2C6Df2SDzD+IA2Igzk1ryrzarZl
tAyP7aabRygXnoczxtGBZbNhxKYNszY0R+QsPJPsg8Oraxf+AFKNK1bRCFsyMFgL
4ugPMAczuXTjyhbKm5I6i4Etwtp5UwtTzsuy3ui61fZuFeZ5J2niXhBmbvuGhUpA
78SjFdLouzDbwU1KKtnGKkGY3JB1IjPwk3UQ/raB/rGX+ncb+Xf61jzrkq3gk9ix
hLbzUBayjT7lDJMZA8oKd+FL5Tnq8kTpvw9W+h14SgFvw1XIJ4V6bAQgR9QVo1sg
Gog4W1GXYhaacrQWaAg4mpDYHKqPptKaFmCq+mz6FZHm65DQrn1h2bOVOdXTS4Hl
c6Joka5dqR66HpNGCCpT2i9+vNiLTykkGbVeClQMm7inkSwDCu9Hy5egwuu3MrMX
qqkn22ee961iqrPtyX0sUqBqXCe2GUlzbg+rg+evI5hOyadpx3UerzSv3lUrnRgU
fbFVs4IorvgKglPgR8QTR2IQpBiGqKpvCVnZs2/XyjH+mbnsXD4FC+OgT1NL3DAh
BO2ok9TasgtLaFKLE1VGP8WGdygiD3kv1JdLujGVbBZSVKBWQfYYKc4Qmh4oIUE0
tUlSs5WrjVUBJc0JX6Nlwt0XEYiRGG+eJRN/OVR7lOX2t9bnJ/Bg/mW5rCGcHYGO
aVUjJVEtSRuFe1VvaV+jRX5YQVayvEmV+5luTJRbwf23F4qDZwBzKSaiYDMAutvF
uVvauK3XYu89qORGgOvythkoQrfoc0lO71fKFip8GQJWvV2auKjkzUrsG796QetB
y6p2kkFLljmsbukK5yf+ZmPdN2R27yHeu1ppNZMVu4/5PSsdPDFcQWeoyUErHbmy
n5r72Uz1JVCfRNuwfuXSZAXQqzZOojI0XieUIbwrUTIrdoeeI8Fl1ygjriAC/2U3
mnZ0D2eLoqfIZiqPg2QtQSEiCPX5t7QPNGaydnMD5GWq5Mql2HEogK/G5dXAOThs
hBAIsohEt9574r8kPwY+aV1TNuIHjJVgt1qCrFoo1d1UcEivclPoUK3HJX7rbe3E
jkBIonu1issqyBcBZ81/+IUdo3f4hBSFSfNKe1UFCzlK+NSpsCYp0qUMt7OSOf7B
uEaZNPNwkgIwHzshQXXjT/fdFkpz/Qyo7k8upERPoN5G9kiTdjSq2Oi0NoB39Mqu
lS4EhbsgnHVS0aSKb3sA08bhRq2YfRveT4B29AUHGMGPWwVuK20g786x6wqBGUOH
x/eg+G0OXM6jFWpv+Fs2OCfUhpnvxMTE+ehDJ2maYdeGoktbc1q5dFYYDnH/Ofdg
JX7Oz5HzRML2RUy3ZWYZfe37kaaxTtZRKFRcrHxp9EzUioS4tD0KP+xMKjqOvJTA
wC/xYR+NbIcwPfUfeVRck4DZ2JDPXOsENyQz5K3Ufsmv8//vozgEImJVq2D9cw7S
D1IizojC9J4hGGWkXyUpTrPdXSnLtjkXSoVW3NbrSgF1ZBC/Vgt7DNroBNjNI3B1
AjAkAypHqEgJgHryiXYya4/sG2iLuaz8riQ7DepmrAFX476H7MNR6ZAVb6K0w1XU
LScGGX/4q+T2zpCFQFfi4sKU8wPmBq6pr2snzFcnNvU3vd1EY2O6icLPOm04wyro
n8K0dbSl3v+LyXiU/QA8gCNuI5wI+cgbp7pZB09mvxJJAk2G8cg+zsRVkTb7m8Tj
b1S8n2hfw2pB2u91aK3vSxIscSdtPEado3PYmpqL9Tg534ith82BV3EIf1Uc9Ly3
Rm2zDCWjy6/+ehCu0O6geawwuQXf9nTR4YMgkZy1aD6O0Cq9ODB6xL+8bzL+vBRY
yySAOCKUKM4Ig3XBBA4ppQWhPW0REasyZrfnClTxWb2Y3X7VvTdEGBMWj7CM5O7O
G2ottbWBlAv8+f5l0oLMP8brVQm+B+Uv/S9ZL6tLMdrFuiXBxwoHvNG43gR7DqUJ
h2bADkghMBKI7hLlWdEXIdWVqO8N44yL5Q5xZgMdHb2tElbVdCKCfaElu2AAmHW7
Y/l800Edb6U0DQbaVNigBJZgJbiQsHZzTm7r9F8m6SaTd08clMVFsQte6nF2yhvI
1MtRE7I0BE3kPJywIm4eAA1qKxaKJVNliBigspOuJ2c6Pdiv1wod9n+nrVXHmhYO
uL9gkjLgd1aCU/zjOv/LjZd9EGZcMPrk8tGmuDnoL6Na1vHvyA2iaT90g3u6Ei0O
UEseTOu3uocYvD7BJU0Lz5K3Vl0TUlZwDGhcxlyaGCeucpiCqX/EGu8n2/nulTnw
qs96gNuZoX1/3z+IHplAzS1SX5INMFVgbt7zvRZi9jwtD4IotWyIflDEwRvuqYMk
tZkKOSkjwE8AnA58od9qp2rkM/k+o27yPUsB+13wwyiU9TNtK7DQQ5nNKpjHrde0
j6FPFgXwXqbcKtFsLnrMDPBnqZWcQxttBPK517Lgn4+ph3iDDM3g7Kh/MHrnp2Gw
1eMJkrmWr12+66Ha8/srMaX8jnvREIvF4NqL1gVz0qPxI0R1zly+COCQJJhmqX14
40YrlhrbhLdf51qlWhzkl7hFuLESCSEoVGgdQQfvKvpJnRCUfQp39bZsF2RhK8Pq
H9Ru7ioZ0O3MWfPREH9AhJOkUqlI9MehC/UIafFMRMREuizBhn4GT45SAlH7WD8v
zZhWEt6M+sJ8lQpCFB4UAVCTetC6ZBOWSv2az6YGQOBJh3PE6d1sofeWYHKN/v6S
xFcMZhLFHnb5Sz1x8Ehiir9Fh6leS36MxMNgXdDl+cTYoOoGN2vfgMUDniLBkYfK
MOfjODW7xcCNWbXR3hxm7KxOyM2rWHMmQRWIBazVQZFFh0Bhh+Mzwsl+5xJzpQKP
xLUSrHAyhsRTuYcH8U26L2g8q/MisWfdYW1Wjk3GQHPKwoV6Cwcmvgf/tOci/QoF
5WeiGdAp56+2/G2xSXDbdIB5oic54xroZFV8je9L8mLG95GWA47PP/NP0oNNpwoa
bIQgYq4bBoPwJLQHRNiG1F+CS70uVFsGIFK8WoYjXTbDCf2h6IICAiPtmCbZA/me
ElJ7RBcJj+XS35WtownF4Seuokox4Zy+NAul9UhsoqigLI4oQgv7sAHRd9vzEaOU
4d6pZ8ciTjYPeBXVRCA520Ykz3c/IWkc4inG+dG3yM8CXTI5MNlANvTBShGzioo+
HTDe9887g1qL4KncgRNJG+eQ2qBKLxPmZy7dZXtwIFFZ2mn4qb/3vdoLyQUi/I8O
G1vuQcdrrqFqShWa9Edp6Nz2Lh8psqlX8oLWwnaNZ4R5HsOsssOFfftxNjgSi8Zd
GBX9cb1g5rU1ZLbeV3LG0bogYNIb8G052eEO8wEFxiuinu4EqxaCH3W5gQ1Pvux4
avVrADlOyE8EPKLgqz/7aRq/xyChh7HvRpuUDgmGjfMSOy7SR2QtPVn9KLiajkYN
fNMwPSuSLfDfBCuGUbZ6OmMpwP8PtoUX6hZNWMlcnIHifomuSFatOkC0nYQAp+F8
8tsvUm6tDXjzYNumzQj40h3FECXE2qborsXCxOGpOphDWx1NUHAnN27c8UzFEhQI
3ZDi1wgYVuN8/n8CTQgR501DgBcF5lEDF1Kbmj+a4jjvvQDZgp2hMzzjDl0R50Fo
KQNNbqO/0NNkwhmyVatSBVS1wfwM37dHlEA2uMTpXrZ7JZWATolmP2COxFTig1jH
esMKTcDTMUZeqtpBloBhpaOBbFF5DIig2rblSKMU7+dbC4SuSHHpfQhWRYMByvUM
syVQqqxDX0u6YQcGhEZbkCSNNfCBd/nqXbOJsPv3K/L8Ye0mjKaFNv9OndlfqQWJ
psvYiUSmXwqdV+yjlbmX9q3N9omAxGjhQTls9VDwOyJHiMc+3yP8S3mtjzGGB4yZ
ERel/DwRi6PMTYtRHofjo+nY77Q/woywlyv0O5pv1LJj8cmM8SFDkeUtOO6Eeray
Qv9SYWoDJ3sGVtThqNyk2LOhzdbSqbZkdC/llED6fQmkpDEa6Z5KnkI9WFNHAUik
aCleoskxdChL3wST/TnqJE4xMjfgqZNfdHRVFxWtMEA5ApdtlHYWj0ZYlOQNi2Hk
xXWgoXRKCrE8JT0ukfSXkaAhoAVRW7R19WNWIoVs5h/p6fGi4F9LVdTBfQlv0YL5
5eQ+g0A3yQhpU/DgqhWZnX1yhjfiZFxLoLNU+L888jjC/SRKJSlIJOqt56JR1c6a
D0s2C5uSCgXndUP17ApEQ+VKMkisl4K9zdMtNq68F0oyEQu8s9u3E4ALK6vurhK2
7oDjtJaipwSW9g45DgEZgQPBX32H5wtYTknX8UtEdojXPb9HghA0IZjJn/W2/TSL
EUm5MQADZqRETGAeWDPBevNNiPJSnGogmadpT+UIo2eTPOQUMEygT55fDCRQmh6u
C4RNbw+14D77LvYll0efhIHgGoRhBY7908vpHWyFvVQDRWGOmIvEZGBFsX3rY7uD
qkV65yg1u8d8yPN2BQKkpB6mWZ5jDXee68qWE2kHkx+bZ4Qs9P38VqZMvL6R/IAX
dq6QvUKjpAG+QVwDLa/AB+fYlc8m1PpnDE3CTu4MTGqQA0HvFN82WpAMRorh3o5E
7huo02FT1eYCfLPVI6eTDFCDPRzkpSLxQGYdyoCtzAO89CukyeC9ddBxxGJFDSVZ
myc4boT/G00HFsHCyYM23U6nJ8WJp5EBXcQ3EM+6Wg0OpQa92+G+NMJLVogcI7wU
DEN1nSl8vAsmLvYxlTK2rjDm9dmmY3MPoQq7eQlpM7CPd1s1Q7Ygb5g+MoFgTNar
cIvOMDwiCsaIvxs1s+NTvYSrhfY5jbMaCNF89fg6TZM7hVNRH0tWBLCQh4EkifzM
vu+RjRqLhqmqNAWCgy5j75rzy20hegkpx2Do1CsWjTcwxpf6p706fQhcCwG6LrJP
WtGxh1Xfk6LTLDeFWlRtlO3TCl5DJP9BezajWPatTlAFbRlmhXT1aQvcqSEpK8AO
MrQh7pUeTIOSGDrR0Db5U6tb0ltxOM0tIb6Z+735/0KEsVkBx8nap+UV90eh7zIq
E/3UwZksiXlj/31oY+w8tBo94K7rawYkaM3Cn6jWjfY1gJf5dpkkjSbV7gXk9I9F
Vfar0aWwoQpcZsJlvTgV36LwQdxkDEL0qIpIbcZCB6skfbs53xLIGN3DAcZoDC0t
l4ifSnR8OXY2A+NVNWaPQzPkhVUw+HYaLjNW096DhdUgOTOh5HjrUBWHiEWqVxJo
aaBc5fneRakz/iRt+W9d3jcy/6JRfNP3eXAe6VHjtesN86TS/b4DEEvHbhJvvST4
+TmH3bbSWw3qLZqF0CZ6NkH2ZpcQTOcfz3leWjXVvQ0PTrzMO7cHeIMr7KMIWcGJ
wKMKOHc5TJQkfIOQSatN5diBcxfIzAoaVea6f6ng1+z02G2aC6vO0RXLMNr473rz
oX/WTlawStgt9ppmPAbJWxSfNhUkrdBEyQ/zYsVQ+pwDBXdV7GZo9SE1usHxWyMq
nIuakUjFOPmuitrmiSl1gNSNNPp+jrmE8JaPR+SSupxzAO4ZUrrGbLJZ5sDjOj3m
F/GzyXwAWqnQguNZhAZ7PV718PZ4+2GbM2eXTGxD9HNy6w4LMefmy7e8AHvA1w+x
3Tuqa+VCULqQm9Gpo5nWo56tDv4Zkckrvt+u0DudmDffHdwjDL/Z2Juf7OqCf6lr
k/G47bhiiBZM0kRvInq3ea4PS5I/lbv7Bq8ENXUo8QIwVcfC+sK2VFgQRsKYZJV9
uQU8jxjQjvaJiShavS2coF5FamQ/n27NXwKQgHCIwvuamKubhyGUZYO+Z8i1/Do1
3qh549ikuR2o+4zBCvlYmAGFriGNeAiV78gYYhLeRYfzOPV28e5RJzQpn2/uSBdI
oRq9F+EQMX1pffcagblbnoIgqP6gFlY5ASCmzsYHtXW28u9btr6NuSee2iY16Nkx
uJLRwN14Lc+PCZwpaOpjTw4kdJcfnlul3Nn5ufDoN9I2e1J++XzUDBCBKAm2/czo
DdeE6JJioIsqmOw02dCng+fdz2drp5aq8IYXerREb6IcBri0J0ZRQ4m1pWH7DzPL
M3ymrQCkKe8merA3NmONzMQNWilzfj+IoKPmnxQIwq6D77No1DbOoxmalTvktyzz
NXTxAJVZYlAWM0UceVCGfssEdBJqciDIbPuoLRVPZTc+4s/r/dE8czekcFmBM3tA
Dm6I2p5kgq0wcplHw8YUAvedLLXXrxAPe5jKQzIz3SgNqbn7+vchNVlZ8+P5KWkF
60nH1317OYiSsfwgILhSweLkwANaN53RbIyXyOhl66I1aqZsx1q4a+xR97p4QaUs
j//pAZ/TKk5iLxuz3I1qkIghAhr41dln/beVJh/VO1C4V/XGb0wkimVbbwgg9Uau
RXTa39+C7p9F3MOHhfF8IPKE84jay4DHcZDjC4N1KXqF4JUzLv3McAGC9BDipb5t
gSLv/nbZgB7DWxHMs6gIXIOEytBmlnV/pRvhkk/8bww6OrVA8HP5UeNa0gYPREQI
3ulnPrGbReGFY3oT8FmWnqt/1FMXz2Z7rkphbVObfB+u5uwytp2qBtrydiLypDtg
FcrvZ+SBEkTC5fgoFQk/CmAIdj2XvZSbPM1TeNmd40ib+6zC/Nhzs/cFXYgC1Ie9
pbSSjI+LOQnqbKLFZjOdBeOX7V2r9uMzDRt9AwdYD9OOYlVXkZ429UL5klSXN4dj
vbkJIjkPguiC1ViB4yYoFCwx7PlzJg5RjdESuUf7T1+hggY2xN5v1KH22ubqWJL6
1oqJFFLkTXP4bi2tpHC2Ra5PzoOnAjj8/AJx6g+78hGMgT/9xiWwElLr5HWvKZSW
qHjGOCMyS38ucwXPYc+Nrv0sLgCgaf4KFCgG+8A9LR8xrbR/2EVFrejri78p5NrM
vwBkwHD4LCG4fvMmwVbBla3IqMSomByZefzUa+qtOLoh6TWM77Vh7weuvy/HvtiC
7EHKwbacXbLMDGXZWp2qrusO98lKiphwKh/FI9fRPZP1FNEpUnjlAk9H3FSJ9gx+
NdUjZ5BhiwQwaobUAQ3nEKqvt3Jr9JOMP72UpGgRUTA5EC6+lh92+IfUByaXblWo
ZPn/BhHqiA61sDTUwqtSs7nIKCShI5zUa0mDwFtKg+iGI+logwR3IVxSnZPEOGVE
bGQd2EPOVqQAZfQEdfFJnIEIz7WqMEBxljr3MX7+KyQPQ/ZFVT5oK+KuZUfNwXa8
tOnjJj11OonWTL15yzm8OuV2xtnqlszkLbQQxZ/OjfaqzkFffusi4tMDehRc3Ztx
ENjxaqzefodGCL58eS+VM0jCfxs0MflwOKkc6sezs5EZHc6Lv0IoJR6enb65ceay
uSX88esuOw2/0vphzTsWf3XhJwh0mFoMZE9zPrJhxqJIWHx0tYhWWdTL1/vys/gP
mqDyBspNk9VsmKRYk7IC7M7HhqpZ3KbeEYrIEhtY23WwE9fQ5H/ojv+FOnGuZ8Db
9NqFt1Rep2TC7zRFNVS+GREDSYIEls7kfpW19S6A1w1gTIG1vQWY/XKaIfUhT0pH
bqHQA7J86WoJ1ldHiQKh+DrnKS0QibsxIfdHtnt0+mUUpC7PyYuaTofRanCZnnKw
BujM2Y84wrYkCvj+jTdiJ76WKIH0N8kZp6kozsD7TMEjlpthY0pPmw42PnZX+QoE
NGCdyTE0B1K4uPQh/Kxe73OxWw7vtwCA3gupqidgmknd6L9qwkD3d2XFwy9lyvMf
HM9cCemTH0AGnKAkT1iyIubuy9jmrTLDCUrCAkzENDWvKFkYEYnDNIbr9LN7eEwP
3EoeE1wtSSE3IYJEZ4jJDPdbo6wvTeet07i6frjuckBfP93UXaIw8pKgw0fJLOVj
tpQqEyaND6L70yQ3901TfBQu3KbZcTVQTK55PeDdFFO9Ho4XL2FboEgN10sFpxkh
EKzkinKGvzZ1J9b8A1YLGqkK9DsZAW5VoaBNerAiei69zjeqXQBK64QC5fsrPk99
GhlBVZOsLrshAm6UUu1zGJBNz89JHGTBLRUBNPzsztlSHEmxaAMdhNHjNr92Yy5W
F1xSo50lN3pquCdimYxRSyMUJnZxcDRpBoI2R8VC+mDB/u7isz9ZQNqmqUgvrUsD
1lmozCBlOuKLAPg5qNVwNeINLUZyGP4fvuPKZhBdtU8Hb1ktoC7AP+pUSiaOLa0H
h3cnAe9kfdz5NilmcqX3SRZHvXhvnnWcg0YYHix4bhZ+mofN4PpCwFx+nxR2yKFn
xs8crl1TJ83ldwJ3xGdevtrjuMbv3L5HfX5EJ8pRJq9XmqcT2S9ZLA8rp/Sy7FPh
JJ1B+pw1HDZ03xur+qf1B48wLQgJd7pv93GHWLdxt3x2wE2KmWkXEaeWFzQuWDyf
B7UESQB2x+wL3pomNe9eCbJIz7h5KZPYhO4eX2xi55A=
`pragma protect end_protected
