// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Thu Oct 26 07:22:39 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iEgVKgPRtedqOb4uzy2X938jQKOEi2lPYwrE0XwBaGonTYwjcnfoZ91/rCfT/uy3
aA7p48bBuffVevv2Y6NYGcX1ZMP9202rxXerf4hQAoBJTymWpLMxrLqBgM4mslu8
p1z1FSniIXfJwm5AMVtYWvRsxOJrInEAsR9gvOnTft8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15376)
ep4StaPIRUNidNvycbxTy3UQNEl2Y+bPbz2CO65UF1RAF3Pvj8P9ZSDRnPzLtj2H
SSrjacVIYfwSAVT/MjH3fL9s+cXdaU7c0OlTXeO4CgpXFyqS/XOOouDKK9jLp3H2
dRtZyOc0LH0HO1yw2KW2t/OphuktdlZvd+xVVkPOMk2EhTh2Qk7POkz6YMfdTGGz
7rG96KD4G1+KLc/vk1102Udaoukuh7QLW9/+KKFoDFmyppKxNznkWKYUAR0g5izB
Zk/6tJDC6QqkleCXdtboSzTCHfzHWRtCLfeqbPufJHhWhFTN9WsxA+4MuBphJ4jE
xd6UVFKLUCWSpFrB5GLsGx6eyTlCJ8s9EKc4KMACpXV63YpVHaJpZw4/ktMmcox9
m8HeV8qMSWBCgUSXz5ICGtXKhAlkp8UBiYcBfWy3WncuKOWDcZqtaP9UBGBEtnUK
wLXsmqW8KK92j1bmbHc4faEJv6cgO1EejNSwMeYx/FPfSxmFyR1l4SuagH40sFof
rV8kntYrYXIWUKsmZL6LRYJ35o+d7ENnm3XCvz6I1Xg4Cht21yv+boxx4B36luHe
txQJTxB68h33vjmwWMEA+Hs6rDl1dRmSK3hKdH7wT/1XQSih6GQizQnQPhqJCboy
ysFXUfFpvjK5nXPR5YTaGvdDa4xsyl9vTyWp1qZJ830qL3uxz3VHqW+9GqOCsp/2
kDrlGKUqALjHJrQelOd0fmGfRzh1RzuPAyguAy/asXJLGA1AX5NZ6EJJOTJtWZZ0
4MQgkA2LWPIsIKScbNYbgCjZAvkDq2U/qBKlhlE5psbVikoCa1PpKys5RVQAfy8G
TcDCc3H/Vs9fYvHvUeNzHhH5M91rG+EMq5sdNuLEOt8PU3KJ3P3qJYVPVEPVsNdH
uq6wCnZOLNF3ER26S6m3oNdOss6d1RPDCy2fgJim1+szBof4gBHklyiAbmxBeMOH
TwwLaPuSc0NdhLgz2BDi9pJ9YAwSw+hjFVcveh9ivQrt/dzCxfLfpA42iCR7yZMs
nS55cb+sNqNyp+Yskco1dooWa9bzGXQ3AgSHSdGAdgvwGAAQM9lHEqug4hciiYSw
BPxlx+lEZXJjs6FgMLbve+wF9CYzzKZsYNmET6jKCyZMa3BBqyS+4esIkjUjojrz
VurUD8YY2zOkNwoI0Pd16C1H9j0FeD+j0bw0ic5Hd9aq0wQNLfyApO2gm0cgSvoL
dun9LogUex4+mMGS89jNkwp5irR4SXVetQzFeInrPWdsUxW1RohBYtnh64MoQOtj
e8dno/jH084TYK/KWR0urUEGtxVdLP5N+ZUOxsnybbCoSg0dbf8MR+l/I8Ezp6Hq
JFRR0or701Mk2APU2fI6Reo/E9sKCMT7NHV7gUCfFMv0KEFoNdvC3/Cdj0htbQ5i
Obm7795LZiVhQyvu0EzgwllZKluDQ9vREn22WhLKft/7toS50kPQEkoWsomMUj5I
IWyDQaHb9QSzmhW5PYftkAn0KBqBiAdjtRJ34Sc5bigKrP/RkHJiUaTGG9cv51IU
KAbIHy+T8YyLYEb0Mj/hqr/sS1z5YdjPi6BlTefC9O5AtKhoKE0dkLkFi/zzuxLK
exbGPTt5r+vcts5l5Q37NWUb4JXMbghEYyNtJMgesAV1TOPYy9SIsF5qLgrD2IKO
7ePNTqW1BzS/FLxeiF8syyAJ5UbJZJFAA4dKJzVq7+fQPx7HDQWNKwUcPB9QyvGG
KSQVRg5hRF1r23O2Ppz1pkndrNBDssN04LvW5ByVXXkNxJ5o4k0bk7LOb6Edatrn
0olga1C8m/IUherzE3x6Dc9KiGZIjbk3T3iJTBE3L9D+T9GaPiUtMCWFbFkCv+E0
cbaEH8ZHlqV3DHtIGyhEr3/sS5JL+CnQHDDxBkOXaG5xopFuut3ZttqVcQowF7Zd
nQFsGEymHSSwxHF9j+5jyMxdWLHnLLyYKw6MaWGw6OcasFKNkZXHAvj5Ojn5FKw0
UgnCdeJVfzuzbbxhwqC+6RYIaW4KvQmv24+/6Lu72AQlj11pOrAdVCyLhVxByfyE
/inkyhryND3SAFgL3WH69dKDqGkR4prTi3axArkL94H5e9vfL/DIy3C9gnMTYjm2
fkp7pEEmK3hcEUf/DgewQi623MJs4EU59XJvgcvyi5GW8MBddQHie16NSbsljDnR
EEg7z6ERWChvyAnz3Dy3Ygn745Bxd0zz9llFQ6m5R7skQJMSJzQ1idgKs1E4wuGV
jKyYzdD/EG/71DMISSEGx5xEDloJwkhoPYlE2ue958KuuE7KnA6vOqE1p+L2VxG0
S4ttYZ3U1hWTnBP586y36vI3ibV3n81CPnEViYr2/4fPWzGc243WtZnug821KSFS
FowyntD6Mmr3ZT902Er2UcWPbELBSR3ErElTvhHyzyj4Zr6mbElOhZeKFkxVXuzv
vf0Hd5vKaLbbeif/sDzmURg06hKAGezZwC97/cn0QL4V+n5PQ8yPrLHPvpUGypCJ
YNigy7yH64BpJEm8pXsQLzZm61VP8z8eV3fiJ4r/UJwdwdLHR8xnOJU/7ZXu7U20
RQiF+mvAfpMkzug/s4aekACRcnwRUZPJ1xInWcaGSoXod9rLvGhAifuFp0D5U36s
U5cIhfyiEQ+dLeuAnXk1KnPYwvE7664d1GcIqPJ21kN+fe5koBbQ01fW6ULbviLY
XQ7EUhanIE/DGf5JUUceyI8TbQWI1d57LCKmXYgWY1fej47lNiYTY0jmR8uT9goo
d4SmRU5VkgRaXRVzzqriMkCPXxoKIBDRffzEFplLZYnGV1Q6c4/Smbm1B4FE2fdm
EjZTGGEG973FM+/g+Ormp9eZcRbBe1Af/vx//ONeuCL5j4TLK7uOMltYWev4BONn
Ceq0TeusyK2BWLa4IBVCzKYr9b5rQ2wvdc3ejUqadiyYW7HNwz26NKoZ16psL6Su
r069T9228qC8kDn1mJlFhcTJIu30EZ52qS6r0CIQjImGcTQcVuWZgk+I5uN4o5xR
wROQ6FtgJliOjjocJ3pfbJ/+832rbEx9oFh3YkluA/HT9BoAwtqfxJg4K2sW9ZP1
jMf8JBNN/TxDRTyO4sgN7dDugUzn0xwtelVHGkomF3tUwQO14ezl/HTfmXQuBrCU
Iu0CDtxumE3TtwAwb0bVTyQ1jM1uw42On+LfckDdwXPm7DLLDkKuwMXNuW+2C3Wh
/0pa82etczHCz7gxAclbYOFFycED4RRMM9/glHtl5zbt8idsfcZKhcPK+yPs45Aj
aoMbct4CqE4vWNRd5NrLz1xfhEVdDis009cs9yu5pf4nGZgsC8He/fxTOi6hvjVx
sfSad5xs1EZg3cm2kFMzJ6DOBWZ4UCDHJwdao2XP6kKpFhq6NvMIzTmGDRnuW45G
AW9qzdnMEhFsaoGYfyL1ICp9LQmi0WhPd6vcRm0hZ4Q4wT6KS2QfhOEXjXVpD+Q+
p3I7OXLmCpzxQys5vs5jfzeEYlVaznEzuTSSqAKnid86S+L9AtXWtxf1M2NK4MEo
8IDpgpqJ2F7/kFb45QABEgq5JnJGwbOicLZi7y6y5X+9pU7A0fwvANKTq1G130F9
RiXHQZP110KAmJygEvq8qu3e7GEfsOwkNdSSW0Ji9TsHPdfmhxev6hYabTVdiGxV
FLKefhseOvbhcgY+l37Rf8hB9LGFlvQebwz1WH0qML3Pviv79Rkn0HTXTsthu6hF
DXp2lneRtklXh6XrsI6Ko0t3IJAiHqpUk/vDfA6n/NEOsoWd4vD9lCV6SzCA/FoU
6I6GMyLVKHioNrcls95F9vgMaylKR3yaRYmidrfVuqsAVxpxQKi5kvlmhvxDMusQ
jn1eOfNZwX0rM7iu3rHO44DPOpIvwXD7nimldvUGoTDhyorvhMSzlSN5bh5h7yDN
88lI7oqOSsErU25y6uLws3ok6+LEfeXpVB8kq0a50lvhw0vm8A5qyTUGTd+Ba4SH
AocX8bHsG4rtbr4XEblwjlTRhM3e9mK7ltuvzOTYd5KQt1JVjr099cjdHqIkA30Y
RVRchWl27LEHBSfCSwsWpFG5UR3+zsFSwUdZqh0tYiP0A+ZOldMgpT7+fovRsENn
1NCTSGGHFjBazzQHgdOL6QcaWl4EHNV0GoRIJu5Rzd6gRUhZISxy47jt2Gw+zE+p
jtvjk/s2bk2AFxxKi80IJ1vx7+998ZW8eAs+uf5UEihzasmvzFGlpaAYA5nklSjW
zMtoMOK1i5CVMfC81AwJNsaNTj2uiyLE7qcZF+1rsqEZcl0zJec/flUKfRU/m7Z9
wSQgV0RzIKn+wVDsMzImHSNoxWUMRKOHPuphd+H1A9CS+vJG8nZyEeNihH3WUpPE
Pk7TF08NzBhQ7AaxpiOaevXJNv5xsLdvX/HEi5u1p+ClGbZzmNM+DAIxu1T7+Iuf
bF1yWJzVdIWGG20YU7gUoRXqoX7TpfYq6gyn3s9LWwVWYOuPOrgyWKSWj9N1yUpY
jOGCUVJjEpL16C6tQN2wPNm/u6nZWFoPNCnHdSGfKtEMw4WhvKGRCrU3CQ9QbppR
g6tt4YFFJ9sAyg933qSykggzv5Sj599Y7cL92VlTttFX0laa48ZGvS0ebclfsIej
C8MfH/7i1ANDyehhbN04cp1USkbia+XomNwmW/G9xbGLGGe7/XpNMmWczK5v+G22
WwC20n6V/YmSSr0UZ2QzWpRHB3FQyoNq0eAB94IXghHaGpIWCg+W1Go0C/uA9sv6
Bjrh0VaIgQbNz7YrSInp7lPYJA+FYbvFEYW25fMD07UnAd8onHghMUXzkYh+Wxbt
hZnuuX/MUAFBB/8Vn6eQOvI19/QMufEmRjaf09T6ghs9/+GTcyWZxVu9xSJQlqZ2
u1VAdv8hAFB9PLopDb8vzSwXUW9BWHxCF8olKseacm1ClF1APV0cUTfRFHnRXPC9
wxdFlfajdlg9WmQyMiNafj/pwOzNJ29HYMA6uNjdDNbkUWY0IrchlDFm5WTyUBG/
pdu2QOxmkLu4jCm0rZb+wGtawjuqI5z+hxDDqC2O1cSfOYBEoAOiZk2Rvb6T1CQH
7oThecXBQThibKrq57XIugb9DAcaJjpXmpHBEVOYha9QJgOO6pU/XywHU7PNs6vX
TYhhlvdQCcHwUIdkDriS5y+hwXgDkEL4bVOSH0/YIJSR0oNi+frEjuOmVut7U/R4
VWu2rCbnXiI4M3mSBAs93tBoPpHtmhe1gYRbbYq9szlxgNXJE43wzu2itjm5mKyO
iG2/sI6H64eTe5prHd2cPixI9MKcYlMJe+0SeFp18NcH3AVRnQloQCRAVsWvB8rS
m1f/ZRk2lwEd9NIQUbSaUgvmEWvR33CEZ+e9jrQfGEvdyMyFEzvxTbjsl4O8xCYb
0TuGvHEXtLa/vHmsHdtEFqvN/azndOrLwReqzz9MhKao1Z+6O5WWuhh5DooI4JT5
OcFhg0r7khZlCpo1iicdH6sFFb4FhBXOPqIrEQEp5QzVOQOzdSgBjwvNuuJVXlgA
kllZlVPUXaii8z85Tyqh6pHxpi+EJoPJ2x8mOXPGVdwkRtUQ9HlRtR09ZuJT0IYK
YVJHcAhu7U7c+9p96NaUai4PxRPx633YOmWysPXHdfiUAnBFd3mR+AXkD24J9EwP
FtMaueSQrTnnRElZZ8nbV3iFOb4HgLuqg6sZX/WQzF5E4INqNBlk93zFK4riLs1w
7xPNieZTIXLBVKuLmUO/QPXLYFCi89hKF61KyruUG8Uv3VFKFULqTNGyBmfrVtZv
oRy38sOxKHylz5VlEB5esaybiIbRfRQbwjMzlZVUD+3Wte21+v7unuuxVLLdm9xM
Ta0fMqNOMwEeYNXNTbt+BI+Q0uTXAOn+m8Rov26qUkEezyyp35W6KYC5EogiX4aN
LgIts3S3QPEwoUrHPrvuYi5tYCEsRXwTsyPrw5UHgBUzrvfni+PJgkC6Nxizddzj
bNt8jMM52gt3e4yNECxkiybngD96SY3DsJxddld+q+1FOC/ACzwAIa1dx0ajP5t4
IfH9adcKnK9dxaAf2fOXy145OnbmUxnqSKy4kSBeOF7GWGDvbC+Dse7ZY7rDaKC3
PmfG5ebNdR3Jhp8Xu+B4QnYj7ONO+3PXX3UG2SsF6LB4BK4M6FSMjx+H4zhAoKcP
63kXqD47grOtuDNxXC65npJwPxkJ9QMH+qUn6V+lmeKXIDN5OLERFtvSsxM4a/Px
uQwVcAZAF9dl9MNvSvKJmxdP8QQXoD7yVEzaUcpHSbYWOsdiARwbIbjbFUj/+af9
wTByvVd8xbD+nSBRs0g9vTqLC3rovGjL/TQwt8DyYqIXwk8SWIDEYxFJ0OwYHB39
JuOViRk5m97N0EIC30SpuWUs4H17i7LcLkJ8YUwHarOcAKhsdgTErHg2e9xei0mb
UR2zzsiTxjbXHcWsskrOfUlyZDGc3rqlwT033Oee6koWumwZSl5z8JlnjHQaGG6B
q+rt1jBE5H8edi/rzRQi/ImVEQ54JQwq4cg1kZ26xdvtPjVCtVAsQAuhYmi2vNJx
9gChuNoycp+A3RJ9A/PcgimG+eE6esNqmpBFwxWwbea+4E4e7cGEy9wI1x1aH8sU
0owMXUs9IuqfYQxJQHVKm5SdK7ko70NQJ43V6cYZ1PttwMz/CwXZQW+XsZG+lLn2
IUrWkchTO0flUdC2N04BNZfa4S32/Gq3m8pBZ5rl/nedOmx344P6QOcOm0MyCNIN
C2s9xluCah7gzLUjYbSD8n7u+VJKLQ7VN/Y9i2hIlHc0iz/qh9EU2GtR4EUF/SKF
F4e1GTXIWPm7hvbxWYgzyS5SCCZS97HNqlAXtt2m/7YkqPI7Ey4p3QS3gZgUb7O9
SedxykaxnmY4kNbeY4pxk90hxyWyAxaLnAsYlcwJ5sxBuQb6bCENqgMyY9/jZJYO
ZKRms4dshsH5DbVwK3b6O6SmmKCbO4tnAh1GUCCHnOrZyrQ7f5fB5rwtolfhhtTc
RooJemT1CAYDy+YQTQDXYsHzDVn7PHUqsn6vKJ2lc/BhKsIzyEcBJ9nfQiRl8eOE
nUtHRw45sI62mDvundW2On15GnicRAiOUTEh675l34serwxms/FhhyD1YmIlW7mU
8dH/xKysLOAqBi7wHtkUWKwVJuUYxjaZkw5Y8azyJvB1jgFeqxIGg+y8KPYMDU+h
13EEEyEYiuS1JAJzWycNg5+b9HSLmenZ0f0WGeSgY85QaZvCYgrZxR8YLRHHtERn
Ybq+6t08S2KsIZy+cpbwAede0gQf06A+eEarqOcdUbALDoPDIrJAWHgOnEVPzMZ8
3BydraUsXwx9S99PmpjaIos+o3DOif5DPjgRWi973er6l4HtcLLVL1nl7pyBQbT9
pwicxVG2KY5t0wcWC1YTFg+GU+XuH1QzPT4SA7IkanGLlxwLhzsI4YPuLEOmdA01
JVJyjayrXEFDKIooBi2EG65DODwt3BRdqzMXjnLUOAL6IenEAEUeU12U14jYgtzs
7VBcHYBkoaXzw0j10yeT2ISGUcIwf20sKgb2HaGnlRXuJCgfv87d9WsnD/Ak9SHe
yi/rXivk5hN/BZI7SQcZklxHGq7Rm8jV2SZP5WywxV6t8h2VGeKmBUDDPPbKFlJt
FCONjL1vTbxFxPM+szpKr26YyMCaScr2val4OXQQmaSorKve2AiX6gROQ+pd2DHS
pWWoMRUnRQcxxKCfD5EcdiQ5bb44kUxkjTE5V6Y7t0N0kXL03qNi7l1mnJtuoDUg
0ssLMNF9qrrzR7oSpAfIJJxQ3tlfncyFnrNuSv4AWtWOWFqIKf3H8EViOQvc9+pA
X28kJbpForemVmOEx4SKrL2gkZLuMM8abdtc3AvEgkmVv6vOaCVP/IMHQsB6MZ5I
CAUn84+HXB65r/zJFAlHaz7d67oItCzge9KD+FtcYl5sUAsNlTzrt4Gp/CZCJiRh
JqQ81dSa5GlHeBrM2YR1O7oJK0nbxBrBoho4dM14+NCuxdDOUPGkzvuNHzpLweJc
GhFm4fVI137Ee3xcRKjZCcFlZT3elB+B93KTKde2M/bsmT0J9RWypK11zSDBBZCs
E5NPo7E18QlWG+OaVulLukzR0zPWAbPX/9TnwcxQxeX6ANZ4gMSHPeNNg18c4UY9
BBm2FwIp5MgjAZAcvyASlc/BHadfy0hujhnIl7awxDlOJptYbiNYrd1yAWpmybkJ
4rPFeQhe2O9PJ9mXuf39Y84bIb46wacgbMXwQ4Qb6Ig8uwwea5Nzoti4m8/sNLMi
oeagbMsMQ6Ukn4cGYo58oBSRnBISOfs1B6nQiDPvs6i868IqYoQHw6I3k+N8ixcI
XYygQKQI94Uzn5xe++LUQV6e6dFBodMi+eqdPDrgGvmRIQ0fZbDGXYkegPZDT4Ox
OvqDf4o2VXynEVBdSKngpjTKaj8RMiE19AACFSfVfKFgxX1PNYT3H7DupBDxQBen
dmodhQTS/ppdJuat09WXY6SG5FrZMVHeR7+tz3wYn3NUGYpgA21SqkhS3Hs0udlr
+BY+sSgK1sWSctx6YeAp3GPd/5OngBm29e2JPRRblpycN/r0CWXFlJDzDsC+IKaJ
I3aePMNv5iyLLR3nOLSxmKxbuTOCTceHxtGjY+mQsXy6roJpXPP8ULfEj9n0jiFH
3N/srpVobTkhm5GZ8jKob51FGU6Iwd8SuHdKRPpNeZEeevHasoyJuW6sXkvYVx9Q
VcdcdWQnAheSz0pcq4MI7wDfFWLbP0oIWS7XHpYA3V/CIBoHDXGBoMK8XuZ9qOVG
NGILpRpIBiLmNnGCH0NlBfHk5lyZ7E675/6ibOb71EmcXJWu60mXkaqNW5Oghdog
gJxeTtgyneXZ9Lq/2yYnrdgyZtgqMcCVBKQkIO41Gm8SMbeIHdWgzHB/75oM1K3d
9vBD57uICqBAJJEDQg7V+rxgRThgAFV5paBFzLsP7j9ceLiEsAolmeOiO2FXeRTC
s4EcikJP8FYffdxBx7BeOntNslDy1f0vKG8dBBl1Zp/Adsr8JJEsCsCDtd1C6cZ0
CB2pjK+IzPjQlw3KNaF6S1uENTpz3AMvGma8IjyOkP9J52QeKl270tUm1cAqMoEi
8UZU2EYIyveiUnbxYQ6U0ntWKxCFz6e50/hECWGMMhGFBtg5BnRUDI9px4EzIC6j
LnVZNY84SzGX0IMqDpUiMr3pFDat7k9JGzhkkY+USKkhZ7daDh8D1eTCeRs46N/m
9nNP10SglXBBnUrVEN2iZIMaZZ5yGXPPjm8JRIbjdtlaMTRxZQTrzVa0R4oHfvm+
9jGNNrlL6CzLNttPUoFyocP9k2lO9f1Mx1+dM/37uPU595Kz9PfdjEHn29TAhy1c
qqKGhRzGDUgPM6anhsW0tOuHHXbz5XFI5thFs4yQ4btor6DwfzGPzh6vvmY1Fvug
IvoFAoPIu+hv7W/7P6YVQ6qsqlHhek3ThaO+vqDHHRs6lx/PI0iJAgKBA9ZtagqZ
bpVRGQ3JGwGZBNMqc4cuRprmUy/Vw0r/KIAywulTEB8dZ+++zNHRCSBqyPun7eG8
4tB7r49J4CBG+sblop83+Z5XdSfuJ2TEmNZKDQqiBYDISqX2Tr2BFdM1rCmI1UUU
K5LZLTBD+d8Ux13New9qD+j+EICwxhhlcjQ1fIv6wYuPTQH18doP1q+Ntrvi02ZC
vmdk+O8gyq+NwkWOo55Q+ZA/EtsuwCfkUNdJqK71J+Rf5mqsIPAkrU+k8P80a5h5
z/M6EAHtNRv4O9HtVemxGgjMbZIzoR6vOk+TCc5D0+A0E6PKuLu9cIpxDlbV/A4n
OEhrU+LeQTW6abz1ZoEdcf1nnM2J1ez4yzaEBCBaqNYVweIG5b1BuQm+kqun6gjP
DBxRXh5ptH01RbGGMpuS/kfIOVlp2M1Y8jsojMK9IP0kh60Sawc9f3xgYWy8LJUx
NM9FfIU/Mz+0wYFLA/kLg/gTYC4Lbs3jrSxbNo6e90i8W4wiiWwNOEJDuSkPp+gZ
au1fuH+UBypc96YKkUIrqEaX5iLdcctdVJb5vtSOfZ3Ap1HpK374/Ufp8PpPhwih
hXJMqEL0jwzmhxiM7WBK1XxAa2jbRCTg4WscYAJr2GKvU4AnG9p99/lofD+xbgad
/05varhFGJ6yaJ+K5YlSOf0JGhNnVaXiIzRMPNwwfWOndeE9G0hcpLd6Eyv30CQB
7a6pHalDV/Xci2k+dZpCQoRMFh+sgE+A8SOLvXePRcPLSV4jzJhB5vCsGCXZjj5V
Op6vryyK79oDzj0wffgsw38TMUG8POaEgdi2o2bngQkmxudbn6oc7Gn4HywBWpAP
yRkGeqgMvEga/1Gr+VUeRgToxp9Kvz/AXNZyxvBc4ZjCIWyR3RNu35a+8RtvSzZh
/6h3bfuFpfXeIhZQ4lCtdzQjMSf9MnGZ69Ag2jaHqk8o9rlr46EizHchYzS1GEEw
dju7wHFgg7lqWjeI2g86wSbFrDW6uA6/BD8SuES2gd9iZ/9kU7YraSipGUxxBJ7V
6Oe37+K+KNefjoiMqciZMW3z4IROBAUbZrJj8y7fQxWiVfM/Ear/ByiC3J9mwMWG
Ym57iaKSmp9fhehf3opW3UGxc/RN9wXXcr6M5Oo85W5OTODeEToPc8kxFmU6bhLW
+5J9PoxmuTNjocx6MsXCab+Cx8/W5zDH0192LJM33CDwFxEJPyYptWRAhmdIYuU/
o2/oYaayt/Pp2vBYakzgQYeSEgFZGK2D2Lhn85alFwlUPSRnMLQE21qo43If2mY9
Y9d/trHqmn438iQ1qZoMMgnlcEeQ5eqvS1VNSmAJaSAiCcO/4IfYODcNYM7S75t5
CyUeOaYWmdyXa5N1XNYSeekYo9C46hPmQY7/zOJZ1XSb3VdOPDOocLqs4Vw9CDNg
LOdWakGAKRhsKMLm4+RKZ+58YuVA69gt1O/bSsVMg4RPutNoGbFpwW2Aon9uDZTx
tydHHrDMRE1kVQ48z9joXyBKM+cpx1Bze188A+KkNbT4y+DvSu4s5SnX2MnoQ4iK
mmEYUMgvj3h+HJ1I3DJPp8DAJaS97ogGFkz6VpfVTszOJMMnF+YRBnxkNADZDMKU
EjCp5UN0mXea7tYLc/wdGnADXubkntbAjoZOd6SAEsHxjIzuDSby803d+Rvqlu5o
IK+JTWhL2SirCBKDKONQ624eJACCv2wuNqHU+osMfQ0sWfXpDSWbmOvNUw84yd17
74tXVy4Yk0uYoQws+KgSBNHr/P3ylFIEaWH5mKLwW+jbov7bwtur5dWDnMJ3rzMo
frw6fmE+SrbeCfJW/CWbfEVVMOitBc0qJr7+i4akSAn6jXS1Sag+6drCq0G40K5r
eBsFREuN7gwr4fQgGP8ArekLfMV/40ZQf+tBoKPG8GM5YJHJUYgI73gl3rJL3x8s
0Jv8oboWZxN+fTG7n4La3kis3nGmPccgBBpIFeYny3MQRq+aFFFACOoOdP9+SWg2
wlm54Yuv2mQQQJKqa57QzqO1Ox5yDoaTFgOc1jWlD0su1mKIg3f3jyRnn7oBmU3d
415Dzb9Lq/5/qt2vfPg1lT6im6tz3M5RQ+i3uwRNj+A+p8nl4Cl8c0jpNaB357uP
uWMuyGI00X/FIPIK5GBj48jFdQLDS8dFHPhIvFo4EpxTvvCNCd29HFp3N68bZoHp
V9Lq6aCT2YdmoqCqDBTgSn3B523wYERpMuiH92qvjisvq+vzKdHO8AoJ8k//LqWp
JYQE+lktuJSGl5fGnBv+LNAlSVb4ug3e7lUWbKKoGBDeroMZ7eGxFh9dbWcg3RfV
N0zO1mFfsObX+TN17nQNpf8w2BAMLejx/hOg+2/otlwQS4tucdP3c+i5hAw6xNok
4FCeDC/Xx77YOOzzp63SNhSuUv2Rtq+xB7aRY7Y0fQmaHB63MG4k72cpQHm7Z7XD
MWRonN53Kt8G0/+pZSL3xmFY/pskED7WY70dfS6/9Do/qFKK0AX3kKn3wKUG75+/
W++MADabrNT1e30vIFbMa0ORc7IgPXEPk1Pphb/kP2uTlZ1xOOoTggEF4KX8HMgG
fJikClhLJa8r5zeCr9cLp3YHqsi2At6HpXRVb7s+uRLBpwT1s/Devbel69pAu1+S
vt0FoDUNwNdzEMsGHuVH5Ag9TkFS06ijnVYoMICSKcnODkfG55fjEj/OPxf5dRX9
ZDykcLRWGhBxKqWaYqvKeB5xkRlyyhog4YAvtGmd3Ed0r9zytBSYoUzS1YKChIIy
f2Prt/0U+kDvQVofDpURXpNg2m1Y8QRFyVWeS61HhbA1+b8d3fv+7PiSdhTq2sXG
jabLDQlj2z5N0xXuSu1YpFJVpEm3sezvDKrYyYNqr8pNERwMfoL7Q9A2pgiEtio2
nz1B7w1ENLPAGfyqzcffQSPoGuXhJ/i3R6r8T5y0TaGrQ71VhDYnBlsxM3JrET9t
CC7Ksaj2qwvZmh0y+UUoL+2+cjro5c4M24+ypZV+mB0Pt3raoEhj8uZevr32Ox1v
l93P7rOV8X6IIjgREmW0ZOoM65Tc4uo3slOnWtJD/2hSoFujz3hUMBl4J2emxqgx
Ggq+a7uctnf4GvFoJiuDZpe8ercD9ZU9s2sFV08YOGz4o0K8vDHC69ZoGmHoyRwn
QwswdaYtQxJAxLaf4/zahTCPy9RHuI3H2CxuaqN95YvQlt6hIc2N7hlkQB5K9lQg
4fT7VsWrFiToxSiIh2i5WCw8Fz9x1uxqYIBF8n4dNEapd7NMNXAzHAoLXHm8GKST
vn7klkn3TFAenGjSme9obeJq+Zze1V4jtIUhgpn/YqCCWr6X64KFW+vIfDR3lebX
aCAkq/qhFKOjcyhRNIs4uDwQNBDcUTzj/SDplF34kSsKLMjLHExBPvJXAh8fG34J
wz0NsennV0H53A0/H8QBw2LO19Jzu5vvo2Pc9z7HpZTl60ByhJlcrI77pg1olpBA
A0d41265WF854phava38yT1G9QZQrsojisDsE7ScHGULyRyjPjOCL9yUJPJFRnh/
q0s41ni52VhRHBgvP1cBXlO5aSSfszpPBlQ7lPDlR1WxrhFjlU3XnHFF2aqrDa+e
5ZKKZcqXzn0WT25ZC9TShPwEeQ+YpLlxjRwqI0q09ifj3BJl2OWlaU6AVflReGPs
5otSORKKuNhrEG7mVKL4wtQU/+7q7Xcsp6o4DnTjH8S/ueTIFsHYeI4vGbRC+buE
7m0gDSmzQXOIHgyPPHL53lSI+oX8fSKx23eU42bDDcrUJHa0GsUJt8soJb4ssXxv
2pcebfpErIqg0tuVaQqYxQB7ZUtzc77Y+u44vuJpMvG+8mwkMjKCAWvN86wJ9ouV
dNcO6MJtKoD1fTKPU0pyuM87Vxe9ubcvi5iiVbP/jsIbBk4fbod4pw6Raz5Wl8Bo
WOgZryVhDphjlUYWuJSq3MILZS+yIWauX3+pBEhWLL0tZVd8as4HegRouraBOLD7
w67ZYtmKMMN59fpXxXU8Jl6nnqQM3PXLxhKzdk7r38rSOSrNMWiJ3W2f/inXpySG
QIDr/mOMB+TZhuMnoLyib/kwKzdvasPHGGipjFpEOBrbRM1/n77yYoI3/mIAV3r7
BBUpcsKkkzCntEX8xZfn3ZEwr45EWy1CXh09aJRi8XeDcX92qyrqTUpp9XGzsLXP
WTZ9d34as88T0KUY8RU+RaV0llnFFkVVykKipIR9Yih6k9Og6D9G3cnCmeh+y4Bu
d4gEA3tkafeRL6IIwrbJ12aBD3Mj6CeMYIPEULw+Y8tTb3pDfdqG41HsMtH6tjSS
9ubMwKIWvTZPp7KuU9bQZT3iJT5piWdFyk1VTQq5g+P/ps1Zg/z3DBRf1wnwI6LM
nlgowH0YdAl2K7bjKEflkirnrhxj1FFdtt1v+VlU2k4eX2OK//VdG9jiahopb/ow
lpSLiTQl0Ij0GGFGAQQPjDMhUHTes21kQGCN+Pi7xUKK3IbSr8/Y3GtuOb7xXsjy
2IMQsnEueW8VtGcY+aEdWgf8ysaTePxSAomlRSyCklmWoMH75KoByNO8cArB0aya
9h+1E2CnbY8W/E/pC6rJwjdqpsZwMlRf/iYGv7cazsz+yfYHuf5/+uocBEBq5TsL
DkbRSEJXAeOhEJHAn89a1x7UUfoMHlJEFNui+5rvydk9i0jK0EjmRqZST3bwZ3pb
epM/FwepgRYFHFOco0fnKXBalSbWSiYbYqIwsYFJ9ShaIB1lBToc6BPAP4BCabxs
yhly1/G0iLffCSOfLV1kYlSfzM/QL7iCjCur8mCN0+6eOQQyjMNOxQeeeZwOi8LJ
NWaSlWygsx4FThrGwIBCvw/q5RoNvGDnTRZ9NyL22pJSj/byc7q6bS4J3iD10M5A
bPyNz8rweT/G8PRX4lKtD1Juz9IQPbdLbKhHStl1RMt4dzftVtuZeDqjJ+ydW3Sn
FME5DmV7lx7KodZ4K/on5k//pdyZycDF4Lz4O0IAq0DyAUMK1mfODVKUxWgJv5wE
jyaPbDFdRET/Ao6a8IGU0DgUe08GtNaPKlxm4TyD9B8/XYrjPAnSwGvWCetvSjJN
Ac8txiFrD0eB9KRRQi9s4scjec3EcPL1/71dcmf5oxYV2laTEG3uHbmq2AXt15of
TARTvx3Q43JHA5ijyBe6TXFneqTXUGlmqrOp0gUYuTaH9YUzeX4q9dQjZ8VLVFGu
KDHapojfCLX0pOB8/fOCE6YJ5QK0MrrQrdZIGsX28Gx95syr8542+MiOHv3FBO0x
jwnXkXSzXNkmr1heTY/4cIJEUYGYHeI/4FxEJh8ngQsCOhY+0mpd9LIUw4Lg1RbZ
fDr/8UFc7cgOJdVQQKLtFRnr691fLSBzXcycb1oy6VjjxCkmW97A3/un52ZRjiml
I+SW6Hhtqf09n2rgrSS5b8659OjRZk16o4BzBY7F2KCfLgHgEkjgrOi/BVZ4D6hC
uZzNDFySg8BsyQIER8vLK/ZrdOBP9iT/DlgDzs+HIQM7MtmsDopyKmeZk5ZWn1Ju
mRdmkybMNglzaaq4L5rm6rx+LouFCJXNCrcB40keqya3C4mzn9eCb+gaSL2Nj32P
MQymCgIXymVZzSF5VzJ9574KuN6wgmLJrzoQl984LiJODQ+QUPcUMNVFiiWm4Yr2
dpfsmGIPW8re7v0ThEMGRWJmY4GH/pN2oDvvdXrGkccCYyAPCi8vgA/vLMT/Nq+d
lMqNPWXaQxNbEhknunb0h1RFhpwe7y6WSpPXeNOhjqZm91XJWZ0SUc+QhZ6VUBAR
qdxRmc3LfSw6LEtJjw7+Cuza8jBJ7l3GVvQETiiepkO+Xiqp+whSYhnafFEYgDie
p5sTa2xi+IoqnW3j/v/CNaDUFIFVFso5t7jdiSDGMIlDvaiVKg3JqBrbBEGtzMRd
xUZx41OCfgz7hP9R0PTNjwI+Uv0Rl/ymN9oUn+iurWyU9ZcCZV5zxvHsvkfQPZ4g
SPjIAxkjqqikvignHAvVhSzjxvCQFpdkywFlDn3LuiM+2cF+c1QfAhVyhOJryaOT
bYyU86KMsT7yDRN96ggEFEO8dEtAEUstYP6Ku2pv6xIeIkKCP5wbz5B+u8qxJCsD
oqR07PEMi0fVbF5eNeRr5z1z3MM1HLvQfk1/LQmKThrK6vRQPV9ULMpJ3PxJETwr
Cojr2ZhqRpmVS2Ed7809nKgLBYU+nl/Fz1ZkBAwieckNvFHKlZ59jXvwvB5430Wi
Z5tqLyMdbqfHCVAqCLKkIajGUuQQKzLiB8H/fROEBwpAp9ZbCF5Oo1Hsew2pJRnX
1XRTvPC0v3QDLnbv6IjY/Vjw9SSjc9wnxdcSLNAfYrZigI7b9BzlCvjqclPjxmjL
9kAICgcqu51cfSVoPMJqVw6XodHLdNic2nRCwLaGutyiTvatS8ZyVuuE0uGKuFR6
cbEAksBGYmpT2I4lcWY6YrYQGqouCtdojzAGKW2IUBRkSuVoUGAdgl1Of7EKwEnQ
NRG+eUJReWBP0jYYqzFsIC06ThFDqaIfcd83hp8oV0VOVbdjrd4/f2SdE9v6cy9M
WDaiO39bBl9vgxWhMAZLCvExDpVJXl7RBu6ZPsFPQSS9/j21yh0Z54THuSniYsOT
CUizuYsA5P/8ofM0lu3RGmO35EY9uN8kVMGrQhMQphzvCN/Eo7XA4mhU+2amGtHa
0AnrVmSYdBMDGEgMqJ27J5epnyLfhx54c13Rdloaj7x1jmJVhQqtFMoLJsNwV0ju
C62rC2vURSPoeKsqcHLv1SwN1HZH4Xzoh2LHepGh47djsmT+DuQ7MXvT5hkhIv2X
i4ruUa5wLaBAbdRABfJtOK3Gdnpo10uF0BwdAHsAd5RjQ1Muko6p/+LkBwgLCXM9
CetaeaczlYPBhuRCKfKY7LD9VFiogwwxTuXwv+6A7/aHOxqjkIFltn9zVp3GdLda
wIm/usaFetEcYaRqoQPG8OzoNBXwKc6Nqm9DFwZzAYiy4B2vDdaFJ6GVs0h4hEfj
Rhv+HiXSZj1+tLsmdMAf8CFStsqaU9nCRg5CZuzL96ia52kzE+QEQxpt8NTQBqdI
Sf/AMKF7IdQdNiEad6U6w4/LxO7ZpAsVhBNDPkMCpU1wRJEaDEVZ9BUVekUQ1YoO
hBv8yT3NcH79ELG7da8c/SSKXiyjo0PHKA3rL108QT9MLr/CSFIzATBA7LqJPbR3
CnsI9mAk7Lk8owzFgqhpE15ryrXknkcJ25RfNca1QZ+U4aLBP1kqdCR7YGIEacln
oeKLr7pNgbUsKeDiOXNK1P0q3xo80a9iasEMlPNCxcFeD1Ttj8uezBNzo48UEEsv
xDsajKd9t5X+tGpBZx1xnqGvoH6uR+qzXzFHhqCJNAQhbkt2xTJQgukTKCMqDnsR
L8Lj6w59M2z9WLBxZY38cOqpbJtxg06kcdJUeWdQeRKVyTsKuBrlfJ3bK1NNJOjZ
Z9aEFaFECMCTHOm/sdhY1yNJlux/5yUWsPnNcntrXTzjgAUmlu42hS6z3j4MLUGq
dTqmY+sS8tfdlfOBZek4MUSww9wOD66joGaOON4e2My2NIAWSmFSC4A8Up8nayLj
9IlkCy2zoCVxDAMudXxeNDOhWXzRISbSJNWWWH8gLdC0J15NGRGdxmDS9U+GBFxZ
h+xL3FVdxSSXHJqM5svUjkEV41maj6mbdndX9DNy8Go0NLH2mH7LBGTYstiariWT
i5E+Ba7gWtrFVC4mV1o71Xg1wW6bD/OUh0Y8Uux0qcyFfXNc1wk79UMT4fRXRubN
tetj3HM90Gm6vp+7ljwlaSfy+9+GoAg9A1b/+vaIP6GE3kYWfvK1pEkLCN6pN1M1
xd9zUZQ2rcCKnoRWqOzNixzGsPWzwEKDyC9z/3QVqBVqRHNwbXg+DvDrTW7+zE6W
jCLQ+4E4n/Tlgpupl/0tqCVI5bdtCuLgDqy9/kapF7vGRSb0f0UcHDLiVxqwKMQ+
Mn1UR7HRtCx5wAEea5f/OU9uT1tWOgIgqOz+cqI2+d86P6OkJdQjnCqt/897jrQT
VlmpghGUUYsaH5k6rDF0pRjQbDUllfaF5cw+jBzUX641fqcAg42U02vRPUomokiq
nBcTe5e+LQRNCxqpbyHElXhX1Qs33YX2UzwjTDx5Bv8CwLl7OMC02ZJ/RC1Esjwa
d2sSTc3T+JhwV9148qqx5630QxPzq+H91+tDlhhgR/g0RsrYJ5OSoUwEuS3dnOWo
l0QW2qo7YiitKQ1xQYZaF6bCe7lJDz2LZc+inA6Z+LZMUw4r+O9nhaE2xbRRF1An
4Ubb/tVG9YKAnJVI0hBTPsOUFa2SNlau0xFhM5Nij+ai757W2Om5LoIzHG9HrmMM
YPnMk1wwSFL+Fqwr8t5sAk2gTzosQKHqNOaHhqoMW38XL9jgQdvtEjE7L7fQcN39
2fIJMise4peoThETqHLj7ze50cb56G2KTK09naHulRV6nMzq39nHXMnETtto31cs
kPDZNJTXYPJsV6Wk10sgtQAdxDqczMZPcp5Ff92N/pM4c2C9KnGqLYTlyJjjJjCR
vcn63pl5YI76Lr1rDyNB8GZfSSqCF/fmemEckgdCDMOO1g64/Dmwdyp7fAd9d9lE
lDUK5L6OfS0VillXRAncSyGZlIuqOGqPQdWOFUoM80hvP7JuOU/cYKB8/H/Fo93F
UA00Vi5YzvWCwImtdDzdSO9/wARys8tyOiA+TGTCwvCN7bLv8CnmaSOr+wmT3cmF
eOKPvh/UO0tTZE6W7LzAKWFpELm/Qqs2wrvQue0yH7Cn5f0TnXfHprDMuPZdNzoH
kmyM4J1//CAZ6bb+APYYojEEAGKvYX8W+2aDxSkt6eINct99kGoEtAW0tNUGOg3S
P5Kx1/LnV83zEMjCSgoR7Sotr1yuAsLUF7QFCfCfKeZGK06CSkE874hEvteqQCUw
UPQvlOeLC3R/S/F4P/DeSPFaTCB8cRx4QS8b6uZmmjG70hW9fOs2llFPWvALehWb
W0ZXo7LZZBHUuD0YZ0TjU12PjEZoU91iS7cbY9rk4eQjsIFaEmfjU24dx8578WUn
NO8Na0r5RBpAoW3pnHZOzUkJHqW2IQEq+PhHuE3HLmoP8lYklDnGfdEhpCBgFtbn
61C7ji9jHDH4XFM1bxlSP2dbOC6706bcf59dqtkm/i+u2gJ9HfT37UVAJQD6UjFC
tpwfW0v7ZMF3LrEjWrGJK8qHlIWAhVlgZ51PxI1Grues7oGniScVnYhzb+yzqh2E
H3HdHiajoI0vTeEGxYde7H7OlfTGOCwHF0P0TESfRBqAThytgIZei9dEN1kojWgR
w1cMwJRrdeCMLpfc9RZluxF4Nu3gou0z5NFVJXJplMuhmiTeyjwrMp1a2lbLIkI3
IYCF8Gxjy7t7hj6YpgYMrC9t5REjlIFZs6h8Xjo9Fk5mPJmxS8+/ovl6QnkZQsTs
thEawQgermnJYXU7p1KJHEQW8Gb+6j5IcgZpam75omFGcrfSVT5pb6q2IT+ROuZF
PvbwkhgaoAt8jBAo1HqdWb9+lsIhZClp9l6mHyffUNRigj7r/o/GiwZJaps9+vTd
p95I6cJpldO8CfhAx7UUEjj4xVV6zWpdz7oKX/a0By4EOaX9SBSYsaqataTeFMJN
QlaNzIsvHasdJfD7VrECS5k6NGNGHvL/Ict3EC6p92SeIAQEtu3nhfDBa8vPDPar
6DZ9nmX/yTdRx+s8gh5C8u1wkJBiHYIWduDQwJ+Pu735ds01FW4B511blRg3yOlh
0Zxhw2GRgPL8cK7ySJeEDAzAG+338Jp3WgNi/70esNx5SIRZD1+YbhjMaXD5qp12
YKpHZ0qHXv3ALYhA8/lF+DFtJg6xniQnBMhtx6iIX5j8Csg6BoQELCy6vc6YZ2Gx
tyfElzidVILnjNgkxg9NTe0NDqE3j7ZnRZqdKqd/9vF860DPLTK2Nyth0WFD3g7W
yXzrweMltFNKBRm0vEfNiU7hY3nGNZ3Up5l/mP4mHO6CtRIB/OGdSUnBIP3yuaUD
WMl3Hd/ssTZKKvlMcfF0rMiXY+vc8J+mYWH0i9mpUieyGCVz5DYxAWi85hhQm4av
BejKaJFxRqKE4TxjUy+dTZVQ1VSEpT6w3frwQjTEqIxT/8WX/iM+kzj6BKrN34yw
+6nYIWGoTTOmOKQhGkE7uDcBsslAX/I7KViy3vlLOZ7W15u8SEo+jH9KUT1OV9H6
Vd6s5sRIQWRH4M5ocl8rxR+pSzfJd+0ibK6POkerZlJivzfeAcBjD0G6uLxsKx/w
l5pIoA6hp7Sg70tmSReuswVkiB2FOy2N4vJABWrcigxo2tMffDssqT3oiEQEt7f6
5OJAOyfW6WQwW9ktfc23jdDrOzzn1XjJC87DjITac40pQs8l/fp03QTWuxd4P694
5ZMDtwQW8PNP+Qi4ZJTzjS2+znvpmxDClRqjqYLSl/fWB4QE2GRID7vN8nt1Ru71
HD2L/UNKHlxblLPSXW6Yt9VVhFNrdZFNne2n7kh8OoB14DfaEvv13sQzdfhGePV7
BGUiPRmQVpCEePNyjOZGi5jw36Y690AiE77CDqnIFHZh89QOy9LM5VA+lp9LOpOh
jtTdnXt6pZMJ8/tc2RPTxd4vX+xayPShdMjDCTDf4lGLxu0LBEYDJC32nLMBHbCv
YG4bjXCVCjLbIFReXLyT8bbW2KdpRdxNV2oQFpIBL/DUXiaz/Abmx915BcPuPHkf
nMH+4vx51mGIrec9X7h3MnVdu0osQJ0g8xytwFTbIaFmzNhrtKv7ewTT3t48oC+4
6AdKKKBFW0X7jEWn1q8OfphMVu2ZnK9HQAGkeyICPZCH8PsqKpictVoYN+d3j2fj
PJvYqXaqLTn3IOQ/MB1Cyp3LwFRgeGBqudDGYKbL/qM06clu7Oapg4rCBm7suz2s
LXAui7I26y/nzMIlOBdEy0jSi3nQfX1H4hHw09z1xYNMe9jSd+tBMLcJPvIeKLVL
4rKX/Op2hGlpFfS6Zue1CZiaitJUrIP1pW8HNgogs7bH1MTRhATShCsE3EhrfrWn
4as7LAWZngqXaRoj8E6NAQ==
`pragma protect end_protected
