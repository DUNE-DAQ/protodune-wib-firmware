// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WKG5ccUNK4wpwidRfT+kCii2J6sgH6XmCd04ip2h8Nx+jNGo8EOdMMdB0O0eLQgm
3B14ct2u0iw2fD40PcA4QD7qTgNP1CoLx+vvYtjRlS3qGhxD4FkThqWRkGNAN++B
Bx6aBSR3iX73rToJ94d7Bx6Htq1hd+5PN+uZblzG7Ts=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6944)
nqlAVuk3HT4R8Juulm5Hs575tCnt5UG3BwAYhCcUNqQj12TcVXXVh/rgOphW4/eO
Jmqr/5j0/4ih9vDcMUbqMNh+Qza9idDsDDlQ6IC6t51adLpvJb3C7gs3fJ51wAPb
DAWW8giFGyzsnaOmznUao77ikAIT6oYPKUqEytPnsP0h7vUx5zip+ScYlN8rdChG
plvmnk8JSsQfwoqVThGTQA6SxdCDVukbg94cTRF3Xj5jrzxVI7afZOH/Kz/L84Tj
YvPZaLw4VZUmnArquusd1uqkDjcgDjQ3eQNbIr2WLz3AakQ8YZMdyxLf6ugQIlc3
jYPmjMhOWqtGTBUwCLfWUAAMYYDDJ/ONIYuUcVRr496Z0BUezZueZZL9C+CspJcO
XOtRPtngRVaNwIKWDXnOYw5zGDgpgO7xsn2LTwBBcxEERxpfQvwbd7W/V3v5wD6w
5jPG+FaCec5xM0HZh9QO4tqEX1LP27tPWGjaXFAS/BXFOVf57FL2AcoHMOPRllKC
vW5p238NPIVv5Y5C6RNNxGkQNIi27Ipc5SGhZB1DCGdxlHEZypLXwMex/m6R1OYL
C1HhQ2ERrq1qcYxb6aPxCNYHY4dOqYnBzJI/F8VKfREjT+5xLi/T4rYbkylwfnCN
RWpJm9pfA4VbzGVA9Avc4aiYLHGjbjR4UD5eI29/rSljp045FiqZcXJ0E8gewo3E
vtQ4Ong+3QKkIplfVgNqW3TggyugUNxnwKHBB6bIhqWDlJdU821pDUea/vSnrZJ2
FSaLldJFt39QmEQ4xCt1jVNKE7nbOp/hY3VSvleqX8bg6fFeK74p0PHSfEycPQDl
kjVD0CwK7/z+6ArUqFC10hRCcP/dqMxxgk1Wnxo8qZB3s2U5KWgg1Csfk8Usp+iI
/WNfJHPPOfV0SmYomhhu+GJC/O00PYZU24m+QPlG8MtqGWHnuyLNFfYbH01PxHmB
4W83hExYSO+g468CM/O2NhKH5jbWgx5zoaZSXTEByQKsEiYDLZq6VpgaChBek+LV
61VChYqLcSnpJeTa44+1csuR0rUXJVc8t2NcofuARFEflerb0FbWwq5b4Z4pe1eh
yj1GHgZj7Ev3JTmwqSHEGT6XTYrZD9eoIXvqiviZPxXlV2ybiMZ498s2M2+eXgqg
1cnhpU9HmyCEoltsMsDAHBh5mMQDLSJnfFFmufI29JzzUgk93bBrOqLrTAk0hJ+H
a9lUBcg2KZrjrUNplEkCBzc+lM71m6dT7mIePs/rmwzWlx6KEy0OB84hlWDSYAxB
fUTWgX69Wkpqm6DvnKInt241fQLQHhXFs8XAePBeHDBLLfwQQYPDn1H4vmACv534
wfYboy/pL71eLLNiJNxBGXvsnsWdPPrErJ2O3zIppa1E5usQqwSySwCkyrQgUhQX
pqfOWfhwlNThJI4ko+KuuACbqqknU0HIUaVhvaUV+9rO3YqEZxBrQ47w//kuwA6+
TbxzFuYt5Rjl2QQiC+vYF4MI18dXUf+DUGutZSKNR3tYCXjefMzECj8d71CHiBI1
MU0Pru7RKZ9OPMHGiLaoP/J5usxDGSkG/aOOaGig3vO9k3lWQNjtcDGySe6V3E+q
teYmUj69ZZXPTm2wVk3KpkdSEXHnEj2HdiPVTa+XzlqPNZicEsQR8RM+bl3jqJ8I
CVwAzZNly1N5M32a7ddG8itbqWM5UDhLWgY8PZDh2cmE/LERLSyaSZvta2xrMm5A
DwBH5k1UNk2Ln4/4OtsAJo0lCuHzf6oaB1RGJxGfU5Pb7e4Py3CySzUeaMddGqFX
KggRWxNrMgt6HkdENJ33aRfCyfhShzlIU8yT7PX2hAxtkJfPm2jA9fwVg734lI+c
5r0OWobOOvaWAOmGyuZFEeKmtSkoEyNRyzRT3B+uvcAeafWWdkoLTWysiTiRc92s
vHfqgPNb/EY8o4O7If6DDERDvlCrXB9ANAfZInRHQ8JTnqwF8kpuwjalezcjv/Dl
ncLon4inkzr49hKilri/TWoCot/2WHWL1lEizfHMfAYeH6ZBtdfZoHSTzkyRxdtZ
fdssajdMKVyOdBuUMbKjzYhuRH/YuZ6mk/KchesB8BwfWohIt8MRC3iBCr+H/uDL
BQ/shYmE9tIWoIzgs2xPLMpv/sBUVAagEny54AbFI0A7jRnLO0rAkqaodaoBn1cc
r+yUwYdk+biIVjrYaB3zFkYm/8GnwBWWqk0kFYLtyPX2zujbWwPwNHZliF+OeQF8
n56C7SqmxV73Z0R+HTRsZAZtxJ0c+I6D8Mz0eGadUXnl/HtTopxHsnHCRD97caaV
xCraNhQCslGPy8Gi2jTwbuFVat+VKLSkDuC4jddACfJYaWN9/NDp4tOl+ZgzGKUH
zWJnnngiIoxXhN0osxkgvkK0hvMJLS5fUQb24HsT7XEpHBbYvhMExZW5AA83KCjE
Oef88BxGvHRfgaXiXCQv+l/g14W+itaCakZ2Ppg5qIhBYOPzTgSRtY2NaaxZTral
UqFKdSSdEeQPVoYU1lbhQDk/R8txntJ+EEW7oLdunA21UJqNrDR/py1CtwW3Vmxv
Qz4cJVjzsqMS3ws0kPgeETGmA5ptTELb3j88B0v8qcK17TS+nR9lzQqJhgwxMmD0
yK0Kh+GWeFyuf5+YpUsXNo6NTbwDonnsHe6YcvvCSw9iAZdQRJMEy+ZP5g2sazg1
WKEjmWEOAVzDeH/fW/Path0FvKW4jyAo4zzZwZiGcRpMUiqxGJ9Z2UTnoM5Fp1HC
tclqEuiGYo9q131p/hz61V6/mTv6cd9vSBYtWMCn/ufEqQJWzZmLHHfRmY9vg74v
JvbslkHic0ED+KpAcADWZr0H0GIflkpONFmPcfM13KInX4YrvvSzBBMU6DvyU8OB
aceUGrdP/RUOMdBJ8J3vHWRFyYfZ++nnxMl0Yxg37xK10vZdiZNptrnnCjHrVfdW
K7ilol+k07omCENXw3Zh95IEYGxtu7jf67OP/ikiod4wyoH7QsUFJui10NM59q8S
grO1a+D8rfAQJEi7LcJTZU+SNou22nUmGMGlpsJ4rRAL4FsNwy7cAbeMIeeVlf6M
nms/TIrSPBZuVX7L7dU4lMLEVCzBs7Tu3DfYEWd7L2ey/IFoIDT+pODLLVdJ+RdV
vKKecz/k3bCggpVDlI6yYWJnnZVKcdrHsYrBdpX6uOp6pjGOutYhpkyRTaHnNySY
wZmP/xMhMiQOOhdmjvEGp0qYBrcJP2pqHxYg4KAcTgNUhGdJw3jvJoleWI0B+e5v
W7qL5NnBUyi3WOkewRIj1KXy4N468eqKSYN4YLR4VXqHpwNyuZBAjfGdkB8af2lj
JmhiMxxtK77bomGCOiJLUTyBCP04tMHHpmQe3TV84JvZWcQfXvKtUxkWPgEQ/Dos
Cfeviy0suMR7EGMnzfjJbzHCGsQBdMvkbfjeNW8MUkZK2X9TrYzTT/FIfes9eig6
qR/28ELJ7dmPRh51vv8nnTkYvkvcRxU34CJYyuCTyvhtG8v0DvAoN6m5WJuUTxKH
gP44DMsoTmidZ8AfJQ0vgo2ahp9nkoqi6OPba+NWdTsfZNHk6fg3IOd7/s2nUgzt
nVwM49oad/gw3rS1ERaYhem9gL5rPG8FDAYwPN33u/FzVgbU7aqN0/+zuO7prGwg
qCn5ky+o+VD9yBdnN7+NpcLLIMb7cfoVFw/38U9LnvdRyUQw3IBZycSqa0cnPX6P
NvaHTnO60BphCb78SDtC3irqTIxXLlXz2LiZPKNVF9NPtL/+xHilin/ODIFlfpQy
BIgicSkGTvBbgCjc4fNxTYv1aVkwBZuC1aarAEYLZ95moLXizBekP2K1RKWDl6WI
IuOcbnd287JY+D2hFaayq6qfkVMips3Q2h8HcEeEd4bwnaN+dJA2ja+pjzzr3sgc
YqGe1GopogSu6hITSGBNEuwoRow0uz+LbYBjlGCzY/MLEqBkAC3na17q7/dYgOf3
0nbKdguACulOfnizlapvK92QH9CFzC7/JVXLI9CD+N7wn9XRRhqfPgjF0hxK+EM6
TilgvC+PTA31NBFJoS1c2W0X2Mvr87xI6b1jG2lVGYpmoSmPLT1Er8n3i++RAD5m
BEh8Z7wY/xjZcHMxmXr+5UI7KgIzCyCYdA5seQ05jLJBfBgmlfWopS+ZnlY8C9/m
3X2qBv62VGh2DzBoEb367YYQ963Ep/sEku3gd5vY6QeDB91ed1AzKvs2R2tf3BbX
ZgkrDsGUvHt2Up5Ku7ynHo3duITVQuIKJTe0ycbg/FcX8UtuD6BpZlVs/LoKJpRn
MPExfh0kXlyz4B+IjXZnPC+9xsUKFGDs3S54yDvj4ofnueju/tazav06vYed6ISM
yn0G2F5G0sIVhuqR4MNVdNiiVhhkhx4JReseQE7l1CbCfqH4F8T7XMdgAMFJU0gx
cgjls1Erfsb3ay8SJ6dXY9hw3VKbbDMZJWhMPh5tXxXKGTllOntDaxs2MYlbEvum
G07pwNGdJXOX6/U+mgUorcYomBLqtKwA5QIAfcuLE0A1FEEHeaNanRXxcDYgrnLj
VDDKAoHYkAG9CYEpbRyATpZDHGcuIpCOSusmwQrv1cEvKs6fWGvUr3i1JNh+yg9N
O3RlmPsFJ2ZDEDWcw73Vo3FZxIn2oE6d8SSazqXGlL/Igd9m6xYpn/KO8iRcOS0i
y9xb36hN9pcJlJom/fuanSfKfxj2HCw5Ge0M8EgrhxD4B7Z0C9Zbvi8VZQRyoYRm
ga2AOIK/cEwC/BzFf4T9ONngCJXF6Y7HM3RBXmtC9uvazwJp0hUb/wZJMEBvdluZ
akbvaDsYvxizN9BXMJqjB06SUIzK1feEgZj0BITjw//Pw7M+hAkSrQx6SuSKLA+q
F9YVPrDvcdFJBTh1A+evTYmxvqdTKMOhRmgN5po8t8aU3hDl2O1ttWVlSAP3gpz6
AEaCwkrG5BlRMv9aATqVyMSHJsFfLIRQJYRz4EFNcFjKA0pcyazcP4/fbkk4FDm6
Y+MCAUz6kukTBr9LOgUUavECJZ0aYFaBrBk0G39xEhoDHL0sCYvdFWSuRbO/A+JA
oFcll1OJ39IS0XN2n09hEc08lTYfH1qQytKAV9PAS/Tt1XtrpqUrId1/229tgPlr
OT1RomQ84Be4+jbcJt+38XswwPHRxBNsLBE5/0whPj+8JKsgOV34p1EDQ9WMZO5W
v8uhuQuSFVRn00hvM0BvEiPiZYV2+PKA65EJ7I1mi6Hvh9W0MPqP5Vsl3G91S+ic
8/yRCDO0WIofBVqZAr2ocosXRYKoUByy0a7/S7A2yvUB6O3o3begfPQixijhG3SD
bNiAN/aubCdfr0ZhHyxiZ9Ndg8/YTioBc5YPDcQl2JTTRE36buaj5rshBCV8tUrB
MA9878RwAPmEdHhqIEH5C1rLaf5pWc7o0fNLeFTUaAz2g/e/wlLZrgkotj+5dCYx
FKHGiea8pRgjYi+g9eEdQv/dWb6pGDabgCfwxP4sG0Uq+GSreHumGbnksI7uiZa/
C+07Acr6SYWd3MF8VXQb3FcBCYkc+gF/HFfYT209F8jFlHk+U1xAgnks+jp0kQeq
BkOyEUZpjLhlqw6dDQaCGvnW8uUO9eF/UMk64/D1Nk+AuhnnXBHZna+voz1HrVBE
qmZWTdU7+UPK1zvHZWQGIr+7CtZWiNvPoNebp2piom2NB/QS4Yp6CcuXsEMRNcMw
XV9vzkJYxBI5vV7cstKp0mtjVHAcXGAj2ihQaUYu/n91yYvI4Euww4PxFBTA1q4t
+eIBHEssnVNsYrD1QItubjJasDOQmWJvlJv+wmq6uocv17UgeIxYqFqOqO/+F/W9
xB7+tMo9qkp5m863mP2Lh+M6K0HypQjFSc8YD4xlb7OC/d3cIMpy4hiDLF6+45JO
BLwbVYEO0LM2TBPlO75yzZHfKmNwPaE1BjvgMS/1WofGIEKSV9t08GqzCssDekIT
6Acyejmo7tI8B/PZVcP3IyU+q7NkjJmF5+OJE2tZHPOHkEr70QmKCm0GfkQgd8li
xETnQpABn89N8MdBO+pGwwFYtQR90qNM6yoh8MbjPDpAF6iMz0fJywJaq+PN2qbF
lQokoFFMXNSMAmY9a8eqndaBqLPzux5FmxgOshMjdV8SjOVX5BCZnrUr4Br9BZ8U
IUdiwGm9DdEk1RHxbW+VZ5GQbYqWLDprew9xng5eFdbT0YTZ948elt/ye6Ft/EFN
0iwKqTp3oa7cU+2j+yLozSpW6f9ley/mJe/p8Zw4PH+TCtLvFSvor3y8/n/54f0Z
hkj1UEcqc1A1QBeod+ug0MDroHjy1mj7uCq0cXxP6lSY2GGYjMlUmjR2gI/pCG/o
YsC1HM5PwbADnAIyK/9MOm9+EBdWHNnU+XeuIzycbS2O7oowa/d+MtlApFTFP1bU
iYlwa24cVWgRe1uEggDyAgUGSCs+LcNvLeX7AJGYgg488xa7bqoNUXbSJirR50MM
MPSsazI1sWkzP5DbrABffH1SSzU1iFvGqvH38uUB9rG36Q4McDV6Z42L2kMW3rx4
cnscUXmVUUoi+kkuLrAVFkBVceZYg9dlS0bayNqJzUtP6qtmJxmQe5kCJ2vPhLFL
m6OwyLIfxhDlH2V5E9Dv3c39KlUsZNytWa9wmz3oDXJwZ7Jl1NMLsgUbQ9q1VChT
TPlmEyVRn/NoftxYMBou9vp+oDtzhFN/UuKg+x3obxDsMGAOysLATcp9Xp1z8QCN
1D8XpItPAZb3gcw7lUCAhdz/Vb3/fNmJhRoxyiIGTsYjkkUcEPSKHyjNKnYwVlF7
FbehLqrm75Rbwou1Y172uEzxE4TbBds5FSGXcwS4XkpLSLCA87r1LUUyI5CEcake
7bUwsu2tIijcK78++ys26M93e9UACgNtuRE47oHNHSPpfCgS95ClUYBJFUGjvQcy
Aul4e25UAF2faeJX4hWSRU6/T1ERN4B21SCafJnM51LDqYZTcAPluxIZ3lYcHF1w
p/0Aoo2ejK0ZdQKYvY4uBsZ6P/af/WhqlpMjyAXZ/XpJkTqPuF/OYe0Q+vi+L4QK
Bsouoqy1g4aVxWYb6dlxbnCRiGL0OxoHV22b7THDaqRODdzI31UDvTTzPxZAEh+B
ckSoSUs2JlRZG2QmZG18i0M2PMRiNshwDS8V6oIL8+y5RRmiBgTeCZRDk8BAA56w
E6nbuAzy0ah5XVxyaHI1ihIBjt0aq+xzsXQkS26/6seQo+HUwwo5dHE5ooHtoDma
8J3eLDct0JDehfyk4Rh0Bl+FVtUytJCeEE/OZNIWEvm+7XAVMbwaOm6ONmkoIrjV
nUIFm/qinE6AsI5hoZBn5tfMdLDdtgN8zSX5Zu8esL13QY4D8lgqel9RF9K5Kff+
Mz3LFRHtf8Gus7QWUzED3zeZ3O4/SU3YkgD5zbxUC8fdx76j7QGY9DlDmqnFZyrL
Tmlom5K2TThyHAex8nUGhV624UR/uTaErJ63c/l5JLq3qiVarCBcDV6v/E5J41zW
blOgzQmIRL0FI259P1pSwoRL8DQRk5KJls4gGop26cU7cadgd9aVvlrsY8Majxk/
uPvlpYdrkE6gZvYI1DkxNkPTDM9bd7DAB3Wl/HyA7Y0zL6+OzoTCzo2aBbDDOVj7
DMxcg3nVMS0QvqxiOX/e5dEsIQQhVE5+zXpwGnBAYDFzlwV6b5gmawA2UsKE0VH+
0PcQqNEvKQDQT/3J2weO2LrH5ij42Bk98l01aIB4sbN8bxGwgM+qjq+dbj5Q+UvO
Y4bEWoCiA13TIeAnL8qqGIYCFoxlaIkAbZmIDtFxFpLB2X+DUQHEQNoEQJshJLk+
/b4nG6dUBbWTKLF1rd94NSVO5Uz1BS3HPRFIdevrllgKuMuaPxWr3NH5+9/8UCzF
vXVNdqGY2THSfe+pAtg8NwSuP6Mn7NLs4CU7lIqWgMr5FNUn/sw7cV3umGppPndS
/2KjW0wE6D0tTx+xkBEHcw7loOww0rknId9FqWZ2/n6kNankfjZwKOjUl1oAA+5k
K2aArmmFig/1/PWAsN0KlumYXFWfIY7Cx77fck3qhPnQETBKNKaXCs55WNk4FA2j
+CAdEefg/kV23mEXkkSUa9zkleL60c1q6A/ObCiluIMbZ6BN/ZNoHvFDAXJ2nlQ8
vgcva8R44HVY0KurL01Bfwy4L85X7peWKuBvxs8GqNe/wlLNzPIYRTHvaxgsgLas
aDyi0UViB4gsMzmzqdfBNC0mK1sPzFqeVOdZMkbo7rsL05XPmj3QwzNHT1cMGv84
u5cs8JeN41kO/0wZowbAByUFlSMIR049ZC+YCSCZDiLJwui50Uq9Kw4igqo0nsl8
rkAMOoltLyzlOp0/kc2k/H7PN4+RTXddwd8R6kWgwdvhbwYbijp0F92ObMvjMGao
BOo5q4v2wYkch8/w4e1A4kc1d0bO1O/D6XfSkMsx+pEq+JTyivulgQIxETKb1nFM
7L2NV43iZa4NiR2gpPukm41ntYv6zF1ggV1haLv+Nr+mvooTPt0r53NW4THhhdh1
CCzOjiLw/0feiO2wzP2Ltrsfl23DFbHzDgA41oJrHZJ2sZilnYvhZU4kPlOQc8Td
l18zCDf+72L0bOoWoPwTkInAyMVeob8gG8RFHYThP/Uy9sg1zDNQqb4zcot0Isun
2dyBkwsPxQk7zEumv97nMoyLIAimbIpb1DehXKeNgqy5XcNlBUakcqYA9fakDtId
OHhsWgPVDvRwSGxmKEmBdcF5wvepCKQ2t9ydJAeMc/uNlCVPbSyUcw5jRL9JHwBg
stgoLSlhC9d41BHLg6ofCyOpvr+DE0pcfynP9/IcRRkymGlJCp0ejlnQk/qEHUXj
+kALne6rQqXaoGkV3s5ksBd64O8sfnFh9BEpG/6/ZdMZYDZ8rIqKUF9hhy/Mn2mg
yee3RebuUl1I39FC8rqfUHAZjleSwdo1GC0yNP5i498RAfFNgFwGLOcwuwi95+fL
UAdb5RwGpueO7NFZc2saElbNmM3JOaEUhW76zHEgSmP8upuU9JY8URTZAF8P2Yqu
nsYpgzDiks7FIa52QtZxumLhTVQXiuxw6ybUIS/UBCgX2/63phQ6t2bezNheC9tk
bPHEWe5fWGKSaX8a/O2NzxpnUWC6I7GOk3x1J9Gp9HXOd6NDBf2xpsLVPZjOjX8r
iGm3sXIWL4DCN3FIXjCNOtQ4kmxIzFrYiP+nclRndH1BYxORUh3kZIsEY73tkgIT
GGxkRTqNe8ewpUX8gpxRSTS+g8eqhJnZMZkqGX7Ycgc=
`pragma protect end_protected
