// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:46 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ckkDuK/CF1/yZrpDkkw2fNkgL3obZ4AP/VRn00jbB1WQAbvXy4DPfxlDmhAraF8C
gmCQl9B9lHsjMphOw6ZmQDIdMTDGw0DnpwA9GHF8YFTp9HfAcwo6jeSTah8eOjKJ
tAu68DzDnwddWtxqN4q5Orv41kIkfT5+Hpb1LJVvmrE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30160)
aRK8irf5Z6vrJjTU235mno0P6MphO+76D8wEkUQ0BodxIQY/IaTCrSnLpmvhATDf
eV/oEbzMSXJXC7uUmaYgzJNsCXW8QWS/ZDQnbC5l2SzR7T+wdH9w89uqAfNoXDS9
uhMLGFyYfH/Hgs3V7kKMM4CaHNSj46twNygo4mwHy7vHKdhgsXa+YmKGT1lzUHxL
OV/QkPDmcBjYRY3SgDtdscxIihIZ//A9hKEmXdXcuBhVa3WX6i9yZ4pj6YLqFLb7
bzPRvNNJ/nqspPTn8VqszKvImlzbIXd7Gqu5N/myv1Vhr/jIJUldS1NGVdUzmWWZ
eZj/Eicn6pKcyY2V2sXROUrxpjjTEcmVQkgFcAL3Q/jMn9XWhIwhOXrS/Q/Kx5xy
53sSWq04UDc4drcRIcSd/zC5GpgCrIBdb7puPhPVjUGaPWgZ0m+YNwPAc5dYqGit
T35o/DDVi7Ypmw+UL5LpTQozQDE/8hvOUj1b8sQM0zieDT3Qlal+w/9PvVQ1QTJQ
1Ddu0XRBi0Tkdpqpi3MA0ktpgAuP3zPqrpwKHGx376BDX3kJkIWQcuYugldMIp+n
IOVlEmsW2pHPdxDu6XV28FpV6v05osGbF3Q71w7JA8Gi3wO5QiTW24Qvpi2NyFOh
nBVbl1ZzrUrF6gtdhZJaew1QITsGk8+jexJqPsRy05MquiMJEdUzLTcfHW0gbwCq
ESSA49rYtvd5Hv56ybaxSry2mLHAW5P7Fu2hWTiNQA0769GEGPrzINHNYzBp9VVO
6/WfYgh4UJZqHu9u1PO2LVhX7gySkfIwsR8KhffGqWTDbPHcHT6x2u7kSL9T2wyb
UH2vEsTPc0ZXc6tibzOtuA8RkHDA91d2QS2aBQB0LAzcPN1/k2rIFxb0yqn88Td9
X165E+76udvK0k7XBui13wwuAgY2FycvuNT/CpAkeKPnF60djL6hn5BI73Iwlmf7
oZYd57ZumVfov7ZnTfvTeuucCW5j0kDq4GXlCZzI0wiUiKuT9bv2P5AE+dgmTtvr
k7IHBU6cYnCpCiB/mzIkN410EJhfr+tdBrAVSniVzGjsGemZiS6MaqXZMXV9NaiX
XZI8172V5NitEBSgJSDeIGtr1pglS4pMaytxCTjQZeejysAqJFP5G6nKSgOAxDGs
38P1j1ewU34IBvAfMMnEDPa9gOTAz4L46zAOU6qnNXA6IaHB7WV7BE59rvb6w57s
Ladlb22P4KvwjlwpzK4meWWa592GmGS1tb8ABya5PF9AaF7unAg3jrde+itAPaD6
j7bnUDaV/osPzVEiV+IgNe2eM2A2WFm6jUdTCoK9o+jtsDCcjD7ZCN24ySPtJsHe
5PJzzb7qDEh37mwnDyWRW4lP0o2vYCbpA7/RF+GiNND71wVL/z6RylG9M38Fg4ta
lAgKjHIgmeBl2DNAIE3SsSJZrzfWdSMEdJiDN9rwt+ZvV1586RKfQge2pyq9cyFr
2pOf0ZmmO6cmXCyiDFn+ryC+VjRegglp6V5SImSA9bEqa3Jsw14d02qF56pLUDLT
0DGQYCRhYDYvr7WglKaP2UHfk/yArOO6K+5Kcoxs6N1KdhTBMl/gvYa+L1z5odie
mlmqnd4sQhdMjyRoAjghS+suP6aUIpYJoCAV/KlbqFntESWEa+AhZ4oCo67qRW/k
hy/tjJ7EJg2i9xxfIejSrWJCbJdch6ieEYF0F5LWGNUzJggU07IibIvFHz9L36no
MkZVejrrkSChxMGoih4jzD9bth5hYs3Pk/ZHv0YuW2Lsi2NuDskJh6ETthDGPXDg
oj6T6EP6IgyMWqR1Z6pBNEsq/0wnN73XWW0KsrhqptlG8soPklc2ArHfCg9WpVKt
rbCTORcvNw5y61y0q+FKpi9hpiU10cOqj2ZM3ThSxYtZmgfUdlL+E9ef+WnAVn5o
RqFg+DaEkxlVlKDB6h3IuPNxpzFievjKw0sdHXByE1NL3bE+ZvFaZTprrMR7DDtO
YdMtc/pn0dJ4b3a4MgCMORauElv13mieKULxK31LtU+k2R85MtEvYghL0w0cwcyI
YnkMhs7eUJDipVrz2Zc9t5y6J55qLszCRgriSMVGmazAvG2TmhyYmmzCA//elEkr
ETJ00gNa84Qo4OjKcCx0MdHikGKT1RNoKBfnRRw8IU4MRTcNGW7IzY3R8MYmbX1P
VLrWbmsy5+utbLS/P/cXgxV8eGgNd7w6WZrEQilcpxSDBR5NK5Xv7XKhqFOclJdu
7gia6swFYzkynNNKIPGYvtkhV9ko83UbNEH0ww/G2HIsP8rQ8nSWbcaRZd3uzbQu
8b2emPHioj2RwTf0Du5D8g8P8gttym6qJdpEl6VU74BdjqgGcIuNxaosSQz+TLnn
AR+Ubmkc2UexHfzz+bbUv7K+ul04FOoZ6txTDdVcHChg3mZ0S6DmmWmoR0z58R1F
dqbaEf4aYSq40xDbP+qDAfR8/y+rE4o4cLxBbQqbtxrD+xUUG/9j4a9hCPRpGp7S
utbdZZ7wNS7kuPRtL7XWIlN0ZeM6nyqoYTu2nTQW6o3T3ebJytbl71xTQm26zNR2
L2jJDMjY51ftfMbIxA9Tu4DQMY9plPNQ3wS3wiELfJuRnLSUdSt3561Nn2oW+3/6
WzbqEoc1kXeWYBMwkDHxAIGgMRsufIzd93Jz0+siK0NKbOiGLdQD7Z/QdGLBCpdV
OaBrzwRsLOiDSEedv8ohSfFK7rSJOT3Zp7XHmZR/GvsxWS6NmEaXTkjr4IMZD8Y/
9httN2zhyJLGAiQipDZdKvpTe+ouAHLGT+F8BxZ8IGdBnVmT726D2PgjuJT49rL4
lV3Y8dO1GpjkoCEXOgNnXlRPlKaNAOs0ygpiIX04jc3sQ1hAGxaqUEHbim09wy2c
wxjoxlTOTlmIRjnJ03HbzFYM9X1uvAS4zuZuFgrnP6UoYkQ5880mbCzi9NjLpgIh
ARXGL/P72N96Ct8eXVIF/DTfKTNgOjAWPJfEw92965W3ZNPq0c/D6ycSc+j8QF20
Lz8UiypXKcdNuBOboZHpKK1jwN/X+pr2qInvVPOq7MYIQ7vV/RCw7r1DMgxZYApt
VFSLCp6dlnuuDHasGcc1fMsubMAPm3l2gBGmTsqxCRnm6QsS2o6q+jengG7MysbF
u326i0GCF52Jdqf7SLb1xJe12MV1vTzN7WMF1itqHyLg4FSBC/9QiOBG0JzLl18M
qYtsUnm9jMLN3p7PLHJ00D1UO2H60Vnp5yOIvQ6SomAm4j07BuipOfijOirj+psb
ewuSbRjFz7NighP6kTABd/h33EqgsVCDcSaZNlpS6vum6uIE0rOCXsiaxjnWP906
sP6WowCKaINn65jvHkMpWvUoMU0J7PGx4kQSs7wXHqtGLLC/y+4d/arW7gXm1alw
5JtHOmB3tI6IifI85bA0GRyapP6dnHVkWjMPhkI86yKLfWv6vIO2wf7EGnah+IKN
MmaAx4UQztT1qdIRugaRXoYgvc43c8PmjiCkmijwGK5WPYPgDp2s76yx1I1bxjDs
4AApMpujTplg/1GBElgyKru8bIlXWDkW9r0YEeHaZ0fs0JchzgfmQE2/1mlcUSCO
j5ocdZ/0av5l4ZChVBuiLzHsBlUNj3bHERP2u/mMSWRkk6viLk/Ey7fgbfmLPPzm
apquj54sZN1JJwIjRrxeHg9lRbP2lyzxkNk8UXlaDSykf6bn3k4360NhjsIOInJf
VGu/q6IDa7c2RdeTC6IHlTwVN3Oh6keoDBJQxNrfRhy43L2e4Wdb5ew9vhF2whAy
OFiztLD11XJ9rZY9YFYQgKtPPDYLFUV8mmezK09ZGx77BnWCG0AwtK6nm6iko3Fm
wieYxb3aFtusLepnxQnLREbw/AD3Br1Mtj3ajwgiK2NkbI4ejfHPH9L6WxCFkY/A
uu6dozypjagVBjVSPDROzfkPXMo9c3E+WhqWsEfourZwsN1P4hfIVAGKQPDyR49k
u+BBUyoLvxF6k1m1BXCWR8H2ID4mWA8jP0Y+f90yusqRsUJMMPauY+HxcORoXtof
OMdVRZPQVgy0LCAx3C4H0rhBvcfoOiDRBBlvd3pLA9q4S0YdGmq1tOjRgUdl6+Zu
8lEukgwZeV/Uj4HCnewMiuvv7ZgOuPsh9YQI+XTkZ7AVnI36m11OD0LBP6JbEOAB
C6Ui1NEjoGuXE4Gj6g71c1R4WuDyG9hxIQTz9lUILR58HR4byNbWLc4eGFkPje6R
EZjypeHu2R4sUygCSFlojVBP2+S3Mun6EqSvlz8QuHgB0zkUhsFK1//Z9CcL2yNq
pxge9vRkXEoXmfvzzCtQbKuqeUv3tZWGZEXlt9/b5mPAL6r+UzSdWc3khehAA7+v
IKA6q9KEKPvjKSF5RDge/i9X4Xv83y9+ZTAC80QZWd86M2CMN6k3RZbY/EfKw5BM
rtRYRZmjF7JsLpR++zYBs27ZvPsgI3OwM/K6DY5lSqAGPo7Rc/uZsdgMo7L6dEy/
eMeG7PFJuc4GBSxBeFW1HuQnZjVtdR/5+VVe1TDGFicOeehysK/8WnmPHec3S2IW
jnImmxbIQ9moxshmAeLHa4DQvrXCPl8ukgHDUN5G6o6ukVEjnv4gQfkeiKnrHRkb
9lKJy9JyYiqYkjhUgHPhJvlKE36JtfzQZquNbNS644Fk4coMKMyvjDuTvPWJHO+Z
E15U0F46yyyIJ7gHomYWi0hp2WgqnRey5lP7g/fofzdKZhA5ww5N8Ch8mKJIN/Fo
rjiO9JRmPsu01egVCHmky5ogShjx9fFea6SR4gCG6H0QPpl7N4/BoD7vTkaCSC+W
Icpo6+s8fAHMrT7jABANP9JWo3gc+j5izyCS3/TYaY35QhOnlviwMx7zn8V1RoRy
hfmJ2DX7zWzg1Wp5fBPRNiolkC8oamVKHoTa4bbej7b8V5R8RDGW2MnnXyh6z0VU
O5qSMfwIPdAyyeE//CJWruDsvON7MUOcRa4UXNiEk7dTn0ANDlW3yAGA3whBUNJN
pxnWK+1a8z1h5t5Hyi/T3LY0W87mfwR9hIeWpfhTXvI4ERSahK1jtk3eYKRVXrkd
nSdmxFIggYca+wo8PxiPiKm6SzpM08xMg40ka0xNpdXSu396rpX49l8/ktX1506P
4K0L3fvVaAg4NEmr+69xQNomhS98AlVpyXwyGwoqEeoYfGkPNOsJjtuTT4waCSbS
EFLHsfRBiVfna95krEhK5MCTU4JUyNebQ1BIIqoplQle69OLf1pYpFLakiMmNZBe
DGIbq56RDwx5jO8D609OzSmYJ4uDg3CqD8K6+0P9Ucw5bAPCYPVof5N5Dmb4FQYG
bdVyxfGqUwXKHebC0u2MF8kLH420j6iHPrcgfDoj+w1rCW9X06nBuA5sYf9r4ESk
CuJEOBqZQi61Q1ZKu0amE3i3aBA1TOCftzG7JWNjbOMcSvuy4oL9jbKrLxkfoma5
OaWQeNWuhEBA6EamsBVIL5mIRsQv3Uj1TBDOjs4m54WKP5cKkVzp9zP71suQ1Y+E
mt2np3Wc3zwbkRH3kRjoS3saK0KBVD4x3EfmT/oZkLRM2RSCq98ONpDoSgr4nzZj
kYcOeWRnhrj1HUYsMyortx+y0V/4odG+UDs/3uTyC9pDRJaQ1TJG5zJX928FRsIt
ymVuwTKZx9X7PMqYcHD9SfxVEkJGM/bN1T/XFzasg9zhxtNjy1Sg3lEn6yRh0wLT
2enDLi2bnIglMR04LLc4KejE51lenu0hLIUuq6B5mBEoaS1TqIzzFoaXkzYBhtVG
EUpM0ak7+SOUf76UDfvch3CmsR1mzuOAab8zHHh7+gm8+vPOFCr8nJnnyFD2GbiJ
NuK8WxiywpMnpYvF3RFOYqsiQpVEjmlQ/RbjGGMwyQx0CwUnhPtxm+2IB3/2hp9B
FPr3BayD4tz6Pkn8lU9roifP9eMei76cf2r12vpxY1TlbvUNOqXusVO1HlXQMzrB
B6el3qT8ztuLyDqs1ath5xMDh71JJTvKeywrVma08URBm9kiqdsgSAEjFTBDSGl8
n0JhsA1vqqGKrF1oJw0JFu+EQkBQJUMva96T/6/5JsvBpI0rBZprk6wBD0+eVomq
wP9Xw5say8iXY+gBn+Sjp8Sr+VkMEJhL0YOOIK/Aeup7kBmhJyQDU0vjyo7GuiMz
VCrBECtVXPHmO/bkyS24ndOWFIpaR76be60hpQwOgq2p1CZauwuyVOZxmwaDFXLF
rb0ZhDFivCIF60hqSLCOnlbXvTd/t2Zk4qxRu3WbIZjXTdiI9UhnRLMzWjL59WTV
wDB+cJJza6MQqM66WYuzO1dHPmDbw/TFGEh6mf8G3fh4LwI1h4ZJoPnJUqVWyXfJ
u4BHROZyu6BSAYjZ4JQaaGG5owz0pxZjGr0uuaXW1FOyQpzqpxN3HB5m/9gfjJjI
ysALqxHiMaLhBruO8Pze63/Af3SwL1rDiftDb9WTIAXmvQCsTTDIRpOZGjAWPCiW
Nz8edMsLDXKBrBcIgz0izYSkWm+t++Si7c18lSaROc2R928kMyk5JsOIvyPUFOjc
5l5OAaVAmwiDqxWlLwZXxxBrqq+zYPcZpiUiYZmtQC87hPBhA3ih0cuYdeqMlblG
MUcNEfLhHnlVMZLFop8N3UqdfPOLXyvfuZe3WUXxHgLga0RjZMfJvdOgpYrn4VEM
GBKZD1sSuDq473jcBvuhSDbvJi+kjYNh2sYYRHFJBziNndBKXzNjeS+Lcxe6Th0s
LS6LKdA7P2g1v0INF9WJyRZcAeMJ5CuxYsCziZu362639ZkG1moHaJmQn+nCkrTg
46gxhAqaNhHCkb7MuWI8PmTc2a2CPPETqx9mJIR8XfmFqYQeDVYOX67GTxgQLR4D
lBiH290mhVhScAmsMcTO0lsmUhZ6x2Obhwo5OhrmVNiieeBJNnlbmQICUo3u8ZKI
AIi1IceM7oYzpscse7gEWYczAAaQGs+P0BMkd1cISq5U4E5RYzpsZAzo5ppIZaqa
72HIeaoCTj5efY2Smc7VxwzETYV7XoOcyWDyxV+1i3X287rI+ZsIIvyfYvCyQubN
eVR0fFx1JQgQV1fLlKZqwhkEi7oaxiKBH92/9dpHbcsOHMaJZrAp2DRqAbcbQoOH
sPesS3qbnoeo4CPsY3KFlNJLHMYE0XrHScSl29zTx6IXJVZZmR0AHx2rGuiOlU6E
I3PW8enRGIiZ+SvMXx33gA7NBVGUnkVPCmtq4E1uE2IGwsYUPj2vFkru+ONZyVEZ
5Nm1saJPEqGcbu3BXj2GqaKSbnDOWMOIlaVMiQU+yUGguF8QS9DOdZ0ShhUgE8mF
iANQ9jwiRPnJ1RzPkzhUg40jW5kvSRot7p6vladTFDbEAJT73V0Nc1/8qs5paXXY
hq6tEwemFIMU6m8cG7rpd7mTvui9dqZG4kNgnmr+tlO6glYfNwNPlRlJWursKuav
1EwDgIAPTqgw74ykGKf7Uoooe7vbHYn85ySAJYO2aFSe5UEfTAujI8rY3U2r8kg5
deKIEqZ1H+hA+rXWlTk4AwKgxU4vvW8FiSQirD69LlHaw8CQ2aFONSm5JhE9d1T4
un2KMxPAIw6Wv3KzMQCHpM1u/icGJHkIV62HRUWzGH9pZ7vomvf1qb72l2T7qGer
gqCqgw3zd+XlYFTWZgS8YpdP10+QqJnbS+rSai+VyDOkR+8oVvO66x9VP/LR0M6m
2w6b8x5frO+AgTidVzaoS3IgFWxPCPKPnWtVr8LKPzQru17lrG6t10RpHN+2vRLB
K5227fJFOFsAvtnHe+mxpfHoktvyy5B+jPU6I/4ktw9sM0Up/kO1A+W8JM8XyxJa
qEBoqnkHJyRuFc7A7Q26UycwyZHDP5vSPiaDNIOQbcElum9ZBNF9hoBgxyNwKuaL
BSucGmhnLIjhUhUq8bOv30ZTuP1FUjTaWFdvO08hm02L06zsibE6Nw7vKMBQh4qJ
TBcI24WTdFATXAyBUc8OxaS4DZ1ZlW7fcFbakAkVLkpV9San4OX/2f7ZZN9URnY4
jDzUYGTkO45xyQjdjl5GVNPuyrqaJ1PDUFgtP3fkkEgXSDRaBfSB+IZsu5ULeuss
Tj+xOPJk5AW3Ovvx9Pnoy6gda7thXVHUYQZdHKq9gUvco95P0rvULdCmXSgMb/ls
P0z49oIxUQ5S2r2myobZv+0oEltJ8McPBQu90IJoNkpvIzP+3cq3qNc3eh9ZEf52
x66VSYDct0vmzLozSAN3WJ3RTNrPrvznnLYyCj3lpCgFhIzduEgBc8vVBw8A8MZT
h9CA9JWX9FkdMR2FDK6YYvuU+hHv/V+Uripqn9rfz9rO1T0t108rPEoI8pDpl3HJ
+S6SFduLEvSx4oBMKLzEdnKKo2we8Adg1/l0Lfwr9v1EGpujXh1GHKBcH4w5Jzeu
ETbUlcdjRzVFwuoztrv4FZZ7wt98KcfdYYr5XbFFez4CFtaBm8aGNoi9jDQucMU8
ZhJ/QsSM19GtUo1Aauk622MhTvfvQhjS/zBDvUXIynr3Gfv1beJdxHFkgS9hqbd2
kUqnS48FG5t0Oi/GO0lckFl3ELeEoHJuR8PTLXjpYFGn+UvTEmQfLNPc7zPRe5tQ
Uu/yhpiVtr3ULW3Pq6t50DtO4bFNpxON/dYEj2nsU22AcP2jdixoOV+YfjmdfRL6
fVon7KDPgEOkQ2BYJHGRFHDdi1zD1oVBOQUWgswsNQz6dUX9rIu4eOXvP5ow3LtE
C0CT6Jw7j64aa1Wo1kTo2Lc5SB42FbptYUo2f/XkFevziuwIWDREPV0mYrJB9dVh
dGmUm1pZTbL3XTS2/ECvac8ukhxiAeVemKEQMj3Gmm/FMVqZMLYW82xr2IhnOgUO
jHtoc7GHl+IcgOveTSUrTDhCDBOQatmfPP8rseKKq97JtnYiUqIUAl//AAK+KzyP
gU7MaKJWPZgHBC7n8Mdf6SIyJGwVEjFDjgMjv64BYOgsuMQd8xVWZ0jU2LHRzcyD
a9OTF7w/kHAZWFPUHXejDiGcybUNFgwLM7ouy+bGqcvk1VBQMEvxzHBHu3sYizaC
52NVuqD+uTIja3EdH48s9XuVQZ9/GgE/Xhp7WN4w1BQnWwcvq/ajLGgLfoK53YFL
JkqOMrLCuZoCkUSymet9LAGXSkm3JpFt2Ya8lX6AvOWjw63dH5mIYh3MNGQloFHe
Ecvf8nLF4WEqIsFCqD6zu+XUmcpEU7QhbkFA5K2SvImNEdRPGWwjKVypbQdSZAwe
JLbbAzQRhYHwKZfPfIXKCTpVZzSNCqHRTWS3fwddtU8al4oIM/7CYWCetSxDpn2H
w5x9HCs6oEmu5oATbTS1xpFAa5oArrv7yt6qzJ+b79T3hEEJAsr+u7wXANosdXaA
n7In0TxvNeTqr+4yCeB5xpJjjHF/ix7pjypXXNAfvZCVhm8/XcUL6bSn8HuJNxGl
fTLKaMaPK/syjFAptZ12p9RJ3kHPhE48dGB60FweN/mBBkmxPvDmXFG/bMfN6o61
klQTEVkisRAWwLTWtlPlXk1mZ6e5bY9zHXJzONO8wBie6BpiGRd+SZ6SKXhLO7sp
sTwzcLQbMOAdC7CjkjYDQDrMI4bpG5hAtOMeyqIP2Pkf7OYO7RC4TaDM+kFLn0mc
wzVRLNPQQLHrbBJIfIo71R4nDIw7Kxjs2f9DyyS8L4NLRJTe7U1PhlTaArTZO69s
mqu1U1hRyde8IWXP5Mme9glhaYHJTGKeAjmCKWbzjIWzRnfAEAHypbQMjPHCMthy
aXS38UiwUcdO5pIsQGqdCZbGjmxaZuL201t5ZlxpMKx+vWymKHme88tn4YTyqFpt
B/nGie1qfUtusRbz+N2NWjrdsCRnkoQaHPbb3TulH3R3RhkikJtUjJ9YaVTolKQR
bgzAN8KWDvFzu4Kvp7RffsCQSApkjzYVr/fZxWwVu+4QVVcV+wCUerrG1yJ+aYa6
zTztEfQVl4Ah21xSn5ucDFmhtL5G0s2vRt5VaFc/aFxDab7OqgxZ/D2C1rhJK6p3
lXGI92pZNiUZUNmLdJeuZTlSqkeyQJAkB7XT9OsidnTfc6I3oIBwTm4915XCd6F0
FWSkXD/OFFhzvylfwVML/Ku70FF91txPEGQgHgizLWfKXh+DonvZOZoXqQkDOqx3
uSEDTv1CN38vzjXaHZ5LIbFcEtIOI3O2AdoLfiqB88OMkyWtD0cuL2DvPaWoBr4Q
EMH9omx9EPM/MHNfvAVILbyP6nLO54QK0281dDu+eLSFqVqgygAyRocsbeZIjxL4
leMT+aP0GAIKO3mARcdeafvcDLZdNMn/anw8rz+a51k7OosJDru/W8lN7C0OieUe
f0Dzlej8ERFG2n7pvjfaxOxeh7hF2IzIwmiIMEgOaW7+QM2CuSu0TIXGroeAm97f
6nhwp7YDQ7GI55MQr7AZcDVSKJgrGNpCMi2SQiB4OoJb2wJDm22cJ0Z48sgIC8N1
SAGd2N2BP9sFmDNscmdsJwJo1l71hjsHgzGtmbcosqB/X3FcGvOcmwDOtwToh8oT
qZz7ip56ozCiuH6u2GL/UR6ISg6Yfn2okFTkxikbOUWF4FDkSQ1Ic45De0H9Ps+0
013RG1naT4EteOaNnj4lInsIwsMZHfGHz0Gg+uMWwbja1Pb+Dhuw6VcqxiqtvR+i
kJ2rDLX2xfKIYqvOMAXR5v2zpujVas6z99x2nnomIf/1nKHolzF256b6zOoPnmnA
Bkyurb14SMUVanBd7LM2tg1xSLJNE+z96mqyNFII1aDid4u0DKeJV+4ZucRjZvXk
uSu0GiHQHk5jCOhXCSs9ZI5EQHcXpaIqR0RKphrpIycrjmpcRT6I3w3Ge/+xvXuj
6N5h95QHr4O9Nery0tlL1TJtqAhcF563hj1QRC2pDkCdS9yD3jRxbkAVMwFAao7/
BJttGdSVqsf9lFD9ZeXiO4kTQaDakAgsulIP6PeJ6kqpcDC7WAZKyHfsQ+fSMTM4
SaCOOuyoctfK3FYrR7A4QjzONjb92b8xRuZY4rXjgOFH9fv3uT3n+cW+NOlKnJvP
K2WJsAPasGDppmVnkMLqa0zSWYOFRjH5XZjGdclCbJCDQVCn2kYa1lanU7+kE8B1
FkjmusezEQO8qARp+2tOPeH7f4UE2hJJRXJNj0r0fEnQKKatUTz80IblBSJCjCV0
WYrubRDCTtKGzwGNEwQKdc7WGkIMXtrbUQjtV4LpyawDD47DKxlSDc6UTaDsfC+Q
9l0L0/LP9ozqc2PYJY5ic1kWw8cDScMSpZYg+RZbGotUWaY5JgEjr3ROC3Gxsthg
5p2kGfabeoyp1RX3LMZei2rYmFmPOOrDt2tE6smo8qjN+DCtj5nkyvEmGtAh2mmZ
GTDsasX28nSFDrwn2nrlBDmnhryORmhYG9FJfw8TWwf15IMqXhpeVdeeBFqdY1f0
M4qmAE/npraXDMDEQjUI/0raie5f/aD3hhBreKIE6b9/iX3XqG8x/2ZoV2I/Tfny
6JeZiYgIqmKD85wAF3QsBpym5AIejCluUDAE7NfL5nrJic9JjaPsphtc4aCqDT5S
x5/DQRe1Mxw90b8pUrBNo60IuTJbBbNd4jwWzbRqBv6sXrh0vdQHFwyuhMmXw5yF
ytTcGxxNVjcTFIKw+cED77eQUVDOA01dcRRlzNBDp5qIWfCVfLvS/d47zN7vgPU3
jb4BMgNGv6xNpf37FHJFlHH63Z4NmDLLRptfIgiEQA6kgTjcPjn3CMY4JdHAtLEW
ltd8+jZP9xpSNtvzS3BJ6EaSguLX+NvOv1YpxPJ2CUPhDVK38Hbkqvx+msVioiCA
N60/l2Ub4yPrxEzH7g6K3tRjZJjfbdhN9g+XLrUJiWgBlihphF6ypUmnsxZG4Aze
roupGX5uw0p0ff55ypsUH8ky26lV5n1XVtGxOtPn6WZAj0jBZHYcOQRqzVf8yO76
ABk7Xa4QWDSrrlZa3HdxK0jXUa6ohqSiEKd0a8I8VeVrr38ojMAE68cK4/zEP70H
g+DHQZU4bxAkQzJTgg3Bf2DyyRjFEmIFhZpi3M4dVCJ6eTzqUgh4LXakY5ClcXKM
eDvqGa+CDSiVemk88JfoVHPSMaGL1TrQPDqI4BLKj00NlcQ+PO7Fw5FusVBabpXL
Mkzjj2ckh/VHc1dRuV0oTJnkTEtCszatRUhxfNCPwB7r/B+/HZno8XPHHLxnErA2
YxhLNQxb2NenkR7YwQvZc5yraa6Wi6Kg7Se0w4vFzLG6IsBx2OQAp66lP+bvsrl3
/3ddYvXRcAeUhHhcRs5d0YkCre5LRlIEzYaj4BwGokII6g3zhGFg17TP59Up/Yq0
AaPIaG5tJg2vy+4AReR4sc/LXM5/Y6gDYgE+yB9V9UWwe3kHIDQ+6iNGcpNLm1jZ
PtirvWK2spURzlEbSCG4uzOkwKpdaSeqaTaX+8UqJdu2Lhd28zjFtNcBTb9EgR9V
+mktZHhNNeeav5Hz2EUV245ys6g2bppUWnx9rAlY2aLViK/nLLFCjdML8TlwzeVD
A9NlgXxOlpdfuBlYVjhEJc1gHeqodme69SJaXs4BsErdB4Tf/Q8upAlUyU40haKn
PrpHK+2ro7/8SGNQh0pslfVnaneIW1URpSLAiQb7rsmkZP2vzdvLmal+EgJ5NbUD
kOSuELqZ5AEahKYm9R3Y8dn2s9frUdKsPL8YYhwucDc9Wp+0jKyHeWdosxdV6hf/
PXzGQQdNUCY3kO40Ank6rBPHg+BmXs2Elw0FYnX80xz3HuQLuVFgWsl3My49Fupr
USL6qvTd02dipYQPsqo3kTmgTuQi9sf89oTctU1hlVXtYkUIna3jtRV9UfPFbkvk
Yo5R6p5iaTbCL9Ysj4aWeiAQdY4QEtrAEsO9Exu09Zo+bC1wRqlYGV9mUlJ3o6jb
yYJM7NHqLcXaZH0KJ4YucMIHxgWrB2VtDR4r7jEFnrEx/hMpEM1CBzSGusT3uFfx
p+JnVx1rDwvawDdM4XuOUHeKhQw5/R5dEy1OwFa8LIymc8V7qK2wO28dAdx+mAGQ
0NwQwczz3FG/wG6fih8ZGgNT3uuh+Do2k5CstY+eIkQ04iqHgl2Tm3Ee1W49x6fI
wMnR3b16DvuOLrAT6nuRSI1seFxbaHV6jgFfJyGfJFZfLkW3+R34d6clWHLXX7NO
bK6W7XbqKxXfMj0o5gHCbDY2y5s4B0+d1KhbG95/OzpH0zc6t3ZUXETHLrSITBFS
r2wGiGucAtyBINL9QBptdsgPnEhhWQQNy4vFwIeluBHhj23BKnOD2fsn5KmRshkf
HR4eIfTeNhMUlS6MgMqJ89sJIu+RbqQQOXXZB944U69OxDqcu7XSicxBOCk+K8K8
S/brSh0dxvvfXlMnewDzdKkN1z5HY2FTGOAq7ptZvur2i6FD4N2APIVm70W093Db
srGGOUdKySGz1ehVQKXbIFLLKldSE9XMA/EsjX6A5u6VE9e0NdAkSD66UDCphDW6
c5e9zOgREzGVgKMrX/Uw8Pt2bhcnT+wpSixhlLk99nJ7oTxBW8DRj4dz02cMFljq
Bp5wNeucBNewJoakjy6MKOgttiIa1IUmVuQ+Q8P4WwzNKCWz0Z1j6bKwHAlvuZQR
Vz0vIx667xFYodsH2un4rjHskKlcX6WAi1BbMXRcmK2/c/xk3DcB255niOoUa4oB
awoS4Nek/m8kMcs+Z6uBfG19+kKQ1NEv7mmWbAT6GvYeybIUVOF3asW8t4h37y5e
1QtCWZUJ+I8ZGBFss2YPlFPU1/HI9i02qNyUvOyQPwCnxouvWdshQGeGBQox40lT
7EgdwKWYot55CzFNep2f+lH4Fdq6Cn7zdvoIsnsBcxT1MvUuOw4C3OEZ1Bsk+YkZ
1q3vtUtGpA/ZOGdEN7IWgsLIOHCXDiCu6ltgPGX8UGQCme4qO0ixxQrIiC6UZwJP
5F8dzC615qMFQ+BqUuQUFW/hn5Opfp0iUtyQcR0g7z59uTU2qLviZNn4sHrjl0Go
MD8nWSp3yTCPmrbSUK2Pd43/HLxd6ugRG/brPob0iuMb+IX5CJN3SnsEkgrBaMDu
V/gD8/jVlmRmWzwnvO1ckjU5BC8oiflLN0JQ+WRc7ipGn+LAlnp4vpJhGYb71iDR
w38i4TFwswQRFRjXCcAvkPY8rOzHC6o6owb/3daCtZOTggrK3kteHQgQWmGU4iRU
QsTkx/ve/664weI0SNMJHX1knIPunYP8whbKGS+5atFhl/dOnz4tJ8TCYzC/Nj2z
8bF028iVvcwr1h9mUa2r5MJV9cknmo54z8Ukectt+Ih30VjCQPTASiMFs1rsSUW6
xFLPHxsUKG2iepzqyxGKGCldfWL5FKkBdpCpmwK2NrI4yMhGiDijTtcaGLspusXx
heIVDmEXpoSJl26/QEC+Tl7zr8U0U8+CD43MKVltVLIh5usOm6hL5SjZxNmDhh4r
xR1pvWTOdnoHoCk5h0/+wV2OCp9Cl5pPla/2SG726XqwtrZEKvZzy2g3URG41Cub
ti9usbUjpvUheHpUOKCbQH27ZwbfKgVN9Kn2virVRhhOu9qR8mpuljOZFNmJnRUh
6OWJ1UZWgLjEHss0bBFeRWnAUWHosLsMfG/ibwLfv03wUYHsRfJMw5U59NEz9aUM
7Z2hct1LUR+TGbHmx+9vamud7i8y36PXz80b3D9O8sPtSEycYU+wOcWKqGyza+E1
UN4qxIsAkpNQ9BsxXMa/8DIQpgYSKfFcCEi2nek9vVzXIWKPkjeyP6x1a4I+QEPg
wvYkKNOnmlV2TvUYcbVxo+alR0WedBfWsgMMB2rwuBgMb+RsbKHQ+/H0lk2zn0iV
D/RaxnI/ebw/DWEyJJ6qmEu5vDFwaJXFXYtnraeOXliaanezlxjf84MVheLkdj/t
owv4CVJQw8k/exmhK/lFIQkWuJ+GrLJA0IEyeWIxbYypbSZG/uWwWMkySnMKk5uE
KOFO6DWXGQ1yfeEBSHlzbLzLhHkeHGRO1f6A/WRAwJRrrBTzgUP4LLsKz8fUC9tZ
jJhaQtIF3kqGOVOmaMBG317EGZys+2oNNiH1DajJC58vjCFl0Lo1viz1KJviFSpB
XqsvIbNA/Fnq0l1v+291h1aNXtsGl7pGVY5r3xPOhDPRFm+takdKRyGJp6mx8oB4
Z856pUKDU7zh+mNNHNGx+BA8C9aEIwYqOWxFoWOzqiMfYZLEHJ0cq630axxMLj1J
8lnrDbJjLnuVrXTdSMHXtWMhvtLnmZTC9SnB6tQD8laCgQMEfPWL95KPfGfUX91P
waAxalovLYcZCUOHoAQlCarN+cZHx+MKiz2bLdk+Qxtkun4MGwxpNR0qvNDszcbM
mqbtM/fNYP+A4t4FRO0rzqUHv5fOOhA6Y69qEF1MSghrl6X2UJvpX5SCUDy4Oc9n
yJGK/Gf2OmRlHim+GzGu4sF9MI1kYM3KDax7pX2hSejJLl7UTQReiICSdCA7gR7A
TtBFEZZhwiNpxt8BITtK/EPNp/7fCDg1shf5AhVfj2qGWLTPVbs1ExAzKF0B4cuu
F38z49pCMGAS6ozolbW6NTp6Sh/7O7l85pMTMvbE0xNnk21z/yIptYgbSi4lrQSc
+SLdTp7+eo2fVODrwNyTA1XTvzyG+MCxCewVURlCHWiPPpuxpZwGmVG+iHuTtGSc
2fEktRC3LC7ydD1vIkmdYBzpKC5fjl2Z8na2DoMSwFsZp7VXxQXcPPibh9gc2GCG
QpaZGVGnllSjLWcpdkW9FyBPIhc53zjX04vEnlusOMwcCRHFBot5pEjoX4Ntz1Z0
95Wb+qUxFjo1vhgoMiZS4JvEhIBMiaZYtf0/ZHaz8JigRDM/iBpNjDln+jbzSHHQ
q+7jtEt5gLGDe3JvCpS2enwujJKv3Ibo0HE/wtpph/eSfFpzcnkEbF2+x53OP3eX
EaSIU3WXYR59TePC13N8DhBxX0WXCb3C8nA+Xgi958Z6k7FpqV2SYtsdrsvambY0
N762RS3GRFo7HF/5JhCq6lkZrgmoS4vPSy6MUaDK49MG1Hr5azNTft/TDhJkGhW2
GvxKxp3rGLbyC2zg0RFUhRwzXOU4pYMFWd+k2ky9YpExN1Vy14V1jsf6ZwszJsic
GDuCAVxV5rRW3/bQu/DPb0HnVq6EwDUtMFYnSAZd/TidqzE3B1k2moZ/SUhKSzZa
7YuZMb/k1eCVd3EKY7PEdusBYMRwZNlZYwKLQvCrEwXlr4kp+VS0Zi3YLEKlxXKN
tQMKgyUte6Fo/BLkz0Ee03RFWngi7sqHOHrZIdU0y5rS/UkhT0IsEKpC/b2A+bwF
4HLENKPDT0LAvDTGpun/uhsa6nPgBcr8zYLryKC6VCFSlwIEw6LOGPHHZR7jP2tZ
wMcRl1dggxGU5whX5p4iOAEv0sjEUR0v2b1vL9m51AyaLYoKe978IJ+ekMKS15iK
VN5arZpNrNyZTSYMMQ25TTokM8+ACPa7HlzdxbXW4+a6l29VFQsh0whntAv/+Lsx
FcmlZPrRGgI8SKsLJUoCqxxcIx3e20rluzOkzskrgzLnrJoDuYzhUxdOmTrnqyKD
yfcv2fiMN9gBUscJi3KvaAjQ/kyw5P9iblpJ8z9u57P1vf7YqPyIhjXxWwndCHx5
UR7uQN0o1dIkO4IDvwsdVgO/mZGIcKeU16at8Eoqb4whsPPZzi0bfuS7KvlvUd+L
wrBo7wqyzSO3UG+IfPzXFo5oXo9gRVX+Xb3QQlW21gXAlZLM/RhuE169E+eRO5Wo
KZWloFCPvhXAk4ItrYC8YWm3WC86cteerlx5aeKSmu8VJbE/YUeNlADzIRm787qU
VLDIfuNDKUBsJ/GU3Lgj9sKP2svH/CYj5qr3yu9G8YW0DFmjuFo6HdDOdz3pKQDX
4baRRgxRB9gaFkACtHdmnnQGtKRCp8ByN72jCbhcDA3LbIqmKcPlOouqx495tU6M
dI7uBmVCnm8KsDwk/lvgFtygg2f3KExqrRbSFjr0EJhbY9OO4rxXh38ioUcVUqne
2ZPcKKksTE6K87f2bAdI1YYQNLMAVG9ISaczAkqQuH07H5z1NQ7POOXh5I5rHEuq
EgRNm1RkYIjvTxL0It3P5jvdwHrYz8y+uTZ1INEh+qpzXSI20F744zG410BXWaoU
EMo7PvPbCBgVkKLQJZTObs3pEDA+iL9LKth3Qb4cpMm2V/84n5V8FzmyAMXUWLrD
TwUOt/fR4KJG+xAarV410sO675ieO00HdvESpwV6rm5LGEVWQvBTZNofr6nI5/Fk
GhsBySwvkHySNMbwJynVg9wBCiI6iUxdSVfDSu40nRKb+Av13PWVQ4SybhtSm1NS
eIIrsJmb7pCRNAuajKIxJyxtBm5wB4YvA52W0aU356u6z2N6sEphnVip5nhOacAY
DJJbbVl3LaCBitQLlVT6ZQ6xCG//7u3/cZLUgqL3K1tMYe/SXkB07T69jkUwW+tA
+DZO8SwX7RYXpu8Ay8KVU6bsW5Nve+XtPjTUj/tj1T9JWnURHf/mCI4FcbmHO3nJ
Jw+ODJm4LNSh8tvxCeOFh75I96yhHmv61a0VnpAAiX203jJVVeSUo0Vit5KbBc3H
tfZ+Jwc09UB2v5qcf6bi0M73UpyGn1QOeZo+TQDuxIwu/XjT06EesIYVAiVlRaVT
vF0Bfl2pjGw2BvaEllpHnRzfl6CY3n3TR8y41nRvV0jfJ/KAyVRkLZrkOInhPGu9
hYLTKhVywQftsgAXQnBoMFNhjXMDCEFlWMqFHsOlrjXvb0fe6PyMAbeG2MkLp601
5NrDVya/EuFIwy/rB3GX2BOHRe3Psz4i1Py+Qqz5XvTNtBXy8ghUeR2SEZHDihW6
mTl7lUeqhss0IHNp934JgBoX9DNSnnQcWATJiGN/pzDy2R1m8COXnzNiWiQguntO
fLfr88FvcMgmfElwLdrJyJ3LhHWENF6HdQY9yfCGbwk4ZGBaXIzgg7UbwRpP6y2P
9fqgviB8/LFhzmkC683GUH9e5ZZSfuxZJACgHnxY7SO+Elrr2pmSflJRrUVHR06F
UgAxm+6ym+1plgOL0LAyMNSnbJEvFv3nYOCHUQZyImfr52H/k/4PyeNBRtHhU2UK
uEzZsUTvA83Edg32ggwdUCi2gn9Sy18zyh8OidLFROk54o+4x/1ZJq+7N8Crc1bU
fcQ6LrnN6qqjVcqTRMr29VxzJ4ChZsbfF7CA/cUqRMCIF8f+v1OUslUAHQuvX0Gf
PP3fZAtAYfWWIvkAeIDbMNr4zwVyvRP3iDgmX0cZ93mTK+LZhrQYQpm30yiQgjEy
6hC9YpW2gO0yRaIYzyakFNBKsCInnlaOX5DlpEPLijtcAa2Ao+05Oh8y0UJX9Joa
qbm8IBpVjONQSFiXVK84/e3jRivM+eM0uJ/gBdS+oDeQ+Vsv6BeSR9FNh/zyQnY4
4Jp+2P/+3UsgaF+Dy7BRkvipdQjyAtqVUimP02VaeIKFDVXRc5mb3j9k/3Gw3b+O
MBhl2o1Ap9TqiVY92WgaJYC2578qhmfgORapdxjAoVVyp4TpM3AZvpcW1QcN1jLm
evg3zhAAS6eErFKhEIU4MWA57GHGau7zX2IE9VU+onfjummUsXyafRc93gcaZnkj
Zu0ojwW42RrqXsqPTCcNrHXT/isxNfnhMjPn5dwvhabpC2vdSpeJ/BUnmQ145X5d
oxOnaJiDVLBA0pE5JcM3X3+4m7OoCi2pqzRBS7hg3dh79zzlO6eRMOowUOg3QK9/
Rtur29zH9PJD1UyDqZM66ge/ctnBiL5+4aCJoO/H7pjyQjKGiCYrCu+D1AOQ7on7
FfaGs6S4Rv1RrCevjUNnuhGCEecx5VzhSbnewQZLN16KgNhB8aKEB92a5zrjC2js
nM8PKNE/qAJ4ZhekQtflokGewYRuB7AVysNNWshTNQ+oLJxNxsvS9iGThoogyyY+
Ari1H/v7Ilx++nTJDU2/Xo7v+IU/+weR89Fv+tO1WQO6LBAt5Peq+68pmiB1guzj
/pvBGiqyd2Lb3M5WqqLKtVZij4rjvwraaMqiezCP7oNI3kM0OfrbKP8eAa3HVGCb
KvNOWLTPSQxWlHrYRzlqz3jNGv2MNi+PV/nA+XCioVOBEACvA7RHENr6Li0QpnkQ
M6YIWhmMvtNiSHkdHBNcYgKuLvaavyhYVx3d8wYB8LFpN4lYjSRdDRthAeaJU0Ei
NvZmXOjKDJkVwH/OuQIDJ3+lUmuLK5rEQfrlAt9rh62fRwhAo7nJzuJeoZO+Gt4O
8v9lF/7oWd//LbqqDHidR9RTifpF4b0PFkzAlZC/Od9kSZ/pGnVmYTvZuUPU1e0F
5U7f6ZsOAEMnK2iEa2bavwb0HQekAOCiw452MUaPDj1CFV7qO5+eIyH+a+bcnrx2
+3L5Dljnua2Ibc/fPFyKZJeqoQohZuY74n+zkrJ1QsfDOShyF6Sbcab7Vz0MU9k+
1gkggQkKwm3uzErAyR08MBJA4IYifdFrONNkL+tQUiYLWWEmO+NP2mmlswB72xL7
aIfbDIC8tqAfl5uhE1E9DIlC+vDP+TjY+UZ1FWcqq2lQIbiPrdv4VCmTLgp3ts+e
v+X+umilKPYAqIlKRyt8zEBdJq4ycHysPuz9yT7V4VWwhZVZV13825/JO7xsHfI2
2D2qJkuuR32DiG26DpAj0vVxTt5X1tB7ymZvSF18KG5cZJprgglBONdG9K/BYOBM
H02DWyj6dRCzz0zDXIkaFE4MaJcsj8/ASOJmtzTyqxtXbonWFmEF4TMUcn7ktnu4
JYsUKBqyKtOvfOYFj4R3scfuFyme4XoHkVGZWpH+Vi1T7AliuX6a8vc5qAFBuqSK
nRb3eW7bk5BDp9Fi+YO4ubUk0iG/fEQWy9eARWd1e7D+jUFx9lztWrS1z2O2jkY9
M/GjMcCrHm5Aj3OpOr2bELQQvemfQK7a2YgkPLjYq9MQJopZ8zTDjgk8d1/UGMgK
9Y2ZUkhtuenyJ6Y5DmCRQBr5TJPj0g2d/fUiKmTFWQ9YS81EO5ilTvgDoI58epzG
2WULdbCpRb4xyOjLOOyIIs6d9BKKW72m43asUowpmk+BBCR6upvv39Shb3hXlckZ
K5bfafsUFbR8fFRgdJC/IQZPsh0d6T/6IZqgu1w9r31PcbTJW+2cjuQhqYZwMYMW
ruO+DmBy0vWXsEzc5XxWN9iBYc4JROiFhhLWiRDbYTXUNA3CNzDGhly7M5VSSsPa
nN867LVy8HjXXjQ3T3tk7JlL+7HO0jdsoOkl3JCz3K2450qdsl1thIMb5KyXYufE
5+OP/HQe43NPsMKO+tvAe88HD1gqKK0dBnHYuSEOO8GteglbHziwFLYr9QeH9MRe
8dhMkoiCpdJ4OuWsGt9HYlZoiiaF5vmHz0reg212LLANO80zxSMNUYMrFuD2vEVy
DEase73P2BcLTi/D6JTf1lE7kIc8GWgROJULxFlsvH89ohMx73al94AKATB+ntxR
yy6w0vLQlHsPwEZlKuSaxV5YoV2S4KIFW4c6MRuquFT6quScBWYbfFVgCnP12Sa4
/vmrAKx+ZbAi+8BGh5nRmWz+3F86Y43XU2Yob/kT/esq9cTKXYge0PW9r9zBIZHb
dxpTJLMhq486u4No1JlIaeYqTIUYATNDB6Zg7N8eaW0kJM+4Nnr3e53hRZEUmcBg
xrS0+O1JmsBCgbRG3Z56i7asDjqVZvgfafDq7HBmZX6NyYhPt598Pd1W7RGW+iZw
6c4bJq2KyJaoRu26+L09Foi/lptwAKy/JnEuRjGdH4B0KP0nCBv7bSSAeLdL31/s
2ZJ89W1EMqlcdstNsPpldFXVRAaiR96iaayRA/hB6dtMgXym1f+bOKoS+RTHG98Z
FLlgtNalNSxMW+YN+5KrmLd4rhVoWWnc0eu/MvEy+TyuOJsV7UQFvcxjmTrwd0iW
2S+5GT8EGE5wFfgvh1u77GxmsD857HzYQ/qFhAdsTfSLW8fqdv1XmxB6WJ4qLaPw
0hEzfcI9rKud5KzW4+kL55IiUtFhSCkmddqeFrk8YRXORvOXEspT9by6iXmbl5p4
boC3ZqD7NlCnglTYhxpA6rwX6A6OM1oYsvNqwN9rQZPPhAIBJvQiY022GSHnEWoE
sSCeBJBfLjgyuPW7QrcI6cqC2QCdcgx3RROGkeY2ZCI34cq8vZq/TxWgXEAsF5vQ
RLkUQV9q7GElCqii9d81B23Mm3mqvXvXK/KiSZZuj4H3x1KBf3SbiEwDBSmZb8D7
6S7FBpSA2+Z1qAPowHUVJyb7oCBLMzYckAUI1ZNuUDsepE6Mzuz5Zqf//PQsxeDu
py0aOKlABcJJjPc0bEfX8lSK02Ns06dTal0Sigom4FP4C2BzCLFYPPQUf5jL+MnZ
aD3xkAoA/86HZ7ybeYd7vTVneghjTqelrUnkThd8C3kv6BVixCbSYYgL2Ihe38gV
h8LyNleJdc2Y5OSIMLaf9U1cp6DOcOAjGu+olEfa9xqH6M68Cd32pBlDRZCTEkKI
sPENkS1exOLts6LAvgJhujwl8qyKyZEsXUt5Rha4bJ5EI8YeCC8cAjB4idG8V8fp
oo5j6j4I3p1EyNNr2IS//kT5sGoDPMgz5XGehMBMbJjMg8DtdOaxhQQIyEM70Kt/
Ou1q2JAJEUsNAWY+rurMKSmvzNCzh/kv6d1Z6pF3Mt3IiM1FutKB2maJ6dJ8RNFe
Q4dolc55jk5ez7Suatha889D0vYGbugXmMMoWHeGU9em2rRTFk+2OrzjWVgJlA+J
3+US4I6+7ANU65ud477yoLTsaOHyBcsMu/iim4FP6i9uXpSBcWt/RnnecJ7t929g
Ea45JvhrX/47QXrk+uS4B+WPzCgXdvkVNp1VjV3RYALVjamFYQ3rM3sG6/2CtOKd
i8boOuEjLcR8jLdwxsU5ACMwO+9IK/dqoGii92HGr72Rr90fBPjlAUw1J9sgftnT
P2SVdu4/I8hyNXN7ljo5NVcCUjcs4E4Iah4uVMtlkVUN6+/Fr8jSmZ3DzNShnVOi
WjhsJc1yjFD5OeqpaEhGt28XYemBrnLkZnRNhYPpA3GneUreiZN2WeyqlA9fks7K
RRfP9p55CzoUdIylPEKlXFy5Tt8gkPOmKfOlLsc10d7lTWvIlQG2A0tiieQ04zR7
yrZJWMlq3r8Y5HDoGo5/sY9DEHz863bUI3ZZBfvxgSI0RoGAz6b1RMlQuD+3QK/6
BXKlAcItvdVak+fGqgMD82M4XQCLkV/aKKwniL+bz/22KStE1aPpIL7XSLZWnI+U
25+hxaau/eUXKh/93VhGeC5T1ae1cDvoOf5HrYw11CnKTs6Oux/l6TmivcDzj65c
v/MJzECWiNQBOfZMzq5kWdK1puRS6tZnyLPeT+I1JqOFFHkA/oc+5o/91OlS9gEh
TUURzUs0awsNu3XUe2vEsA14DdcpT7YgykbApQ+TZLjZLIKRImXIcCkGN/WVCxhZ
4EJV4Rvsz9Qrrjyp1pRNCUAPpZvIh0a2FzPVVTUfsDTSEK4efouJLq1N6zX5XZpG
Kvfa8MYq84bTKFLw0i7A75s6hOROUTpVKlpyTR3BdF0EskEUc7sGg9Sgs7cJbC2n
ykJOGqu/dTfBBw2mBWButM+naoE+yZe5JkRIOK2Q6uscSjmt31UOYYmtKB9VILHW
P468aLQWT3GW/B5hFjRrk6Mbu+8JfqZnY02HEnf9jAR8D+p03ZbB//5pBrTEoElV
vGvl/Aph8HdM1QvL9TYyh7Z5nHa1RZXFsHH+XVArJDqfstoWimCQGOQmf87pZkdj
kmDsVqYHbNwsR+aeOsXprKVwQ92w8Uf0RpsP3G5AuprL6esCUZvJqTzdNfVXBA0P
Z8po6j0Lp6iE4rFYovsMA+qvNWaax2ROdWIZ56ogiFo08PagTWEK5aU1HTMYDIwE
1Onwh8/+7TuMiA4m8oiH++hnegx2YARnoRgZwa6+cNgVn9bDsS2+1a3UuAVkAiO2
bRhnIcRbRMZxnfN1W7jTAP5TMGLyVKfwZO/mXhXS3j45J1MJcrt5cnVErHcrqH8q
zlsFOpJW9dQjPx0QoABkvFLRRF7vOskrdKGWm2d2H4uJ21NciM+0D82Ll+YYGhRn
iWNxwU74ZbpR8uhv4D+RjBaGZqqB4l7VuRumiS2lmZXqENmaf0GE54FVebuU67aE
FN70SQ2vgfnCl8TSGQcO2R3R9HmV2LweCSYSXFBRFt8FnwNPPi0tHvXyw3ZOZXFz
X4Qs0TFDCM49cUvNxhWsJzPHfOclu235OEuMTSJG6iBXrb2PM86XDf+3neEECHe/
3cWuXZOP2zlxoth7lX6qdhUqDwcO+vzgaYT+n3PdTGBupXZrS5Ex2PvE0g+MkDWB
Hb9t1LoVYbP/Z7yYcUnwDHlfQvgAZuOkEIKw+D6e0WpRx/ZtMzwtFil73PG2jbry
biSqp45qIJPvUuOtfu5siFjJYLHDIafQh1taNZ/cv9g3L9z1Uhnm3ZQDjrB37Wgg
7iDGfagUN8YKUS1WAn6694vMGThCwaImRGiqUpXnmZxbtVfUZqCk9m2v6Hh66Leb
clt7mJ0f67pLIdlFvbqg7lx5zEhMALGkhsWgovvML+6APuP8+QWiL6AroyoJzP2C
Zw2v4oa+2p/4GzTBIA8A0PztowHGoHYAhlR+QCozWy0kDQwRtU6zIoKMPFOM9Cnn
QnQP6ZGht5p2Lu4uFfQ8+uLye9iHlEKJutrPk9F03gODuj+rjqvVcyXaMZfimfAB
/BoeVJ4p51kGe880Yk9xq01ss6NE1eSanw8ayTXaGEU7bHd4HaqzvgGjpx8Z1ML0
sHbUoDGLJcUY84aCp16+gU9k5wrCKkQbg2ssa5HB9VPlZMI4ivnNhxeqt3lVmGlI
xItw5PdxK/I2RYKeFDpyA1NSogcalbRH7lQmM9Fk7SjrvCLQ+aXoelrThxeuA7h8
fGaWy3Jv1BleoqhfnTDPt50MJTZ/ixA1upLxIjjndh1A1MqJwPb4RSEeyM5HPoEu
uaNd4pDBLo7jzuHiT3P6/yVL0NXAvhoSdLQjOx2vN/AckzE567V31D6EPccpO4yd
9fgOwH8/66TzRjsRsMBs678jj57DAtd3kj9EDBwySYUi9GAQkMfE3MgG33vXT9Zu
Z5hqwPjxPdPR7KhBfGCxBNK+mIsI+eaXpT4/br1JIGLPSgSkPUvN6KaRz6ul1ape
hwKpBZpzJyJTa5ySrCc2UAS42r4Bk3XsBJbvDNQvqmteECAzcJnxFyqLOeR++coU
o9htrLpNtiQl/2wGjPq0ibAq8J8RoEVqrnAOtdbeP4lyOl2R6HuVH8Gz0PsuK9lI
LgJGO3LFxKLzWVRajlLyjaQ9jRD4DvgjkolEi60UkXxYWS5gm+Q2i3XCTroCU93w
OtT2/hP/hFZaNckhB8k69EtJNwzpUuoEb8KHnHuZ8z8TVJlhMiZ+7z3I9dPAaGdH
zc/LSNPc1lPh3SSTmekYVAh7geBiMjUnDC/i227WiFg8PISJox/Th7JVV8YcYSIZ
TeVmq6Qq3ZmybiQ62s3zEfHStDTXgy6Ie1iBfY3xRESt/9QvecFkscFnZPQRdzSk
lLKu8FThOvYqxPK7Aq/VSh+ZkeQo1L73ZXD1kbAsOfho+9PTSl+p/kFlajZf7t7u
ZRuYmuYd66b6dcP45vGpAP/CxWCgQPjUnc1QHcKkCl6hpq4SjsBABRCu57+AD3fc
Me9lqgEAhscfxESjI6O81scDNQS9JhQOqoZkQl+d1DiBoRd1Hufv7k+cVH/P1FSC
3WoWDmDwNgmU7vm86kPgxQeiVHbwTGrmHlQtuLNFX1awN3yyJiFBTAS5XZ4Hk7VU
17N0MVqQU8VD6wPhuRlp/1QwNjOTECggN6jAP38+I9LJDWlUhm2EQJt0ubZpURfg
goajfYcyDEsftPaY8HupXJK+okaFNeeFXo4BGCNaqmr2xLMTzp6aQ7pFAhA4DwhX
O1WBrszNwEUSD5A5N9l41gZYE1pxXx182juC60K5WPEsnG9mxSqA70/tcAf72eH/
6MT0scT/hWkUbD3ggAtJdT9P/CEuyfuf9C0c79LpI3o3pZpQCquZumPcBU5j0811
gcdoAV2n+xrUIbpCfdzxQ1Zw2j/KmojFhu7J5a5YyipHnACj8C2MZuaV8FLR6K2b
8qwcw3p8lw99ba9sW63QQB6Zp6kgEUDgjLqiydpAL/URQnTGnauBEQnMgI4Yg0he
q+yPrl0kHg8tuXz/k/s6m45kvZSD/XD1pRnaVXoq1D05rRxqQZvUQiDnaOqmRo5i
5Q+Eah9PT6+87A3WsI/wRKad9qaaFREUl8aBH1NyQmiZ1UPKWt2wDe2EK7r4HK47
xjhJ4C2mMjJmBCdzrgCfe0PUEvzR613SrjwLUiC4zGXwDHePSTXVLWycRC5cTBin
el0PEUZdIJKSTigVkcJJ/w+XTXMtJ4iwGvZUWHMJacDb5zYC34MQvm3c8JmOJ98u
zY4NT7AfCbARWoUm/5pSKIqWEQUni7nMT8UlLoWrCrp8bJu9flHIkVGbOI8IamvU
LSUhCJD2W80eKybgse/Qk1Q0UPHbxFWvxcjyOW3kOQb3XvGegGx2TRjG+tLzruFC
TK8/9WsCraoq20sUbO2zdGilMNAP9h4Fcxjev1ik1WfcdUwUQXmnCfTHug+psYAd
Q/Fr9K36Ai7E6PMKGbGEJu0fRNEhT2kAzpJTOQCvYK8TVAWKxvIxEVH2ZUlBcMYf
7w0cifsiHnyB3jTwiYUWN3a4s+dd8ZdG9dzYDLwJvFLa1kT4eq6WmzY0Rj5GoxEx
9QuJqjjUVQNZBwaurbiJxf6d6yQeJP4dXmEhBtFQmTKAp+AXjzn0/2C2zKMJptyl
0+mo6w2qcwiyedFsgo3zBrGwhGwaRLoMJkxMkjb9aguUj5stik9nxz1JCtK2s8VS
OPf7I75n5s2frtcNBuMwOZT24DSU5w/nqrJO5cfv464wxXvbohZUJwkyzh1/BFQm
8ztdaGsadeYRMYdlgcGfy1MdXSfe1okMhNKQhmyz336R50EJkZKD315pRQjY9mQe
euTjzZsNb7RGUk1lOGKqMxvMPxWFPKo1DCVkE7Hn+B4IstKtBSaWZSNxHRBo4ISI
WMZi+++V9tQxkHko9Ucf2t6Hz1RnhZrmSCrcWNluKwoCIGneA0ArZU9tniAlNTZ9
fUIGHJND6ws3c9gM9oP2m7Qbixn1xZSiYZYfEcZdrLBySp5Mvw47C6N9WV7YIfr9
/61SmyjSvwqsCb1l+YxL1I70vct65J5nsT4yagOJYnOLL/Jj8vRCaiObJM40mReL
8ThG/2r8hzh4iFWrViphkodC1wPgO7Xb/1YRq7UOb2fUG8rcWQKY/WB9xYVasiJe
XlE9Dd/cEBG3bTFx32ehyXSMTd8uoV/5sAD6H0ZDFmHvbmau6sapRPZu53qmwqjc
DhFcBv+Lng5UV+KOCI5jFbgmaYjj//NVTAhw9Ja2dRyJ/a+US1j8i3kNgWLZXHkF
ctapv3T+wqaawz9UUco4ylLIlupQwoEMuQteK2LzYxB81+9RqNJc/THL7j3OPhCW
RvPUaRE/BtQ5GT2Gi7Q35nIwJ713jV6tbl60/cxvFj5Ye92GyJEwCzjlgALKYVR9
H9crsfJTobXopK3zK4RPuQD2HUERK10S0FYBZL5KFQhurV4EQutUovfeYP7o2cGa
lydupKNEqkyurRdCoEYC2B+YWShIfKB15GaW1XIFUGfkYLNSblYg++DFztFmGOWD
Oq/kW3k9Wg7kg8nocdI3tAdCQIGXruS8796PdKI/V8isQq9AlbiEDnRF7Zwn2t31
fFoT6hVgdfXNhF2Kb/YnPtiH68PSXvohEsz1PR7WdEb+qtZ1Dp3GsS7zzrBeZSXS
m7xwAsToW2UgLO37NusxhkljRdPWi4vbFy2Dp7rU3cTleEI+sgivrgqRoOwxdDcU
zuTYD8F5I5UprZsb1v2JfjtA9aDgrUkGlAapH5M4MfH1jS/RwWdwMFe0oe054L4K
p8bV0k2ZBILrn6hVRSy5mHCq3yqsjcJ33+P8X9wF8i/SztPasw5c/B0PDbAeLQBO
rOTgoR666tc6YUKNGXMSXYvs8FCIHS9qafOCbNctp7pG1Ycugd6C/yjPB668wSbe
mpYY2RGmnVbuiaECrJsmDCDnKMkp3J4Yz5q0j2795W1wR+kjEG3GKkpuC4z+ZZU/
S0hcu2SdbDAMY5i9AKMTipVuMDi0bKfknxSioZC5spSTA0aNJ+6cZNE+w20Ov2SS
sUI52IlAC4K1GOiqIpubS6PmIFbfPA22fECMP5QThwFQoqigca2lmH1UDGlFimWP
vUqEgyI+CVZmMJBDdRD9hvGhyg5g/Qyj98AD0SkQIRZIepUEOo7EDjljB9WBkNQ7
ehJv/fMIShaEOdhQr+0WvQ/Qpr3SSuJNeWwG6VHNFFhh4ZPpUyp/fbOdMCWZDJxA
WMYGd1nvCyRjFbL9lnQyJpvxuxBjF3kudjwUZAD70UjgJkti9g0VcG/f7fakmMT0
ULfrEISKeB5+RWoAvYjohe4Lo0afE1ugmESD1rSpOY1yB+L1JC7ZPxR7AeX0WoTR
VUDS/FyLCxBRtULg3SDNtxYgvbu0qUtkrDwaCGf5zzKKB13H5UCTfuHXxWzByv6B
wyXGMeUtyW+ZXWye9SK8tAxigvl/KsKPIgGMnR/bAr60uGl1BZegqfdetzEOWgVL
MKfKxW+0IZWeb1WNFNjnU8TT/SOodmdVBScpfRha2K3KyBlTvHhKLPp0A/lq0t15
1SR0JEcMvkYVazfx6S64NB0pSwacQXkA7v2RhKAYhKN4phf02IZ2auSuraSabijP
s+R+L7SMU7AlqcMAaan70qTcPhN2a0Bc4+xIByAti2e3Cuk9XHn2v7gW6GfckkEE
UqJ3k4/l1t9Z2Ea/HgZ68H0XGdZcl0fVLxyWPdWK9aPm27UOzHcxs1Hw3yn/x00/
0P/u/l4gN7vlx5eCFd2NIaf3yyJ8Qip1du6li2/aHo1TJrcPejzGvRcQTcuI7LVo
tGZkl6hR86u9mpIvmqQBLOfSzBD91ECQcEpI1uwJTEpH/TU+y3MNrckh9p/ZsNT5
P9xRwR3UbVHN2xfE0Oqzth9D/krRpSpSxSjAIV/BmrzG8kX6Kb+UknhqM/WJw12A
oXt26rmMp8BLBVUWut/7nEf6ktUJGyWV045CUwakvF3Cb+x2Xz31j21RpR+8bvww
YRAVnPVhYFP9+nzgMKW4VdUP/C+DRGEZ5yDUEY4WzsTI6YwehT6/iqh4bLzjAj7W
4E60iLm6V5/t5mv6dEbJWa2eWk5PrgUqnOe0oPSSdP/6BYlcdgEYi/JjFd2gcj9r
eKaep22lSuMS3MZyb6IE1STkB7ccLS1XlXutZKpHrAr0GntKe+sXxmYB5mpbX4/O
iNkm02o8dkQN39wf/q0yPus3Frmw8+22J0ls1FZgUQO+x60DejNlG2qWaxqnhubq
r8YPfCKSSgzuAH1bj8if1tWIYejKj0tjUL+y56Saa5PLXQRbgPxNF5ve3ZJywVry
gSGEJ9mcKONNbnCrTr3TnHJ7Fw166ls2rhcC0nAMIju5fqMBY+zJNchVPW846lbO
OxbE9QtwXMYdQAusIL/k45EgF9xgKHqzc9Jjl8sTjbBnHrTN2tdsvwJ4dS8w5hct
l48//eMQ7XqgHDVf6mDB1AESurhGB0j5TNklBPVfYopX8K51EkjD1t72I0hUlRMN
npX41RLUJJST9aweE1qDRB5Pi39pPFNVXREDOLYleIC1Yz+pW++EFKsPlXO+17jn
k0jnapqqR5eDw/RadZ5YCrZjE/22d8SHs83qmxD0+ROqX6H7TF/WLJuha6CbPHLX
j7hklkn15Je52fin5OJEhxo/gD2jVzBotnrfGh95Cm0kMbGaxpnxLhi5dKWNmg9D
fegkBc7GzqnnzJcOMgDY42mDY2E8SoZyawdjlfAFKpnRVCR3vxe2ZY3N+bgs76B2
NAoO8X1UIYaIUys8w2Cbo3x9DZYxEk6mgDVIBNaCBRRLj2JOhhCbcWJ5vGMVIJJ+
d24HvCERkF0oa4pOdb1X+IeMUSY7C9lfZofJFxd6XnDRIEmIAWvctQZzu0iLQks1
q6tDV9ZVSb6CZ4PwLbQG+NCtq47MXFR6vNd8GbeBmTttVMlnIctwAaR4YFI/Kri1
+bxel/SrREHMPxXWesW9SbSthVdSln9HWiC/cqvV3vQtjin4BwsAIClbnhrE277r
Pi96NXiS17DYiopqUvmF7EZeI7ki2ujvWCfTCF7ltb9RpdUddIiFJc0/GBNEHCaB
LlP2WwmYi73cnaqnVwb2l7eIxFqghRlUR+OnhJS6LoJ1K31yNoDYmbiFcA33AJzH
JpEVz3e7dmL4PSwnOUl4wXYuOifUQrVdd9zYOz5+XkCFOS0BH/PNdeITTMpFOG4H
g+LhqeQOsD4wLDQrOD7GATE6N1eg1kwrFRvnq1Zgr6mWVbFTM22S1gxrGVLwY6NS
MZVtwrB0HQqI5hjPT2bCHu7jL5xfF9MerPZkj6jsNlMhZtUUoRi6iU8mVj1LbcSo
FF6ZbGAknjxaWKwWdj23WhBhAJhb9hZ7ob+MyVC1Y8Uf4uwvXQM99NIR27vtYBaM
ET4W1t7/nXDURNBgGyoJYAG33HnrsGRAPmAGVgazTURShRcr+LswyRKgkNlUc116
xB+plouEpWTbwWaC9XaEzYP4jncP+0RZkytlyEebnrOmAo30TYuzqA12gvy199Du
LnelWGebW4v9wiygVAzb6wyso843dApx3cWqocRQeGg0qxRgM+ABP8alEC6GI/iN
CnGa5iLQxel4vks9u27In8/Av7ADzM4CAmKLYQmUpDeJLFST1JxA4oWAgkGuT1pM
itK4qfIGbBLR3w8FA1glSeiuNbl3WTkUIXm7E4vUo7Vc476sPI+Lfkam35MqAHV2
T35CDi20nqKZ4j0xa+KouiNZtTMBjw4+DXf2tSjqUIucIPMfjpteuMuvw5XqMuE8
5Qs76pchksP2r7NY/wrlmVjYbF0l3/f+dZDlK4JTxtZhOKaPsMDDi6vaD9GQCo4i
gxPPDcfSJ5WmK61Qe8B9zCfiKQsb81VDN4kfqXHM/V6jOcf8q4ddJJR8jd1pr2h/
IwP5x10cUT0/buV9246PYP7/dnlJkGDudtRUNVdUNwUJj0maN2yZGudz/BEZdKCW
JmDnx3cIIRI9wc/1bxr9DPFkg6Sw3xeotbrjOQwpVzaJesGwmDpwwQlEc2gTk8yV
WB3lLmpK9D2eQOzIWNpCvzqQbLogVveNcPItAbkVR4H74hVBTcEvWWYlXWLy1A/e
QVE8+sNPhtbIHj/HFX13TfZ1MeX4P9jrtETKr2ORxATbsC6MKbCMKU9KF3E3V70l
8srD2Twm7rVPyFfjVkIJhOpHRQLkT/vdPQLMgD6yW2vvjBMxfFe8XoNAOkIjsPxj
inAQ4tXZRPZOc4mG3elMWNp76O96trY8UC06NqABgavvLonu95teowV9aRWmYees
sbdszAdk4hR7LvYhRMHB9z51nb2A2C62hPpuN/HGmkvEOh93Gfdcd0/mLxuiSZQT
3mEUE2GaJHTF5DNXGPjVwJlVUqDv8YWitW7wH28UxAx/0P9hQrjBQ/LLrT5brM9R
/4sIi1PJHAEIQmoFVcPLWfk2jM/s5LQ1cMPujl/pywU+8l4Kf34gwXVNwH5+Ql+y
ILhPH8ST8NiGADQERYEgbdBZTGefHZvDXD2+QCAVH3GerDeHXT5afjzImEkQX4D8
ibaiKRRsNX3lfKmx9PlbZDwUQiaIpOh9NZi6vkHAwYAhiVIq8UluOwDZlSGd/tGc
H1qrHVHALPD1T/7csfJZivv94imtoLS5jZdsmOQEyNrr4nJ0V1m/J+OpX1SFAvxX
f/yBdftbqkeL5Sp2kav5EVnGSdWYrVKcmTjJzEriSdDrYd9nLbnlFqiztGapaFVN
8p+33GreadqQ6Pmzz4sr1gUxrFUMk2EcQD9Heh7DFAZgsU/jm9kqUwBwTjbXOHtK
JPYpgcPqiInWjXkGHdHL2NKZRuZjOVCGHyMzEGKN1W72qGZhf5wIF3pLGA041qKv
kp4G2/9SqKkHHXTkiUMLwiTayZRBch2PNU/5Z2p4OP0P97mUjpS71qeNQITeOah9
oJvGU3kySTxpYAtoyWg1wGUq7W9VEMHf6P/gcDcHJzMxCGtxttgD0Yhquv3ZPXIa
WiufpRMymEG/cWsvY97YEK5FXELntXVKIFLD0/nuEMYLyA4Rf2ZAn5EQH+FI9aST
aHlQQEeBxeEfEze5hO9ebuiB4+jGzaBDYskBzDGo2n/ND2xbmx7BCf/MSIQb7YVi
f+rYfrBFfK2pzVb7SIMWp8WSs+ILKkirCxrxot96Vf/3p01lxv2uIOG0DhgOiKM3
VIEcDVzbQTGawK6oKj77K9BsC6Gh+nzMc0hnVhWxt4txvl+ji+jQzH2HSKjmW5nJ
HwDGFh2mw9mZOBR6QxaV6ZhR8NPBsYUPV9/xKM74IO/NVyGN1HdAaWpeqyIEvrMb
uUXtYmUlaQBUDO6D58A0fg5nTc+J0iV4Mxf2/xMnJQajy5UFGvFFajdeSNIoJc8P
vrmbeSqIr2Ovyk3aJhVuriyJux1agRaUzQgKGROycElFdiJUAdR5Sl7695SVAYhI
OuiOKgIS+OGngz3WOBkkAb4b/bXxvnWTnrFErHPBhQgo0xMTIPLUGeYAawuOyFEa
uY2GufH0RXKp7ugPAJoYERLKuAcMj5eeVHX9xD9ktRHEd9WPgTnXTdRfk3psQXmf
Zkielq9D/gBFPM3+Pk9Tz3vV4Fze8JfdwaODY/LZ8E8ZR+QMBmPyGrkQtGpfnxLE
8LwHnLaT+0O4TN3VQlk9CeNQOuNejyfPOLDwbPHLVJAUxIpCswmGYPxoQ0E+aNKK
ub4PDyi0/jhB9/W3Qbe6omD9i1u488335uBIxOzdweiLkhJPLXUEAgB6GA0HKKdu
eBhEFIoIoVxlGf/ptYMxgs3n9yQXK2T0URyIGpXy4FLAHiAV/24zrpcrgOhYch58
CnDEkQNkhPNrgHHEhvLYTeKdB9c5k4W04lWScmORFj+LNZivCP7vVEDENbxx5/Co
Dvpe6LLdocEIZfnKsFrAw5uOLFfCpac4hWd9nD7QFBn2QuxKs3qrpw85JdF4c+HS
9OtJbPVDhERpbZaGdHMzRDUFFVJvMlKXhB44Bw4YswKmYJSPTdCN6wDny0C1lM1s
Js9LdckwkdoHtztG7WL2HTD3p4XBU+nf+r1Zs6NAS5O3L2GSi95Df8jxxXIeuhao
tJb2cdVfDk9GEKG1nwFYep5fZGLLSOITuGbaCqZ4oYKMGEuN/l34JOi+cMnpJlvR
5HGUA60HS0UujIXEiiwUjIO6NS1ADHY1QbHGBvKiYJ4va+8RuoW8kGxiuFgEk8oK
3triXzqCnqeM/stvouCy5gQPnRp2p+HaT/7rYVTynGtyaMvY2E2jWYP0Ods8GhhT
6Y17tY4gqCexkYdWtbqEIBpmbyLMVWPgcwyjqL8gFvdDFsVomdAI+SsU4ehgCORc
3LR0IoXGC7f734U0VlYwZ2E+0kihMVqM1Zk6oz2tH7BrwOfF5RMr80iLH7lEo9WR
s0EI94NCYO1GHWQJppRJEIhUF55NDfzzZXMQhncJfxNEu0Tk3rLCZP2ZjeRIz7SF
YOpgHFaBZS/ylnu4ka268SBccR8Bj9Iq9roE0PYCEe8L2+kQa5kGEwYxnPXiBWuQ
VXIFWfl6X4vYaFBlGczQgx/qIiF6bTj4Vd3qH/mI6kXbu4Or+DCxfbqT+bthTWyM
4ikaVB85nBIDi+NF953WG1PWsKUp3DuAXB883UNS/7okiinKh7EnCByMn7tmFcfz
1MzpMtvkIEUWE7+ACoL6SUkh1nkebALofIV3VIPaJNgOe8snlEDfMBdaQQh7TuXJ
DSF9XVcv+/Ihhj0I9bx8Z/MAnGmKTiLlvRfxqptTB0mlmr/0mEoz95TIISAFd0Er
H9AaWedfpZqJ1xVeAF8s6V0zjzJo8jaFOyyqJBlKElAr+iKFRSePcmG5g6y2ZYu7
yiYwe8RD9LyN4ymt2WTYIkLLEl7wjg4a5v4eUt9R/Lb7E7w8KWwjJG+Pk7GFXtiT
AuCL1i6k+34XF6yHo5Ynzyk/s/50EC60WmpKLOin3ChJ/z3YPejFML+lKL544fDZ
uOd8Dz0H/1ifKkxkApc6jjr2xUBRXYZh/8Uz44yxElUpIyA7DKedm41Cbu+YD5Ro
b3+mtSqPD/bmNjtpChPnbbtizR1geji31pIIMaMotCZGBjKk5x9osR6wyjLpnHZ3
cUJYO7OTBWJFTroLLTmVs6iORB4DKfDAQ1XkxBWxiuHuUWtlmaGCevfyJ82TA24o
xUrgqQRq2SvBOdHGi9iHQEWn65c7thhWAqmV1aYm3f1KorjDNRWdsVB45my37U/s
3Gr0Vzkqc0KgrPzLGokzlh0eIYF5vIOpSvNw4VHAmL/d9kl8IUEdz0gbXlKnfPZD
Gvy8GUy6m5EIPvQNyJdXGAmodS7mqcyUO2IFDQ0L1jRYtsY1p6LqpLLUAzOVUW+6
+ZRPXbgTNnRhXwHbnzKvhiYMJq+NgvHTB4ElYgCECpo1AOrhaoEn80lqR/QZFhbS
y7cbGnnagjsDssm/AqvNGFlHUyWBvqGhbbviKUAjp9vdWc8lGdwjaPeRgThHSxGr
+aMjYqSm3EipLpBUh8uDN7LsoSNvM5HcRyArtjLc7RFSRucJ6uFllZbVx7fEhVV7
Wv57mZKnZscbjTJy+bS5jolA3yngSx9RphBaBb7pakL2g8//WuC72jlOODTS+P3X
t7HXsPix7dD9rxWaWpLceVhhowKTkirWBjfvdmDQlu61ePhJV7e/spxqwGTBFI4F
aiTHHMjfiQxlEH801no52Lt/c5ZK27s3PnarMnZXNrPPa5yoGbhFJMf7lArpaWYQ
14QgHuAKJaW2L0iKuwUlRm08keAxr/NiQK0qJLXlir0EhQLpfOmTR99Ofi5Ved2C
C0rQpof8RqCS6eQP3mCM6Qj2WF1sNZvk4/R3q9+nEYnQ4KRjqS9VQY/BJdROcEAY
kNc7YaVJbugbo0sfdPUwZXFho8SACoX5QJPGBG3CFI8xGmpxzwEhzezcmQDY5tC3
W6G9EIqjO2ndvQ2pl/mWH3O3Tis/omF79L4BlbsBLTsBZfCqN7+cW02esIW6wX/Y
x/plRYqQgaod6DOC43TFKbaXw4zvDiZYtgS2VPe8STj3ThwyQjXiKlHSqvx/jtQo
/da5uyCAfXgD7Jfqwq4VWYH+15eYmPg+m+qtdffgtQoJ4bTPk+WNqsnNfjJnC7Kr
h7vLOo+fisyGb2s4m6BwG9ZXNahVSJVhnj/KGWhUXNQF3R3l8uDKqdWtFKkn4W3T
Pz91nB8O/x3WcbJGmOJXx86Yd4+eF+MOZXRB/XYGG7fCwIVDg1dZA1JEfTGyyVf1
ereQNpoblZwLmafdlK7giP3M+aCleYdjfVIcjOt++JVeACABbLoPEhtanDGEYwHh
h/5RXdqsJ3a88d32snB7Wx0OTzK+rtCCV8vGOuR+3ZzZ2tenk/RiMkqIsArmQN+C
QPlnHJrmUBDitIZdFshNF8ne9i2W06wnEx93iDy3HBP9DUP5x7/VP0sohOSAW0dg
6YjDz7OZs+dbuxceSE3+aUA1hQkqVK5p4DYv5smyRT4wBqPAjCjrgkmvbssN6X3F
dNc4i9EEqte+eJXweivqK91hLxgQzCWEg5nQTPj6kX/WuomT55DaWXb6WIaSWWlV
BX4q7fmz/VjZCf0thdk58N2vKkBNeyEWqbgoSGmafzFMG6so89jbb6YjqKMewLlA
1sC5ywC7/aSeAInhzD5QOl1mwXyLVbc51oVGbp8+uBf9twWbb42sFg0198FdK0Zt
wD0fRJNQqnSoV9x5IlHOE6vCzApkD2+w5mJTEiuNINbQnfDf6xLb/flF+MYH6mXT
1vAQD5AeZBB0tg6eEPkvkHrShv9onafh6m6urPj+EYLpzc0WMqgNKIc7R4CmnZf8
tDMFdHKJ1J4lM6abvnIVWE86QQwcHPLrrBNumFagTJSPLWBn0uiIbziFaxQy9Iow
HsxNE5KokyAEoWSzLavV8SPfBrq1eeIb4UJPkocQuGWDkkmm29hvvQbtT/jMp95N
CK3ZSuUWrD+m4LiPOVBqMuYfD6cTzIDgTkmJEx/IEid9LQZi48d4C2PojiDDYmHK
n8+zxiUQ0828y+gOJ8PLG3+l881yhfaiNAN3hTE9LDK4h0zRGUiCq33Rz5IBqrR9
kweNnykVLAFoHpxQVS9SRpoiwZ6lv2kC1GeWaZ3hPC7pm8cpnUpyr5lTj1d8fbob
ndlMzTCylbX0nP7a/NGZodXVGeljfF3U0gNvDVum31BIunfW3QTeiq6a0b4VOCZK
SHjDLytYcGhU4dO6x9SHklBVKb6ZUiXak6/3Li3zpSn8BvtJ0b6SIb1iop7zgXwc
ILDsd3ZN/d/y99y9Saq6w545Op1u4hwdYJPyJoSwfnywpn6wq6/3xrqANwsnTZPB
Nr+p5v+mvK2R/ERk8urSz4HYcpQNlOd/dMjkfBMxOBSwuF8ycwi3ZMJikGUPaSK/
qvwwsUZMRwbLC/kveqNhGKp8QP6VkrUIH0fv/InmQZc9Hyz6YTr4TEv62iSSXMvw
qs7WAYNkGPaPgetMOodt1YqdBERug9NYzM260FiFsEBk1zZ7ZdRl8QLe7McmGvjW
t8SNc/TdEFzktrQGiroPHSFQRHYmjLmjW3nsvov6jQxELXdFzEGNidXNvvLYSqnc
lMHrQtq7Z+fUaVV0n1DtdEep+NRrDNEyg7Rjof0lG1UvZc/7dy3H7rRP8S9bk2Bo
maJ3gDyim7I45O37bfp9a4QYDrCWYsYAB0oyjnQB5i7cmg95FRPFI32qd2NgK5Dh
Pzyp+ILop4wYShGlx1cqI+CCDa5CjMRm7fWfhZGERzpwzEue3FR6iTR31HWQh2lH
pEr8m9pJBtApQBq92aFsR4fv7y2Axe32C3UMNyoIxgalqJpWhSQ1Phe/ybJ+CIvt
vv17uls6DMI1uaQ/IivzWZpxTsoO+VYpcPrrnJdt1H1Lmt5Wpl9oowQ8cO56kalD
qYroOz0RlXelFXJ/MDa+zK/Xw4J8P3L5XWGbf4zNr0YRi1s9uhYA7zpIkNMUiMdA
oKP8+djyWkNzuOXZX70RbhFHO/AQlUvGnTEaBnWnjCO+PwvG1g1gWtyIH4N2RLkU
IC9izjyFSgYXxMulXGPYruXYyCwknW0LIt6Tetqt9iwgdDPxVmDimIJFT9SoEsRC
7iVQbHvwLofgeSNTDAQlv4PGbjaNqKhFHuuouJ74V6CK/gO9XR6W3OQSmwk6jXP7
bhu6HMOV2GcS7uehOoOmlCrVXykH6O/gNzNfRDHvf/+6slEVhCwj0ynzItWu/Oeh
+lvohmlGvh9YJSVJfqQ2t9J4DAwFDYVm5DiiQT6D8KHYGdSl+8Y0WTBLK1zeSrF2
XHuFWyoyUM/DTto9GSBcxHlas63l8OKADLlt5kx+ySvfQPZw4EwgPB/SdgC0ccCh
gY/MBx3bnPL7Ho2r/6Un2Sp2nUBnmjsQlaQZQSZdZm+psvtuJ7NuICE9BdsDQat9
eGuIFYHgUy7pBso4g7vD7tNys0dhnxtitoUIEcBk6miIpyExpJZWUf6KxpgmPZqn
yhRq+9xoLHUKduZ2MWQLrpA78+TLvXXFQgB1g+B9+yccAWYCHa5M2flPcQnAcld6
GiBVG/K44emn0uXzCIw1JbEoLWrqYXkBNvgSmriz8iEaZT3jMx9oPz1nr7/UGyAY
eeUcGahHGRnuwZ0KaO2O9U8QoEh3Zr0tG8uPmhlpRvwpJgBZEvRWGNtpTvwamHTc
Xmd9vG0emioK7CZTeW7mex+7y63GYSsLzHfAatkyuWacE6ko6oitLDBtG8WUhhRs
ScLfg2HIWeGWdKAP4yISYGj8B9EnraIIrOBnW4qLnXnzx+bp7ds5REh4hiwgN//y
HRWW7+IXb+SZBrl/dSR0Tgfw9cpn0HpwMmWkqx4Hy/mqA0LuMpEm4CwzfCtC5Sp0
6uHRy3L6KMGx2WlPjJlJxU78GNdgdOGLgtUSpE+OWqG/v+7Og0C2f7IDfNYHX4vS
AecDL0ZdXkjosO4IM7fahfEmDxbkV8ghKBgo3BUzErYObIhESZMpKHj3eBvbrQhQ
ZwkravO35lziFoYw2dRPaoHdbrzngupqeXORHnr8ql9yZtOs8FFoYZN3iQf9Hfen
sa1TQ8RyY+IVXa9ck4Ga+6BPAKPH2R/zI46JjXGPvFNwaOjdjSaXm4Cx+3i85Tpf
+S/9nRBOP0RDvJ3iVPaRaSRvyKZn+olaE4hiFQWRvVWtIcRM4zQzd4Blc1gxw4GH
HE8v9ETfC/FpAgOEM+xUlofMBzUgIIr6cNZ9IpHcAtT4qMl9LunBcMht7bXp4rrz
CfRlXQTXKd9wOsAAsciB5PW8B3vR+fboKn5xkUq6krUZrr0fOQbKjvCvWyBuiWtM
Ep7Quwp/Qj8SfQNTPiONkwKiDUQneonnN0xdfqKo1slBDzKg0ewYazLzMp69T92S
PSlnhiFx1DoF4KE4KV9UuTbkWo/TA2n43waO0SHbi0CtlX4c5ukHQNZWHEXqQ0Tc
wt9DYRcAhgn7cIiJig4vClvfqjykErFhcbufUIT8RyiCjv9pPu29cGShWGAbHwhG
y/oEPGbSiGAO6QozwHMetl6T3cYb2AuPli/NZe1K2XMWQdKD0VuvbITReJP/2W26
MloaZBoU0OjcDQuZFY1bSnVgA/0U4zsA8UiijuIhMVlGE/RjrjyLaXzwKH9kh5Di
dgzBzid9oUi/G9YEe86+u+kQIwjYVdmY3Suui9PRQ6eJ3a5KesbsgqcQYYseq2KO
NyIMYKs/t0KWX73kVKsb98cLWd2oA4wE9ZWzkHtmNwFZxJsN3gD9iVxJEdJgYBU6
a08F5nAM46kgKjDqDgwirMjtcnZoy3aw2pl9h0Q6E1CVB4tLRlEK1VGPEb6ljX0W
5Z14evE6NBzq+/M9+MMnjNyeN9jGCtvO1+XT6lLCeJnS+4G/KZ09+Dqu3HjnKJXH
aD8n87+eCAVFjXU/L7dxtqhGkCfGFIGdAwfFlm1v6xxRVVSzCAPQJnNdF7PLRXJL
O8v/QOuzyYCXVP6ZlTBDjGacfxV0oMSo8lAM5K8rwK7zH4PGY5Kkewth7CCE4PfX
uDOmjr2qj692Io6SgaQNOk1cAG78sx8QYgc85E4ruXGmSqf0QjFzhIpNtd6YLfKB
FUHzzxOaXjC+QRA6TY5W/m27B/JfMNJLE11F0J1VFiZuEs1t0uyjCkvGCm3RMGnI
hwwFp9Kz4Nmlp+AZy6cWuCJ05yyyPZNDVssbckF2voueAf3VY3CXQlUsdVOzGTpq
Y97QF42L+rJm+mk0SAgllMHgosC/fBwte43OmObuENdjlpFX4QOkPE7zZifBW/mb
zUpyWMRVKX/3ssWaxFYnnRKMt5mQdK11kK5w8HCnOTDDHSnRLIx+UW/YlBfJZ50W
P+kUeivuE3SUTqpgSxJoc4lJp/4BKqIb28huZ/E96DvyXzWib2kOYAn5gvDWaspd
8xaWeD+bUGASPtZOrCsTncIaANxZaagQxs6vEggeAxxM6QGKdHIBAZlVBIubI3nB
y/pA3oyOQMYsb5Z9Co2gOZpzB517ZIoyC2hl82PVbj4ZPjRYAulkNGVckrPLtEJe
39qakI+Pos1xykmib0O5UaEbJNzA2aCj0dop7xEiV1j62dqyxcM7tXhPQqCzAg9O
bGeqdBCwjUeVgodMqvrKhCQkruF8G5kotlX1XR7pL0oEaIO6AKLSmSlej/PAgc7p
PCSUaswttvtia7AOYevYSkf3F6SUOoJ+x94/0/NXsC0+QdAvxtLgfyovQFW5frDa
soM1zbqL8LEToyTdMH5YzxA0aUb4lhQQptxrZErN83+MFIoj5crPegPyBc34yy0A
8CuxLRx/2tHlV6dcwfj7WAv4HRqFAna08H6XTU9YddvsElNxJyl0YOsjWMBvKAJt
PUN9PKEQTRgU8YLJsPrGwM184YNQeq8/rwTrrewimuhO81jYW5fYHlPVDYdAc7Od
60lnIAihCCU5tBsiTwGG/+GhyHEwZ+lQWcCnkss9DDavWqHFWhZchA5AEfcEWQwT
+gCKEobTQ5X/SQTlDxGwLxIyh5HJELl+h/jzP+CcPFAWUaKZyQAs9628y/P4ObSd
o8xAfZiE1ohW2BdLe/XWfSUpu7iHuZoZ8gtrXp41Q4DPaFsagdEmvgUX+XmWdURK
BFeTo5WAh8joRB8zWXvmMQprJZAdVCRzFTyARXAeDm6pLHTEwLpHQrXBPMkVAJKX
uxJ1EIXNjFHLLpxgMKNtYDRJPl1ha/iUldp6ic6zfjYyEqj7xlFyEFwlhLYcTWaU
IuB85HMGUJ/mh/kWgy9O63NEPmReZg0AU38sCYoKj/x2mIOIaVLcpL0FrxOMdTEt
4SnhSpY6l3nCcLnYBsr7bnJkZvOKd7mOqtPIOQU2DiUEfZsQ8gjaF1r3ee5drWDA
n8pHysk6XpSquJ+PqNPqJjfTXiM3LJ+oo+5dq/aczW0tAwp7dwhpu6TPQJ/YUL7t
9z60otH28bMsO9CGdDDuvFhpliZE14SICaYQLKoTQMUZnQiLp9y/E1QmTQfRBgVX
PpWUaBLJKUFJjZKkiG6+qNLe+mZJsy070L8eX0eFImp2Sa7gngr2uJt63gWumYTw
5GD1kRAFS4Hz7fLKiD1Qupyms+5qzzSD72n1Yy2BhgYZhG3VKg4v5zFxS8UxGLmR
wQU3bzLeJHRKX06qBU9dq8Rty/44Us3BH1T7s+1UVniE/e6020NHB2EWpOOXupHs
GQqTjVHTI1FXlgakMAjZ7VeF4TtN53IqVagEydTwoc9N2FXBMXquEQfIPISe5rk1
gwqDLL6uXE3Ujo1IYGtPYb4ZDVDfsaGpr3up0Y47xSDB9kJ+DEZbnKDCugh78TKG
KOXoyIMv5Gsuu51YTKQc9DXAZd5HcR3IwCMKRGWkl4ryEm588mDBvi5FEll1xBiJ
LZAIvp1L+wdlPY84AZg5RB9mJuNpXvO8n55kqDFLreVgXTUfCsG38JNuHlU24QaA
MUGhEkIdn0s5OTpq+kxtVesWR4cvRKbgl29QnsEIYSoxScagDKGFBxNCBiCi6piS
BthyhMIgSsirr75DArE6rQ==
`pragma protect end_protected
